

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GWT/RJdN/UcIKTAhVxs3scTnM63xEPkso8NeqXOmx+sudHjUMJ/qSt5GFjdXAqexLlRND8lEfssX
Q8fYY8TuyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J+phMqmkYiPgvjvEjlpcdWdxzP+34SmYIPyc3dLXEqt+h9EhMcqfQg7r/svpEBV24DU6CyKyCXke
3gZaY85pXANGRT/lW2K8drptf9l9vYajWMSy/HjvETFYNanQN5XDicKd40/UNr4NV+8K3+zJSD2+
6HJJVC0iWa6RgWieT3M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZrkwjC6jJHChQhf/EDIYzNRopX0ckXH4NL9s7GZmKhZ5Xuu3xV3LqvLjlAq2T+/3AXtko4HEVfJk
jD8rEKHAwLnqMbikHpL2pup+LY4/a45y7duxNC07dpJvYX19IW6mqYLKEJTs330XVwBLE1KOyaGV
xhWwwqThGo1V39JpBwMcpzmL4YnxHaTlERiq7vaoQpYAMkwdoBVpG9MMAn3CbeZJI8pLk/zNkztm
rMeS9pshqNVtzdUse3pl3EDxWMB2hg/4/G9fk9okekAXBV0rv5NMqf0xPrBsTvRJGO21aW42nO++
dC8am+sI7nAhoG4w6z/WxE1BGkRuZGX4CGhIDg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iexpjlh7M7dlTcv5seskQPlqyHreGwsr94b5YKwilWQsfXW7U1V2aK3O1/+pXS09S+pTH0rKoHNi
ofASVdK1RB4/i9AYD0Ihai7zYaqt6eRX7azypmOnO0M/ZZIrM+63BHWcDodlNlh86PWfwaKQSqJW
hLVuOmY14GXZev020lRZWg+2UhI/Cl3c8nww44erkAvCrpxmrhaZg0s2YPKI/KBqZbZHwn0ufJSY
5EPF28uCCS1urKeejeaSBUmimEDyf29zU/xFd0fvevSdWXaFhwjT2mOL7DranIxEzj0yQrN0jiKy
Towa0uazE4xB+gMrElDuwpcw6ZUMyEBsaW08mA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DVPBxTgKjw13z3lZMl+QMKXV/uHfXNCgMoWbgQb15TKXtTCmkLiaCYkk+UNjnupib1FZuwkbZs4q
pFuDW3Z3x3poQoD+4+Z7IIYAmkcV2VNFgSXWGO5qpHWhRfkulPfZcRStTLiN9EUcwXJUsLi1Rwk0
oFaVSUr3p4Mr6zjC18beDCFomH1w+aZiTDmIDtnqdWVtxtresAhXiT6k51hdPESOpe/yPCGrgQj7
cckAkNk0Y7ums+FtMhs5xsfKLV6GQGr8vql+qoCmnMNbYofWKIq3pY2FrW6f7ZGbFhW+vgaVatOo
wR1vGhSucCD4x9efRbKZpd3HOhDW/vOAo1pd2Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uIb1xi/b1sGS9N5+ge4ctTMaXcuHePw5wBb1FVa9aecf3hzk8F8+/rWvK4DX9IjVKEx0PLXI6xjb
IH/rGtJXdtbDJdBaXxCtQZnZ3bb8a74BAJHYm3BEextG398AX1ZCOiiun/unyz5EkREGrSg9f1qp
tvP1wCaUgYbP8iAi+ak=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qK9lK7oKxV9h/658uwPcMAAwYeLmnKNpsdduH0hJUA8HIiT0JfF3YHf9Z/+4sugCSI1ARr9LlbO/
o+J2NPNqOXlyDgJW0FGjeX+G4wdX5LlxdfSIcRGs2vzyXQiAWVbMq15jqJGV+qheK6QIsLI/qwOR
naZ46kfkwSE8kQXhF7WZE2kD7kLSTF5QPnmYFPP1wrSHpjD9hfcjmg2768Oxg74FqPuAHl6cX4Bj
Enf4+hzQMQ+IcGssYzesFwyeHIqJFbufwMH9hDnmz2bOveVtLUI33QRmIvvIjsEuvmQwCu/AC3gG
UyfxcM7HSiPQe9MbxhcS0KjoubQbTx7z04URRQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504864)
`protect data_block
5E1d0HeB6J6AfXvWJcFl2ETasGGXQvta8al9KWrl0emoWcY4zrRJkb30j4gJg1NuiSGEnZJwbtY3
KKIJlZPsF15zK04/1T2Uoa5aJtNTw3jdHZNkHeDqQrrR+8qi9m156Cm9FhwQQm2ITIJnJkoPV3HH
fHM2v+GQ40zIrt0AovhNH5+kWmt0fqT9TW07JftTpuHPKSJtvssq/ROcgX3Ppg2/vaLvIXBuYVDQ
JkrxrleryL/27nFuaFMVfuL3O3ARylYO+FzaAXzplE6LfU5rC2usAd0fQECucK+W0CNnfcNSiu04
/mv9fIP0ME40h2/xBvSg3cRXcsbay6xRRbpmrIbqwQuv7/rMca0JW0msfDXeVxnP+n/raWfA7Yj1
3zgRPaEDrklYkk7Yo8XmWa28bSNiPXsycwVITERgGl2LeIBYKOt5CacSkgeGV0Btp2Vv83p6dzYU
L/c+qQRhMUTn2kS+Ua4+3MWgiAGA11S4+hzh9YzakxJYgaEWCULuYBwTYWIlrkrnXfkjulpk3AMX
j2IHPsK2iYJKGViMQk7DsZZw/J7kM26StFtVm8K01I4nId/E8QQ4/oEKItItb2mWqriiprqc3HMI
arQQSdjX4929RyGSD8HpVc6qsLo4GwPg5dPSswsNAffP9vzC4Bx1A1u9xodqaZTCUJ3xsYHE0+dK
Wn+W0LUjuvz1niTpBTk6VTvg5gBFQr2Ki0nYuC8SUgQsqqKPFVjTcu5SKkWFEqCot5KOLUBr+cIY
q51x8cK3UO8ixt9qBR/WqqHV8vEjB+6DTSD4Ed0M0vGi38vtFbe9F+DP2uI9k0I+c7PDXDbwuNzt
dWBqkwI5qsMBGvgeuScGlvY+/yVHj6O7NFgvKtmTeElG/s/++LTAmT5cyBjqEmSq4apdNOgfZFNf
HemV4eM4V7uYHO/fj1ZLYbO0xWUyEbH9b/QSjDH2ZzGP2S4tVyHuq6zP2Cnoumts0RsHo5Tg0xjc
MXiMHSE/GPOCTPDZUpLpZyffysG8H7sXJZJUFas5B1+tm11Pc1BPoyA4BDYJUu72fvvyXOVTT9Xk
pfLbxTsoMFtfE5lPPv84hiLsabr8icnuJCri3HDOm8hd+YKmRn8bzOaRkXaBHhH0vyaPxb+/Gb7F
mKJgyvP3SMFwWHs1tHHxIoFgK3BUAILzqIA3zDLEzZUn96/WGXF5rbjU6nu0yLArf2VcXsgqaNYy
6cwo36xU0mV6lG1Nui/5KpF3zrY6yWlUFe9b3dKt9jRaw2BBefTHUALPZkvbiydlNZbkajPRqxwM
9X8ZaTf7II4fSnJ6JEvQRTq3vBRQZ/+Uqy1zOs1756/FO0OouDf9zMEkxuUUOolTcymdJ1sBOSMm
mV2k77+ObUoQ1WN0dAoFCXY1V/FvS1jEo8TUxDC1JkN1y2WXPpTjUX6tWLnI2Vs8tPQnXnemDrX8
sNahS0MpAmdg++yLe/mIzOLzcZYuydpSjY42aLiKaszt0lxhIb/0ARI2UoPSBW9ZcRPyeYSKKeMS
ckwXrabnhpvH0BGyxzkOa/96Yw+uXoa0yhtS/Vq91D6Talwk08e0ZPzPnWV5MY2U2EzkVyDoK7xB
dCJcuG3QWRh0VLtZRGX0ZKwDplObT3pwYXwL8AWJVCdvTXEtCJENVjJzEusxOHaBQjyu768IW9iy
CJvhKzKY6xeGcpHaVqmVxhhhRRfAP3Y/DlgRq4F9dqfOpXPHGnwHOOsCcwYFALMXam1Xr9jG/dIX
Ck4vs3vPRV3ukugBTj5IIiV2lnRdiL+5OifWcv9c5T4y9JbG9pBueqjryJSe3C0SESAn/Qd44Tna
oBs4e56nEve7NVmlvles7oCr9N5AkwAWOkZim3a2pxpnMK3+jANWCc+j0GuoZRRS6LZWDLyGmusK
ruhPhrAK6TKqfD4nZHSWmg5LLjzPiQbCwVMpzHw/a8agESx+iu/GSCLdw6Gap6vuzvxtugDq7bHf
FQ1bDZwFzaizM2OXP+1DaAKa1/d1YC67WgyEfwJz2Gb9CkzIwpcEzeCyEnxgiRNvaJwNe7veSSSz
XVtqzcGjhtG3AcUfReIq/05FTJXqbZ5MLxf+nU7sOWCfGia467LOCyIQo4vBDVkKTE/nJ8/MfyDJ
zVSX0/wMOPtT+IHHarw6EbLRQjOGww8xIasERcuvANNbohIhTvzpl+gZakcwc6ExYBPuIdXY6TAE
ME+2kNZ877jpaA0qHd0qfWNSQHo1LpOBkzdzRdwsK97PVYBeVWKKkpW31SmzynwNxz2PEgZWJuf4
1p2PSNrmnCnes0jMdmENwmqD4xUSbYNeo6Zg4sKC5DNpbT9aJo8AQPPQpMp1V+NqQ2GdXew7dxXR
o0jxAjG9X4lb+cgREzTjwwvnf5JpnJJqs7Q2JcqJLAxD5wfl9zFWCb7g7J+Kg2j9Vw6Fa7DV/jRA
Q3RvFUROTgr/F5wtmxasdBmtJz1546Egj/8Cc12G2gSZwnyoYfVl6WWUTAL8bD7nOJm1oAb2zwWW
UaQsVpBjofrEs6k1mcgwxdeuMcqPAbHxbnCm9sYILRmnkk+QagXRlWKX+BO4xsBv+s9udrS1RwDH
QJmJOw2kABKP+ooQX3xeoWMnpxKZqirhJGc+KiDDpC2wsSx5im22ZsG88lkrbQvRyCZvstqKirv8
OhR76iEFE43PyLSJLE664mX00I/weUduCnhKE8UCEobqBradcnzCIfZy/Bl2GhPEJEWe+t5cx++X
GswUq3pzvoGZXuTaiGmRce8noWmY4yrz1nBikazpfAfCsQBaEY2PXqqYoLA73qTJEKSkEF1RyTnI
BY2ZCON4iTHqdhRjMvN4tCHVvfrcHGD2qrVl9V/ZMjfx8a1czKxscwL2jrGOXXwTOPYvcPVk2amb
2aFVUnatfyp3gE2kFYvlf9op5KqTNhH+oouNXJOZ+KC2pIyT2vQvhPcLM4ARfGrTdQUqVFayclSP
/675VlTn66TBPA4uFZbwVKEvpEWoLsuPbRRkXzTefgpJ4jpigH1YoyEy3nQYlVi6HDUBOcSF6yR0
iLRl/JpTPFAUsMGrpg35EmII7U0bC7G4I7xB/VUwG1+5W+hgFy/XnfVvzNJua+ttojz80YcIMCBD
EdaZeS1EWwg1M6r8vZXT3OKL9Am16NQl9mf4/rzETJbDRf1hR0I0rE2vxGWXleKxsgg9gfS3AWB2
G5kT8/7h1s//lXlIm58xdOfZBJrX0MJlWZOHMhgpyfsDFCwi1xXHCqtwmoHD7hjAdPAgQnh5GRj+
8jjpgHZYOyTofVNq/ftFxTdtlBwcP5iwfsVhXmkgZpNnyvOG8FDZsp6UiNzU5rUTihoyi042DbXs
hglcDo2t9KmfOD5TdzFsb0NmQXuebjjveHfmIXolrotMxg6hNccGAz3i3kfHhNKUIpWTRLNvQLY3
KkZOKt/XVTEen4gOwJQgYpmZmeLGjby6pZjChZGLZmRsdWb9eVOe7gTkb8+zvQK1BomekB8RLgmj
PegtsinPTm3eYegMIyPNBZhoq/sBplpMQjITavpFrKDLVjyGYyaLBrQS/xIMpjVDKF1kaTSmcfAJ
V4IE+IiuEbIUiXqk4YeeStBYhoTdNic/FFaF37/cfZ9KIiiVept7LHV7J4+d/lUh3XNSvjxeq/w/
FF/h+UkAKl4X2HQDaNWfV8YlAk41UKYoYGzbldIY1ty0vjetV6/zmBhVCehoq0brxXn3ez6C6x5L
rEQjSLF7mTyBdhSTazX1XG7cZ2LlJHQoALm5jelTa2KN+8n2voDy97SHswvmlaBnLbShfzYW+KJk
qJxYQksBFGmonvoTV1wfFj2REiRPbZwdKSGV1D9rr9I3cIxlZxPisrE9hHvH61B6jtLTmnTQhADi
gY21PV+gX27zs3gnnXG4/GQJJBeYEqVDiDuqeuGDPrf04e29g23WoabF5JqSy8QmIxClTAGT6TmR
EShl5LcKwf5MhNQd5o5rsZJQRgqqeCeCdRPufI509ICRKViJPsype4R7J15z9mjfOCt/jDyO3fOp
RNJMV7QTZq9JLPLzCcBDNl4LQKKGBCQOwXwSzZDW+M/QpVeXfXHh38vQAH+vizNk1OwUcjVcwAWI
yrwVNxWzgqJEzyQHv+iTKp/1eBv77gShNk/DvYweVlU3yDzrBotzOaUy+f5R/CaAQmK4ifLlebiL
UlZ/F2pwALqWB9sx6t+3LdQ99OknkzmCh3qo6iNzvBaeUxNes7gGUXXdCnJBW+3IZ4dx/N4T+ZTY
1QZn1jaBJFiIWVPlxcdh1MkiQIGCQ3/iedOH051zijgMbQy+E5KdtOcmLy2mJomEe8tKyVCTVFnj
l6v5UDzKi6I4It2r0DjbmUJ6719P8Hc000GL6d9XJ2pkTx6izMETvEbwpwmwE6NmgeqkHl5WAP4s
Nd2BGEm5iCkOkJPWHvXHojvv972Dac/W5YqxmhpoeCQiujcUuWiGRKBeVCXifmbVeZUb7PAUZgk0
NdlRoMyx0yyhegXavA5piDVacvn3kpIN6wElp1MudEYp5w0DKMqTeKPqDI3XSjUysfv9JZMZP4LI
slK6HccNwjxqN1LqDQLOO01DejIV+2RWy+VoyAFNyGK7tS/mc9cpt011cwBbWbsiZTD+8GTuJ56B
02p72Y4nMy4tGOfjNWR/YLJoCqK1damP5o8qgHdqkc56biVpxhng/3Y5i67aCZPS0CnVz7p7v3qI
HqdI6SPFWrEJzSHxP1gO9R4WIbQ+WJ/h4WO85/e4i7VrPqpvT5KsMd3Ed2mjWmvaPNtkmQ/VRqlj
YiL6oWhE6lUqXATqoccU0qty/s0QtaI2gp9OuKkh5riUQ9levELkTmzLcEMebw8vwhB3tAp+679e
9MkHgcp8ty5lgMgzJKInYo85/DJUZXoKyZ6iNAYTFwoGKVdnmg8dwCsFLl7pAJD+h/aeTgE3ytkc
8ThaN6O5Kgnu/PlXbzoMqwO4EHcRHZPHq1Iv8h/5UHIPrS8L8DkmV1Xs2RO4bUex+O+kBqMyIsY8
j3KfoEYAbkJjHKuMdag8yvs6ZGU9de7znRipSwnnKF66b8L3SGGxnnn0brxLAJXwEm9KhZwbONlW
yDB6QLLPkteWzjSs+AMYWdOxHMkxSAm1gIubxVe+CHpDgRkoXQ4U9V3hrupUZgBW480QQqxVCBv/
pPtD0NRmQVF6Lody/Rsch4/naU1OL5ywf3CBiJg+7y6IHWrUzsvhaKzjqXfaLSnQxqlgGT4ov1Jm
D8FuWcZlfYmzacSDayAAWz/v58guw/mi2By4oOXcoiL1VKJ3l2SXKMtC4cJZQges77QZ+1LAGd85
Y8fvt92CVsKXvfoQOAgD20bVVGzj5J9AXq2k2N6X1OSY7HpIMbcvune+GQy+n4OH/NS1y4FAQDik
Ni30gyOCymawEjJDYMtxZ8t8OvQvQyU5OGMyDRExc07fAhJCaTUn39B44ZVJUevkyivUM2XwKBh2
73dl2flFyeoMind1CqaU3plEM+L+LbmjvwOLOfVSu3y162qIpxaK2ya+mUC0p4aPMVz9B+pyvMpS
yXZ1F10QMPhsWGAaHPhicP/bwpaSa9Pu/TKLdE6SMRX1NLlR3lZQRmubY8u4WLc/f+0mRrBRrriP
LkQtkZQWEdpiDkWdamAFBon22YNC8QmsPiawSzKODswyt7ciMDHeyaHBFkd42/mQBUy7RnRU0i2p
0B2bP/CWxXDIIu9M3WT22yP9+lZTg5pK8ONgqIFCuGIB1DTcAJsDhJLi5EjbjOlefO1iKxGuGKB3
vOL6uhn+KkvT7vSa19v8pvMTS+t65PzQq3cjGqQ7FbYuS+AqbPtNmWU9/RLOVN6lTXoXvj+7y9tQ
uoO5MfU723iANtxwpJwjB5S3fo4yKgLwkwku89PO9CmtlJSXicJY4KlJgxZw02OvdrjHvteZxJ2G
/JmijAV9thsrxWYPeDolPmf8VEVNe6f0IuMxbj1VKiO1xWatbM+xmHRy2+4uH3LRYvbFkZKKbJ+h
ywHRToPnHW/ab/4a7L8U+k0NQCTUvjBHRPlzgtIru81YpXUK9tef30a6mPoai+/GOxo/JvElfGGC
25i0Qs27EmLgWnYjDowymOwYx10sjSsTIjgOXDZ3DWCo+9+0ov9M3hHiOqyj+Q5DqZwgQowmfECf
7QQqhvCPMUk2FruSFH/8bn6QtVCGjaB43GViwAhW/ZrJhMMghSl5CGF+TyRA2dzkybJil65LjsVZ
daP7frYPN/5/EnubkLGSiyTlvtgMeT+bCw5V1xTgwwixMUaWrM8xYeBfUZ1hv6YWZSh0rKeNRkUy
XSrH3D0yMvkfDeHO+SN1dbf1K9W6oJPQybClBiczuXfr8s1ClWvLjBk1nZVFtxff4+RQdFDTBfES
eXf9oMdODXalwhj+TeU5j/heutOnY2JnzmCTra1v63gYKu0BLpAid1vSzU3FF58Bi77POVDQcZ5Z
mXhSv2j7wC2lmG05NTfWmMkA5uG07CV5mZFjo316oBH1mvhfS1coD+1Iy8e6ubv//wSNrajJYYXt
eulBTusSAKfYyWCr0yLm8g//rJ6rIHonlc+lS15d2BKh7P9wJrXeDeqvSY6pVxfxktjZiiZx4/hE
mBKlCLFW19ZYUwgoUwHumCNf5qGS5ry1aZ9rYzZtvjkFpfDbnHSFKE1wpBC31nZexKPTS7lXgMjm
c0R/jQ5fYpyJzvIhwTZ5sr/MJW2ghE5nTgarMlR0A7mT/HnY1BGrfoEIMLM6dLyt6lpDnytccxwd
YOGEwKGSe7uiMmc7zB9Z2aNAJi97pBQlSOugXOqmb6N9FirBZsyKKfWkz+OYZQ413T2cgBtJ3o0Y
ucX1oMUfl3yYoot2arQ2YSbn8D38XJFB2myPkHKPh/9giBoR+4Ly4ugyK9NX1un8MhhUAe1sNzZx
5aulggVo0hne5yOpqhWX8CQn8LT5zfB0s1FkWzHRwVcgFUU/iHUrkRzu8q2RupvR6/3kvlV3gJAl
IbzF0Toh73IR9hslkQ9xfwexeEXDs4491rXZz6kaWSCDDt8Sb/XrBh3+xFcTXw3gA3xWvljRoe05
E3tydEgwHqz0gFSpKcAEgWJAQIEylpg1nu1DNXomptS6sO8F0Dt6zlch4FkVe8VeTp7jHAgOw9fr
hLiWLm2MEb3j+r2SM5trx4P/HLOd1Zvn2u+F4n4GM1G13Z8G8/1pPfY+OIk7W2cA6rD3Vh4JmyhM
964VY79YPNakSTPSjQ+qHfiIyO/vvGIqRfyOLhAT6cM4N9BXGvuHWG1PNO3oyYX31VwfCpypJfpi
4IvCLkcZD8oBPUiJ764vePTkze+8m4VecDpEgCu5upojlYiu46pggmAgSlsRmLrPkAazpIfVVuFO
2HfB0ofu8LxLVVMAWm1qF+NBiNS9BS6qMgzwZpgi7uvfi53ZKKOhSVR7wjry7fOkNGIcV3TtziQR
Y3PnOSImoHtNytIJ4DpAXC5/5iY/M8Vs54eUgpbINhf9tbaHbUJ4NsAfC5qfa4qcH0XcjsPmX/18
vLfKcNDoORNe4nSP+v3Vm9rcPI3slVoGR7By+JJB0ThcdDDLLVkp2SzM3JUtOVMWL7emfeGRhac9
rm22cKZU8sd0VWwMctVUxMi8g2OqeHZJucrtHldWkUHJt7mqFV+tGfcSKfC2nd8COy9OMIHVxbSn
N7pgfTODM8Yv2hVn/VXfYo4D7/BenQIp+COqaXhTdYVA4QFSiiL7srtMlhgwndmUpyBxFzjhUEfi
0u3xZMaWAbq9Lf/85pIFRA0+arbLaz0n+0qkvuamQMD4mJsx0LdTmfTCK+d+N9sgHbdakhj5yBLv
ETK7rQZLs4Wd+TuCgnKm2VbCaKMH9MbS3bA1xoW/1Mc81mD7qhJh/SDPfFyUXlmSQ0vj4sUrKgz9
E+3t5/UTck2rT3puHZVn88FzRUbPlMgosNA86yuLjNHduT4f+oenVvOMZQSGxMN3kni/FiByi8g/
oBy2IQf8xWCJ+vvCtOHm4txIdkeM5BKKUy6IlWznq2YQ1BGRFC0vA7eJIJPKOaPiUQPgvN50Yw89
Ee3ePfe9yhQgWtOxOI91Bkd39kIDN8I3P7EbtOTBjnHIj9oWXkMJq8JDqaE1XCrMuSFV/7GL9tYl
Rl3JUJHhL2upX3Fa2eQHqweM5XCBKNgv4ZtYQi9n22j2Ox/kqo7Zj97gDk6O6/+ESC7jy/CztfZl
lZCbxhO4toPzOYcjqTSr1q9/3K5H586CFM2BjIdcKZ8WWg4GECTxNGrxK2cX3M5oNHtn3m7vWCmZ
HOmIWANz0XVI6BG9woeBxQfwEjAuOa6UrL4GGQsL7o/GfEuykTIj59ob1DMHeRomULV5YBlcTxFm
zb7Ehp8XnCqlKnRXl52VtQmqFyGGrnBEuDmIHgBWukAfwH3OPwGrZlAQl3QcGGPUU/gneWpOwnM1
yuVaVUZ8eL/NzmTEW9VnW+DfQa8gt0yTanNXvIVXRqjja4t6DX3ymHKO5d2TCqP85F6kYLDT1lWQ
Sjo0mmDhRpdU2S+9nmbqtk3+VvTzPIpgu89RZPtVQTjx13zQZe4LW9/c3N9NYjZmfrUhfSfL8Ugv
Zp7UaEXPnnMseCm8nqgYTI57QeWVCB91kUM6yVg0ibpLAsGM45NtHc0svrhF8ehnIxiw4t1Tjaw4
7hahg8giKd77K6WT3KvHLF7984sJc6OdICu2tBbEgVccn1dg3OOfevk7e8MwNX0jcpRS4ewjryaV
tzdgPPfvOB7xAh4ZXOBQI060jg5mjnd3moB/iaHZqtQHD6R5lsuvG5iOE+NCXwhgfn0TnIn6sd40
1Ay2ZgIDJzZbIWOXdvI8biIVa08zrTq2l7XLPAC/pGn9nf76g/Vtfid2T//hcMHLTdJGnPTGhkw3
9+5ZPdFrLtzsmrxPhFeA8qVgcNbsIKHB9Nx+kGYTlH0CfeF2OuAz8M0J17Wv/P0npn5Ak/CYNnZG
pgGnOHU6nh5y1ElwY4cAtCDPIRnQ9x0WcHutiuPuTz+gzVGdJQZHHCzBT9h+58cDozKDamxyXB63
Ze9MYbslthISluQONmfFFLGjuDbB3eMcd0AFfcXQtDsZwQMBOGFEBQlax+xxIs9zN79UpRLEyBmk
8CJ/E4Z9no+8iYiy8zxYKGRk2ib3uUOJGkDivZWdclZPP4xvvGx9C5UhHlTE9wvin50/KPDe3dlQ
CWEwuVmuyaNR7LMUDiy+RMFW3zN6wKDz6NYil9FreQkgvKZCwVmswEIc/MAhZt40TjqKc+hmbaZn
qmJYjQzya12mHKNsbCTqdZb0+E/xSf3/+vWpp3iz/r/kB+1l0dfvuE/D8reVWmgzJaDO5KLmS+SN
1AzV8cWBJBlRNB3K5Z2D6sR5G5+9gdOKpoA+vXXaAg9PNpFyiXypUoa6PxSIIT2z3CJTgFSa0qSa
mjQyLOMpeFRtp3NKB5/JqGXEzv73YUHbSBGZLl//jqgVxEfwDKGP0JakAtzh6yI1VALeA8S5Eb4S
7b39+35Ca31BGFt/ZR5dVyrYcyK0hChypWaY1F07X9Bcfzz60DS5PMeHTjnGuemd31bJGEwA7YWY
DMx8zaz2yPzCb6KGNcYpeYCmvTcj95W5AaCV0jvGbBBGjZ+ebYNOdOc6K+R3qSb+AwjQnhIfTNaW
a33GFcKNm1bVTbzEjN1V/cxrwCEd31C33Eksn1tytqzJEtKA7uk5DqFBHyBvtwl2miS8n/ubjodL
1Ujmya9kuSadhdmJFe8DuHBjJ3mVDr5WpGQvCee+6Y45b+pQmGc3yKX8F0f6X1drGWrs/auidllt
nuWXCHYuVcgdYgSBGauoxWusNOESWgRjI0Dx+gWhlUgdEsRSRGkFoXEY2K17zHWpK24X03CYt9EU
oDilU3db6OLE6101hVVtHzuAQ7zAkHQPD8kgu/POJacJ2wnRPv3vDLRwB/VTxfyr9oNi5YNSuvNG
WEyVXfcJR0EXCxu9qza6LHJnMcFrHyHSyurdpxj+W+3ZMRXd/4LQ4FOtt64WhhFscNtT4ZYMeKOJ
gLgWm8TpUycY8LhrEpgx+MvZxTsB+8fZhYL2ZzWqdPWKZWqaf+ZNsv7Cpca4oiEhzStnz+WO7YDo
ro+k0pajVa0v0wUcHJZmBnphjJAzPGQ+YeDrcbBXkDZpWNdjFTaxktzpZODXAnte5E54ENhbx92H
8kZ05hamRvi/qvY2926MhTqi1Q0M3tNiuhHPZrL+9CoZxfM8p70G0qS1h4eFNc8MXuy7wLAfwp1E
LMyW+2GE/CHwzaqKGstHRSQqOKndNP+7mYJ7rIff8IMelsWnFLv2ZRs6cM2YEvt2mOoQI4hD0K5D
2FqITjfkF9bU+dGBPHQG0lBzvMZoSfjZVyedxhJH4cHmrM64p4LzDtjkhkq6XR3fwghosvh9XjhJ
hTuPRn51tUE2UhFtevpqBOiOe+i3c9de9fFhVddOaHsPMuRlctFEXuh5ZK4GFUsMZu/CSXZGr4Lk
jHtto6ZMmR9hmDfq9QJnix9hdZmVsXYJUxXWpkTrCHDDAbk8WMUQcKzGOZQJ/m4h407z/MmVmSu3
dDa6SxKtK/t3AQJhC4lHFi7hDE5qHVxa1X6uUrsi+SVQzu+S1OrZAPBchmUFbRQjn7jb/vUS2KVG
gBwGSEXm4MqHFh3+ksD/0UuyhMW5P7990MRsLd7dp5XcZKG+ZPe1YhDpS66eFu2YFC+DLSl1nL08
I4Uk8JFmSiVnd/Pg22I9Rm4ikxES1h2CXVt59u/YhMJI8dgEnjcZgSOUxKP6gdtC59pgq/XboI8A
33qlfTtqLc6kuKThyVexsluX94v5/6dga/QA6oIVnTDlUh/4rG0z/vTJjmtFanr2BWLwRIj8oVRA
u9dM/bpHPkym7Qji6xK+WwOEtpWRZrH2pkJGL4NQ+qJSkVkZRiV6FEPC0Bl4xX16jr/qXJXNGt3D
M04lsP96UWxp57Evl/8OoZwdDuRZT0M7mdO4VLyusTbnlIP3yQt4PNsADPhX1uXh1FPBVjQgJ0B3
nJzbW5tctKeSSmF0F5/mA5UQD9ZmW48zozNjkeYFeSB17UBayr1eoYGhAXa/lqCdaUkzNOwqNd6z
T74kt5kAOSg/KMv9P7SqscakLch5X1y6ESLnVlqr3dkPbKIslp79lm6s+W20b7cmxG9i8Btna9h6
vxKuD+N6WxTQYafdNCxytVQbbJkiJ4hx0iuUBdj9Ca/mNGyqz/va3YjP7XlDiQru4Z4OgfM7Oygz
RNjj8muL0/+lRaG8g68O+Ou2kLKfg/8PfmO+rxcjvSVagBOlAgNk5rmcEQ266rThsjzLaE/xnF9k
G7560qKZKzLcY2nNgkhCgnw5E31fbDKBv1lsAIVoW9nI9E7wZdCXEaefGVSU2vCH0adZFS4TQv2x
283Yw+zPgGlxR/+5thrDrJ/GSe/Da0prX4NoytRS1sxuIM32i+ecXgV+l/mlJwmDz29HYt1oA5YO
KnfntXx80pwhK6I+l5ANlF06SQYOdVSc7XEztQ32ZYDkX6sFAoIyEwE4YSUWUhxXU7759631jYE4
C9S6uyVfbbmvWqz0hY+/9LblA8x3QmebOfja+Pniewn/t/Zjdi6cLOuiMzDebDlt/Zqd2DkwHy+D
OZAtlH4m+bdDseI0P6hD5/edz33gzpPEyAx/0rOh+0tsucZBdgwpwXvNaLEUHvXKaEvqBLK8vT/4
sjivUJntpmAXWcowdjbbNNkYgUOGhjM6b2644aez2TWSdKjC4WKk0+F18gybKPkDydDKIsT1bkD5
twq009Lic4vIRLC3/hHmvfotvJiZjyMKt53Ypl1tyE5UarOHggyhEZ7jo5PoYsAPOim8bCF+XIyN
D+my1rxawPFWteB5suF2oZoI0iTfE7qGeRZVoZ8Qx7PfkBcEO6GxEXR4HoNPcBiueAJ78E3tSC6n
ms5VoAgVzljI9i8Oygwa74fOqiUbY7vvmB0yIpqp9HI/4q/Gt60FFLJ8W2VqgRraBk2Axw8lmKLW
2l8WbIByKdEDOPDPT8vDmbIeciVlvhL0vbArVvDGUzp31hk8mcU1EjcnXLvuIT0gKyjjE5pZuLg0
pBp7/HTW0qeJfwSE10VF1G4HwfJjMQ8xw3+cooETAl34h/qg3ucITnYhn8suZWwmz6f2doefD4l6
cvgAT9kWX95u1oj1FRGQO+/VWStfRx7ioJY6XRhq336k6ikkWwc6GaCDinxiZ1pRcU/Sh1B1Ju02
h/bNXrWU8awdNDDl9HcOj8G86GqBeDZlvap6BOEfbzL2VuF3xfrwtwt+/6NpMkUyAwJhVRaHvFuW
ZWugGzYOU0CuaNdOEiOy6mEX6SzEKmaSpor6czvzfRBoYkrL7yorL8OgzC/Khcyb7aDxBmXOmP9y
9WM7NQxMvfxnJktZLEZLuuvVqK4KaoP9wu2oAnQKIWRlEFQhvPQxfML64psDnPLPsDpNDzKSzYWN
ghVo580v7GqiqSV0V0zrYEBG68XcnOniob6Fm+ipMxoAucRDk/SD+rauNvG2hJnYqQqr+c/+ohFu
wsyL/IKAkUv8jKWkWkLYxzi0LJytpEUgbqxdqp1t6Ah+y8c3DOIMrvIiT0SXh5nmH6YB/GVSOeC4
Fe8sbkoidqPtUWBs3EKHGnkoMYXFwLmEB4g8K+y6AGbo1Q7/ULU8OLqS63tnIH8kBJKzCqj4RWDC
eC2+mS+b0kzK1PTAqXF9oOPeWgIKz8tglm9deV1u8ZttqJRmVHnq3OcB6pjyiUmmxqh9+MyFpHYR
0+Bw8+EmPYWpP/I3+r5EOJvGM0WijdTqooXrJ9I9yx9NAbXvlHWfcIWW1oG3+wegn/P9RRAoWODK
zbpFIR1xo6F9YeIqE5zPpkO/ZUf2l0rNY0wv/DY+co/kglwVsYR0Ygzm66P0BB468AmJ6qS/OKTu
4SSPFeHLJwDan5o3fjzc4AH7PhAVeL7vNvLliDmQz1eqcIOOyL6G6fEVlaaOtJChjTFCf4O2nnOy
UyixdKcNmt76+6CsCfrrBtLILmuLCXt/arUBY7n6T1ej4V4ugKicLqx7uZ6Lhxbi+pdCOmvXjn6I
VOwmqgPxHdo7nuIvHxOrU9DKQinvFTk9ECOEBum6fpg52cZhKwHxy8obhiEUI1o7cSWqCgQckMdj
jwts+0Sjt+wdfPIiqLma6Ik9G32+SSXvCML18J+d2e235a+Wt3oHcelnX4Za5rRIZOHZBmVXRb3S
vFVSO7c+TYVD90+MQy5eCRMW9SzXP4lw3s4sT7Z6eUTmlu6nzt211tPdjFnbozIzQFqo4koGQv/X
Rqer21Suus62SR9e75wqt2jyQoICRXV9AlnxwDBPbdexWA4NbbhAGOBOBXxRVkuJQfR4GI2Xr3TK
Ho1ZV4O2knSKqhXVmpxvk1dg6pWjXrZxI1Aef1woSCRlPP0JeCSl7vNOyGxwe3fFrsCZmNZ79ozO
d7abOkg7QbsOAR/RLKFUIcLUGHWDoPE+Gvz+fPdN94MBtuX4av+SHDt8SQUVK1gTfzYP+uLuzP68
cVOiY/3T9yib7adY3HGl/6u0ArusgVvNPQOnGtgTNu2ZbzgmHWJYWb47IfxRu63nfhH86QAR2PzY
kVuI9fuyFUBcAelInxng05LauwMVv/DxMb9Zow5dwiC3cN5DMdoJf2SaEvKQM/CBBT/bCcYhHUgy
Bqbk3ybflmx6plHBrdt3PLRlNE6rePHeBHx4jjIjLW7CG3uLylvq4pts70aOKmyucOOEWXh+bdra
2MpHNj0JzF6bgEMdYTTuP6IXtfnxdPjfAsqMDgzohhdGpVH4O8op7D8y1C7WxNNgJvtV4dSSYYle
LHFAXvuJCTdUPrFTmMe17hoM5KsmOJyyNqb7NZ3AWDkU8C2aW6MnC6PNovsarKCeedaVNWg2/nyf
z4kGBnusoa1n9VUsP204N5HBbJ4jvHvjyPZRFAjJGsrojrUwD30RBqi+DPHILj5DVsflm9No9/4G
j8PzHlXD6Sj/cXpds13mhoAGXl3pMiic0SjYVSU5WgPqZ4xxydXj+4LZeLrRESHDuEFe4IYnIp2k
1zKlo/hehrts8mbggwZfOn2EJ0L5lk4li8I0INhT4geZcdM6g5Jx/AZkaa8W8746Gjo3HEGI6UtS
r8f4jUhrmKh/fcL9PSOukTrJ6I1XMZEEZPRSGSdT/zBFilJz1IljEjJAQ2jg3znrc+a1nE1dhQJf
+lD4d38Kk//L1ZN770DwPALI1dhCcV7W4uxQGi/SWFxrOscIeXmx31rqcssHyqBrjD1EJWIEV5+Q
/2K/FGONYSg/HXRmFCCMH8SUq2lvt2Y7Q2sH70igdngwo29yFzp56uMG8paN/AMZuVfwMUrY9cB7
uREFI2fw6Aegi5odeU2PVdADZaLg6DbzStI4kL6iVGN1iU5Dak+fAYS9mpckxyYrTsbpx6hT8GEA
Grws3J+F8157vN5GQZ8tMduBpLN8eNZraDsfoB+FuD39CDySR2dK7UrQv2S7OdkJBxp9ecrl5D82
NBTTItwoCjBYB61wWHNAH+aaoNZrNqez2u+m3155xboYIYcpXHSluDeMhXyWkKMho6zvNYwmdcnb
8IncQDDzQBUeh9I5YNlUDhDmHTrZ3d1Csp9ENeRGTgoZLtmYYLBRvePk7hKAp5l2C7f94j5An3XP
7weg1umoH20FxsncO+JKh7IXzpPEChHVx5f9TbBMJt4XR9hwBCZS3KxPvvkcn8yg2Vnh/X8ekfUn
4RnJOJUZhnzse/QgLdgaTUaNY9XMiNPoFX2vCWwHPZIRWRqLjLaOS7UoQwV85VurLyFIwK9dSHd2
IwYshGXAb0coasSUlPn5gm9sK7bNh1HzrB7HUvFCKCxKZuLie3wpd/zQy11Jgh1JJwv8j2XFo5I/
fmc6tN0YNrBLosvN+TeKdUkrCORq9Ce/26BzmUM+h+vuZNZSl9t80Q8vseYDG8rmWfnPoK+pq5dF
8BcvdvV3bLqRD6IRq+sSowLju6ftybZ+Umm2qgaHVLG4VWZii72sX2djlTfY/m3+8WxPHVzQngUE
lKI3/RNZHSdSdxWvqGBWddQtRI/AU79dQIDYYkj+jlqMaRxacLVDiaI7jgQQMjSJwnuU/hV45Dtx
zjkLlGqCTF3orDIq422ywHM1cL3mxzNJ3pjBnKXySve8Me8HDXBbTmspAMfoDMUBh1HHebiXWWM/
sL02jtkAAQGWgGKueHQXFOet9eC5cHaiXeiXK4oSQ18GCOtKTElAeELmLpPqkmNpcYkMDyblKKKB
CQ7kb6t4erY3XIJEPm/+ifkkfUB4U8L0JmX6xwRg1eJ+22m48B3ElviAHao6Ze9I9mUl65qJyXqP
aS2yv0o6nhpcTaq3yL+kKjBC7QbBr7MuWt/qC+mCi74gweJt78QBDKKYPLncMPKxO+1G23+1Q340
s16vUvKXGT/ZI1JOErXpCAL1s4nOOriPYwzOTBKVyNTSB8SrWfVT+Os8ysArWEwVwUh9/eUTakBE
1OWu16thMl20lEdMwb5t8+KI3lRjKt6MCReaP7AhSD9pVN4E41mVB9065+r5MBhXgd6Lvi6FcZRp
t1p157jtpqaWH1BxyUuRL6D1Wd7nvoz2WClYDg4BM37J+GkpD08k7vO/lVISF7gZ/Ftj3Lmpvpo/
N4HoVoxrS0EUWpolEYWQT5N09DkNj/pKo31guXrQOEoBrD5eAjvsdC3jFCK+onIWwa043X77YPdf
xxqYgxT3tRomLML+ehtRs3ePUolcsarbl9Fq5slmZh8fnLW/Ojl57F+golATk9nLunHhxYbYoaSe
gsmrfbiZusLVF1Qfdie0DzOQ1HlPnJc6BTBy2QQtagPjE0J331yrKHQxvSdKnfVbhT9VQJnPaHVo
FX5jMBmnzBrqtdAcxuw35qT6FqWbYIvLsp53n/4H5l2IAm2JIr7r9+RCbVTMBenOcAaqgD7lGWx6
LfV/w08XKdgq5W1Gk/fgNjY4zq89R5csao/XuNrV8QAds910wMaW4kzuMxJDRKKFYRep5Ju0ziEp
aY6HstWTXbqIyBHDtXSqpnzytF/8USfIZNNlSxqXabV1IAomu3O4RDCuST0SAHiRrOz1khJN3LBr
azNfg+0CdmDRR7rRCaeGypztfKTqUCSZCUF0IHTvU09o4eEE8KcpiNwUHDzgVu2T7XerGMKf50ga
ya/JAii7gRoupF4xQgpztUxTC9BgOujfRE4GHUtxxgiHmgB8Js4lkvJEg4nwufEkzidSje0gyF8U
pNziGpC2Qpn8DcDmdmT7NuEYr1FKP7NVKfA5caX1rF8AuWsdUfPT24b/+7toPfn0iFhB5GmUDtUm
0U0O+aIfD+9iVBQj5jDW+DL5QLlHrZLMB6A6vCFrzNEoPXVrngpX3ACAJG5TMRl/u62y/0z2EoAC
FmQGsafYER6Qqy3ulv1ROH0K93P3Uk8x8hP8jUCTuHTgJuhUfEvr3kRogkfz87lt2Nt58AzXwtGG
W+Cj421jCmPIIgKpm0lguB1EOckPBTo3q1EGf0tQvOUqiaNv5ggu/ptjketzyf4IE16/xPxYDAxM
sAEandx0M5C4UGNsFzd8hxueVYOw+fHZYojqetgGZW1bc7I1+C9D249hIAJ28k5wnk4cvjeOV7oB
Hr1+TaK9c+B1BxFJVXFpf/358Vzdl6oGsEiM1zCPakx1pGwF81k9h9ohBmYHNcfihFpye6AJZ2wg
T0Dfb4/SQ9vIrHzCJgni165ZBx5lZ4/DARiCuiP5Encv8SDEf7Blogt8j0HK9/lA63JnCfniM5pI
nVsCWLUqyeV8U0gqLd3E9n5UygRkqWDrDXFLkRaBglnrAgFQ+HHXxYqVB0mnvkR2BXM7GqbHF4bn
UqWuuMkSOlwTmuA4qG3vjXcQVIq8WFzUpWePw4mmEexQVab0QR0Ugi1YpQNj5RGrgc8+ienfSw83
QlKMaPVepIT+A+z2vxmJ21sQrJOA+s8P5Af4O91wvWQLyGSuiNF5xiELNs8nHbup3WbHyyel5Wzr
5YF1C/PbbSfDvxoYx7lJBGlkXyjOzth8A49xdf+RUjo77mAuQuVovOPWYTJqUwZybJEdxu0+6j8n
wt8YkzbSray6GwD7zdvQY8NRrF5nfloYZNpHPsn11oDQNWnYngUYYL5EarUBMgqojXENQYWmcW1/
WoCXv+uTXHa4fl3vyiJZIiBlU1sLK4aKdJkd5byTYRBtyAaeGGnMnReUnrPOj8/H4J9Kfv+DmZNS
jmw2hbwmZsZLAiLdkTSW/D5mzU4Jwn02kpZAnMgAPd1eP8wRj1Bq17ebIq3M4pBAU9bSBTXA89It
0b+gxDZQm2sQlT1hD/MQYKKbDbTTjmaWjOy+9e12sUS+ezKSBRjYWt+vKzgKtxlVQfrsqAPUO8Oz
EDBLHncBAfYEeDkWsHOc9EozbMLVfG01PHhg7PZe0eSENya7usNyGbtvHK7IMB0vqrLd11itBi7V
ygU+lFNIh20fYdINOVsxPcyyxrxlc5efyDeDQe7NmOE+RrxpHLR3oKUO9uMwBkTwrNocS2ek4VYI
Qug1u+Nt6Zw+XTbaTov2ZEBHcdxXFWbFO5f1EDlKsVZkPgmJ8xoWIw0HeYFHa3Y7pDfY2jh2CqeM
C2ZC8yNXzeayAL6kGFuyeplXdIEU5K21KDW561xMDcHaA9WkazmgRj+20PufypdPKJ2mG0Ot0Zkk
+FW4UzW7dgiNaqNMpx0CY3UL7z0qWmhw5FXHPt3TbqKyOi2tWKORucWof+mjlIZIEDLN7RtQ2k8W
K+MCUq+OTZ/P8eLnzgwp8BUwyT5yG85UKH2ISTpKWUVP7EDy9xGzdZo1Xps2NTGsxTSDjZjjez/0
yup0mcjVJLo/Im4GHe8nn+w2kYNJmBZya0DDYkLlM2gh1fJw5Bs+SxgUIDusmujLSRihaNrY9oxu
RWJSVKifNjAsJk9ELZXyfuP3hZZWpvpHObiQ35H5lfkdr1f+cet5W4rutRAnsOVP6S5e4ESA0l/u
8fKvoaoQfZ2JGEs4iCL7YoO9XIIhq9lesqsdSBvwbEXB5TAr3tGYZ2ypyQPeH9FjzZCPwTDtbQsG
61EO2cqw8Ht0NN0rggZnAjrOUcRVStFAEU4jNYE+Qj/tBqpaBM45sMEcrW4Rd7yeX/PrwcplKsS9
DFacyQjikOvWYXBIBHzJR272/CqdwI2jzNOSFy8mvPC9SlKDGfRork53iiw1nu2jlsZVGZQvb/JP
KeTs4b+RP+dkZUvz0N1TUvYZ9OpuPyYpMVRWTHD788eCsUcuScy8Jvr7VdjcDvzjdb8KmLGLdXug
qSbKr5bxuAZebFD0BEbQMP7UryPYw1qGPD51XiRZ2nE1SJkf//F9BC25EiMHbVAcGy9k7xrmROI+
VHAmkFCPgERLHki/kHwT1UnpxvpGvmxio8CHjv/fGZ6/BA3qIOWa22OalVIdXAFkvS6y7MQE3YLx
VFalR1l+hSy5q3pIcZAWwBcKva6FMXG1cIEvnsJhKCsNT5zna6wnv1r5FtIALr0ejO5AEtPwgyCv
VReFvRDL87Dq8nx0mQbTx4wAGYhKgBxks2NMW14m6l1FoKbIdAH5QRMDp7zy/H3ijJCBpAr+MCdp
nuHGzAW6ufpRKgHr5LYFCxPf9+tB1zoJbLQRi4pj6ndP2LTtMOvNcrBzf0Y6ZScpX1fq4ffr+ax1
N0fyMQ9kmelBW0ol764yHfhcIscyukhYtz3GHpCr8/bGVS2MO5jOY98yTaxzUVU9GpfBSdgq1w/N
Xag7G6V2aCGmzdc4awnz0CtkTN0swTWSZ27sZTA7Y8NqiZ9JSA6IxljzbUjzRT1iEqWBQfDKP4u2
wsUHet1VPz7VCkPemzH73rBu3mEeC40iuDrtKGWG01fYaBQjjR78c6dn6bBfP93cMVIGtnCE/YtA
eZOQFkqIMcq+me7FyeTedpajcaxaGpQxb1fIifLBnVFJIpCmuWtN3fuZZmTnLfZDGubbfbzIXn3M
ypQgARin830Z6nA9H1JzpNf5ggw57eFiwR4Av21yMueSGms4CRG1xM0h0OHGopl647atoeZeMcdo
N/RD8NFhe0PECBxhXSNppMon4pVwW0JTmjR62QsVW/RkwD1dQJ6DBILoTLIckVw9mzUlB0sslwWS
VrxtxWynpmo38y9cqtvaCumHZNYE6Jhl23pzHZrvn/AtkDy3T9zgkaDUWrJECQDgStU3tep46HY7
y/OGhqw7u8+3/tNhiG9lEFaIwLgIxfeRSvwllXzgr0cRcunnVLSRiZd9PTHlkyHtJi81X1WeESoM
+mnMYVtEp34U5fctomJnm9epDg4OXC7GKDZF7oMGpW7mch5yq9LxYOXfid8ZmvNYroe5+XkIfHGp
NAORMBEVwpEdbmFEP3u7gYQFvdtcxLkFN1ZttOLOjBtja2mH1rPqvWakagI4KOx1VpegUVirN3J3
clTpJXNZ+AszOidf2SqPAKthHEyhy0Nq6RZksHQqcOeZsispD/8ZbJ9ET5BG5695AqDzkz23wRwu
OOJqFjJBodJxQObDA9Hy95qQOO550Zz0SgXSNsS4+Ubg5GFQg+wyUyu6cDYAFiO/auV2orKTLDyM
dllP16b5E5LM3tf400c0r93/N/YymY0op/sNYx18sTngb62N4+hfQBmfo2XjtCDsgfBOcpAR7Mln
uUbl+AH4dNdTPpAly783/7LE0CVVfy+l2//poUFgNs3KYhab/EX4ZlW0dseQcMlKp+r0xTV4Q6d5
oB5pj86pXnM20+P+Zu2YOUe1luPuJtzyr87P4ZYi+f7GS7ErTR2f8G8kJIaxIO/tBGVHXpcaSYs3
td9r9xEYEAXk7nhMyss7clpP8vNAOtIscwZBBZMul3S+WozafYcmtfEoPNN+9HZulJX0uqmISdLQ
v0Qu7uIsaB1Sn+0BU6JP6JappG36ILxTJHzfOctXrwEgdIl6Q5GKIudxyYwK0mcf6x+rPG024iKb
/Ygfls5rBIzWfVEWPHgGKtSEPNVNRO+coGZB5oQZfCEtcoRPO38x4dHbtxw1F+jmOxLbqOSC4ojm
96oIIN1KtbZleJAZIVgpzyxesqGn8uZJp7/+BEzteG0EMDslGMLWPFHTnhuSHgYUdBJeHzw5gh4J
y3jw+l19/UjzDuJH8SE7g4DOZLd240NCyS+t8Zqk4dlbbxNb3YqRziHPm2Wf22kTz0Ux14xaTeGb
YRlXPpZ+67gL33FDoi84aGYsHtxawXjDnEch2FucV3zsAR97O/rzjSBND5uP5Z5srgHrW/gtTbkq
eSyAaikSkUXcbANCsGtlD4ui706QjxuayCmttMlPctvoqgT83RCjs5RJwnjc3pEYEWzVIDQiBHQO
l1U9SXCOe+Iz06wcL84NAapuUztrsezhHpig/nGNjenpWp3ScQb2G1QNMOLjvsdeq4cLPwMc/lbx
eMulIgZuwJbXi4hxn/Aw0BBZa8tqnAt7svbDKg++ECK6nQ3VLbuvTJzJ1ql9T6Xj+SZIiGW8Ipw8
M8vEYYlHU4Iu+ossSO/LOitFO8elOsgZfLpRO9Y+ifjEOugjPo/tRF5RrTXtHiTXDkqOWQ3tsCAE
K6c7IHQ8GDLr3uOlSH0WXRDMGRQ7tF71cqTpMTqL4dsVkFVQqdZvoMFAt0iR/CpuaC5Y/jcf4Qss
FKfkx0ZIJdPqllBVBCwd8iihx7roD5zh/AyRNbyAXpO019Giagbz/YikFLd/vA3pFo4Jtyccr3Qk
htU/FkDJJ0/HmUkuDCIvxLVf9WAua8xyW9A9gBmVSyPyX3+xK3ew+xi7V06423/8eyDkPnFpGz46
3VV+WSZqR2YWAmhNIacGmFmjDLCYw/WsVAcbOXZjn33um8bPvUn8wT/4W5TssVtJCu8Qs0ZF1mR2
UGxmbQ+ab4wKjYQmoH22Ynu/8F2HOPXrS7bef6EqqK2Wf5v55Tww9F+yXNY5iX5TLXrOjokVXFsl
xOHFvICvMcgiHc29nKjGuaEEuMpdpOuXXqhiHLKz2d+mhF8eaAOUaPMiPcIHpyOZyw1EckKrGp5q
1qTLngVranUfMg2mDLFETExBKXPHABHAJg0Y410KG8nJa98jL7faJz5JRGGGW9T8qofHTdmV6fcz
6ajuaELRHhSlqPEsAAjSJkbjYGihLBGMhlgLRELWAIG2ryhtxZ0G3+62Xi3e7WYFeMQNQ8qOhSpj
6UZSCqjm5FJ+pZL3OeyfxlgMQs931jtDNNI/8btUVecKRjL5tnQGPkqw8wYM3YZ4/Pa5kH/0D7s7
sU1mAhj+xH0advE2j+l+Ez4nozKDSfWID5Bk26hPRGeHwA+MG3VhYEKeJzqbHlFm08djxv/8fJN6
IYvDfEbLWsX2rGJS0CLlFGUjgKmb/nNxabTzRL6EL7TqyzjN22N6vJAyG4HrOxQurY0rMtPpbvuK
mM2Q0sr6vOOVwp9Vw+mWjlBrdnJ9lsCCQPTlcH1/d3FO13kxorHoi2jbIFLyVrGfJi+oXTyXgmMK
L4vlqgZuATp1rimx3bjn3T1FDlckp2GdlLxQ8GiVQ+wzf1XCc3tfg1p4BgrNS9C4n0m8l3Px6rZm
ksYtrfOTgwcMv+ad53KTnFKJKceWS2m/FmLEobqwz9rJBvgEgvOUcXoa8HHuS+PDO4RUFJmgQO2c
CBN8dPbnJY3b1+jMb8FOaPQlzEfmimbyapX+pOgO5viXGkwLjGIMCcSEnOMs2qcpXst2X0NR4y38
i6wKFAc7jLSqLtW/sUDx5edyhHDvrcSu+bXnHfjIpli9Q+iLUGPHjGLEy6xMycqXODMRyqk2cLcG
uVU8RSA0ZRarX1/eycNpb6tz7H7TU8ybXO0wKy3mRR/WiKpQGlhtYDuWcEiZvZX7xj+rA2Y9f/TL
PcYZFFWc4IdBxCJnznrhymxvpkjRyx+4r1aDwC1CG6sVKoyNhXidrW9AxaOvZlXug7lXp8webg8o
up+8l0N6uTdmLOdaqtuU+fiyOt8n57jczYRun87QhhNfiQ4WToozvuPE+E5QKm7wP4e+fZF4cr5j
oODBtKVpmRvsTGjnUbd3ZfTEI9LJOd6Mre56ELJKWESoqsoobVb9mDLN8dBR8GWGgPZXkhdP2pb6
EQ7kxiYtOczWY5DtnDQ9gelha5xiS7S4o7YD9TVK90jSXTPpjihaqtIzeJLT176nftRZQxqKq4Tf
x46FU99ZDnYKSsFr83Pnhz25uqI5yn6Rsm6rrtpxM4aWUv5eTfPtOJ/JCtecVf2Ox7w9rz4CbqwC
1gAuJLQLAaVijl99805WkXQUq3gAsFcke7FZgXHRiE7lGfurysGmjpLZ7rjuilDzmWAzuPnksiHt
VxK0I+JY8W4t0qHNTTfkJixf86XJnlmrLl4UDFasZ+8/ocsTCdS3t73BBRLXTakptKvyUP1ipZc0
bmCjJNUSEXSzynVxcdWrikZBFOqHeWoWDQw0Mx5d2t1n7CPWxgUcKBBWnJ+GcI7LBLwZNdM3YhDo
de/2mY+uyrpE+Wqb6nxASyd4C/y68br9i8DuhMhKu+LOK1J0IowO9WwEJV/Avry/Kde7tQCHACGb
horehUbl5fb4xjWiK9rrEiFkFhXNRs5DWzvBj9q43VOvQxu9X/fOHZh8THrnuT5MvawuycBA/lVE
zdTiHdP72EHxnnpgLqnWwaHpZO3JTpC+g+TiuZ8dMwTavRLl461RcPkrmhI6nmVggUkHMivDhfQ5
bKPFQt0ithx4JMiPZeefTsdSbf3/V5AwwyO/uwFm5szpXfNXqfEHVI4XZa6HMkfwb/H6waqdOoGy
pMHs7XKQY3sMO7Bettw3bvlPGVt4Y7gWqUfjJqr6EUtHp5xuPcGDXWU4jp3xC6FVkOQKMIJnvkHf
FKzastJLaKOAS2pBV+i9uTRI2Ld5btUCncm67px3N6JXeydKxxjHYYGzuPNzY9vLSKDVHMBVbAV3
qnYTRY6u8rd03iIOZR5A8Koysnyhii0lTzsuPmLy4alXI6KBhYeO/cVeyUGECPO3XLL6kZ2o7lsf
vLZVJtevT6FRQqFuwFLPVpmkhpn3DgmzEURDWSXWNOCqUYpMifkPTs+ifvYnddP2mE+e/D6Zm7q4
yTJ2mXhC/zsC7cVGuusKp4Of7q210R+Ex02ADwk82MpoI1j3Bf206E5pRnVupHwbXW9J01jCSyq7
NIgsMeMnys0+ZkmcmTHtD7xyaFT8OBLQUNFJJo3QpyHIr1AlYNIpo85Wqi7p3n9316e7QMAy2guD
g1gX85iyJdi74xGVyATj7qpVHTPTnAp2vSoxEbqjIVyEy36CFUSmTzvxo/nh9bbo8mSreY56W0kh
P3OyuiyE54HiDYRxoqHT1Y5sGTOwTwne58Qy+88WZl5JpezNkft2oHt92ltxOcdNbWrERNQUcfzR
Z9x6B19VABf0eBbPd5E/YFc51iztnCfrXEIIGyeMgH3IGq6jZNPkbR/Zv91VxAgl4xacpeGhhEc1
DA5fhS9BCi41YlNIn5zQ3H10+SFvJZyGeiWScbvTSFBCMawa/Ha7Q/VVOrFJ2VpRAV0264Yarcyn
C/Jldw9L78G2QrAdmDn7nBPIkZR9m5hYlHWEDbFzVxScTmIQwC5/9gnmyC1OWpjFO82bU1n+GHYh
q/tzYr20Z/Umqd+VwICyyuh3ZB/MfWM2dyyb04YiN/XlPQHt3Ny0fkq7j4LofxUi2IytmFxMVrog
/f6Eu18Xyt74FUnc546R42zpB3v3oi+ErqCNs/o77dJHGYOsTQ8k/KfAC6BBvMeM838w4Ugn4fdK
/0YheSo7fwuOj0hwlnypfuN10TJZw6Qje5+aV8cCPSWYR826ER2I+HRE01plbyxxkdXndwfBmC/v
JMft8yvSZMWzo1U48L0xGWdwYoZZMpVsqSZjoQpHgFx24uLGe1IY5AgcnoKrVF7EIH3+CbCooUkd
l56QzF9qk3w460fJMbaf1boZUILjuNw48X7dSjqp5e8YjrTfIuZm6HgpXYiJEuQeoQJ1LzTOOW/V
B9srvdoFHMG1LCv5RkcsqNKDqq55e5z0XQ2HwA2z/4muTX8XPaw6fWluyiel7VGunui4PDHEptso
TQ4KttcMQKvxryqzcisbydzE/qeEVKEtx18o8TQnLgx5CAhtmGg+/+vu/eXHReR8ND3ki9Th4HyH
/aOQAelWHqPA1lyOpyYgHJeF7GR6fFPbxMQVdlxt9Y9SaiE8M8CiqCkVN1Mjrf7yV8TDGY1JfZ10
0nMqL5LZapsOPXb7JlyUofoko6dZK4pfgUPqojJfdudETlW2GTwd7HVkrlJ6QNBQoO2bwJl8UeG9
fdJH52X1vxqCEm7y4US9a8mWF3xPuB7L6kOfop79bQu7DapdUfFv4fZOGh1zRzS60J/gLrYxS/ha
hso7AqfIxkLS64RnrspJ1wTbQmBFl9yFPyCdASFP3u0g4R3iNGmzZjaZjTrxsNXDExzGNNbjMa5t
ng7aSEFOLwT9tZQ8GajIR3UaykyNQ5J7vECdcH28k7u6JRQqOfuoFl+LrWbvN+FJ6CwH310R0KkM
0RcioLDevENQ0iJS4Vr07v4Cyg9Sn9NcHQeMjCUiA7aICvI9wi2GVu4IyBLkfRnrp6MWOjnGZlqG
u2vwXTXpQGHoAmT5rwnHOWWXH5d8V/b2jZJwDgbsvf1R+kCsBT2gE2A8RSiAVSn8PXMmWABiwVhx
u51kydqbrX8Td5B0uk25EyZRTvRwYWzfnkl+IZrsWEKu/wceMD338V50IMdhvDwF7QQ+CPpKNLRG
f6a+GuhxwcFpleNNDOTAU+zK10Huj31lQ0mlw5GL50jtCVYEB1KY5Gv7Bu1de61wP7jjjUuMGKEm
2iuuNccD8WX4gYnMHxHLXYVD05QNsD3EML1zel9PPLa0hrPdFYy4w9kgusjHhwbNNibVmFcaksU6
RF+D7nigQ3cRVRHI4CuqG2u3bV6ZGlFAWKJmJ9LaQm3GMmPgBlO0UjiUbi9p9da2tnRTjeWJcZQF
QJYcAtI08Q36loOF+dShNGdjLezrtVF91LqF4yaBQJnLrhOWLChOmgwloZqeDn81P3krbp4S0BuZ
h87AsoBFMX5i1wTbGwqUZzMRZ/7ApbvqFCaEXlJVKal9M/bH5T69DSYkhos1coA6MORRGzemYY8X
Jryj51uxzxGvnxGpiIH5Ds5efQnTMqn1jJutwJ36qXfExHQNnGfUdbIEBFxFFtB9Bu2im1KTR02z
s5lQELqE7dRd1/w12FvJabgjeJmo8qODiAX+CilSxd4ez2qBCA1Agp1lP/jEaPALhcwfJNnSc9DC
C3AfI27RfDCHnko1eckBjnw+8TiKlhkCJ3aM6zWSevKL5itgPLvVTr73mospzFVWMdmGF2TEcpi7
sLoQJNHfNkCJ6TuCrMDocGGjkZFJtwOxmxw1LSdOciXj9yzIVBIWL/gSvOJH8JOdt1PVSm7PyurM
mNzif5yC3cWooqhWPEczhl3Qmn08J+LKVTJxpcUWGuOB72n/8V5BPvliXskSada4ZBo94F0ZRc07
jI0HzrDpHK3870248JtnIKSGE0m4PTBqYYObtzIyfbR2kvjZ2q8G8RXyUa2uN8Y8oAyjlt6fVa7e
99bSl51uHs1GKE4FTV8SQhbx5zbJYzy37KurL5+pQG2W1VpvYF/tiu1us7SGd+a1DlVCQ2MgvA7s
j8WdU9H5ExIDa3jCkINK0wEhODY2MZ+aUWQxOWEan8/jAgQ01IJSid7pzot+bNgALHuYvJH1T7wl
d1SB4JzK3EqOSmci+mt+/voTBpd2g2UrCQD/DsD+XEdMbIegWEzXy7u4glrO4GjRqRAQGSoSfl7l
pBk3rYQUB1wn6GhaliSiu3K33EXNWTG7T4bjeTNL0bQeGIyl123DsthL6Wxhg7x8Z6LHHutlkkU3
Kj0L13+ZA88lX5bY889EwcZaVJRNnENTatVEP+Iun3jrlme18MjS5qGi++Ge/+g4mqJpwXfkm9/G
2kmfUatP2K5YQJ2TmjIrn9kPqo0842sJjZOM6OEaRoHNNaP3Aa7YLl2DwXegEuoJRUjivS2odyDq
XNrJsfJKs1Umphm5evYi7+RIxRGNQ1oBr6leXspeRsCsT0VWXcEeoY/sG4OlZvy2kaLBZGqwUwzs
x4BbtnAJg2/LhaCdwLoAX4XfHt6V6Mw1+Phxr8gICvk2g/TlcP42XfNKrXJXqsFhB4b8sSmxewS3
IhdUWdJ0lz2S3eeYhJxA6BBaffs51tdblieOLHz7i6GEHGbgKIMFLzupzdMtmpeSpgAFVUtRmXpi
xJmo5ztGG2nCW7le2IRJzMOgZVuL7J/gxX3NcloVMjmns6OcAy5nIV3k7f2a9FVji1vS//wiv8oU
r7xtWyAtABoPvYmsD4G6l7XIXpPg0F/TbjYWlPaTEggVQh+lDQeUkAnNo7xg4ZdRCthm4ExcLd6Y
nKcJ0cpJ/40XngYc2J8G7w/9ncxW438uMWLawDXN4lDkC6mkWOotdfn+PrJ3ApOP+vquLE1eA+kH
aFVjPE4NQdTcpxoHfZUayXUVssb0eZsPbc3bW+PpobUzIyB5JiUZoE/k+5eVxOY94qjdeu9kozDl
mDNdUXdZrRmfDPciRW4ovQp8qSfVJjmzd1Cp4+VKp2qCmct3Nl7Vh05A9lMaMbyv+mWSt/ciJ+/S
/Tyg8AQBCC+ln4rbMO++lpr9DbS9zctoWn5lu4p7x7qSwlSSuOjxEfQl1uDHmZ+ce2jMxW8k2P0f
/TCpMn+GDzEgm9E8aaDXSSNsAK/aIINDrJLhADVQWILyG71opYEa0dKnRYipV/TwjnJsuBZQ+XOV
T0TkGthiFkAPTyeYtDmCu1fONL+MnmxTyzPxmSu6ESTbISUIlLGK3Ium8ucOEhLUAUnX8TeiAgs5
Kv1Z9GRLfmNUCQdu2Gsa83rlq97HwcFcyfum8/mvBL83xe3RF/VQU2mTdjEjkENyYdlAZ/uhumEW
EbAaDyrrkb9d0L9KZCLjxU9gaXjfnHSSIlqCkDglz5tZAeugi20DEBhirz1cISDC+rslhMeGD7iC
HnRGUjuKmBapOFbyiM1VsX92GQ54Y8uU/oURezRWIv6Y/uGyijxN62gZUENJSZDDZo5jSpGf1Hcp
jUVTgwOI1UiOTS7jFtV+uH8JFOthaHUyy6qtmoppETTMF8InoL0JwWAB+rEwBYeEgj+f1pVI6Spo
NWIrkzNggQ/USw2UOmM2TPI/eZYw9jirkKkb3ZXwQ74Lz67sV5QXPjXAV4Zz9LpeESvau4V1m69U
+phghit9FXUWjI5cv9J5xtZb5EbC7O3JlyGJt2yCM2jtpMSDbsHP3HZLZ1xwDzKUiNCKlqgR6Cw8
PodAwOK3Yf5U9gRg7zvBXXHiKbC2G8ekYgq2aIE2iSS/i2ER4IB4GI5hOAaeod1C+0dDXom4VUWE
GBFCTv7d+wzF0O0DKCQvNlkmLvVUrWvlBboX5bBKqZ89yU3xVtrt0nFEpTUniuEZlBmz6DJTuv94
VtD+O2bOuwHxNWxzhvGQDziCHh8ZwNPGYodm26gdulvhM0FkhMtCgxoXT0+oiZoKFVCgmUkc1Flu
dmc8solz6ooCbHy9KQdIS/T56aFqyyMElvG+3UT7Pp7H2b2uzqWTQ2d51nTZisC5lNX3wfnZpYCr
kNaUxXypXxBmcbQzaWfQl7qDjzlgai4FjyEawL64MADer0um5cPe/ZrYDYJhiskzsQMNXR2Pq476
yfj3ma+PFt0YJMToZ1puq9G3JjZodIicKL9GSJijEZPuzWkYm3VK7bGqzI9P/P6aJvnGkWdYRKqK
a+PtZ2rEBEWx+UIwHWGpJG+Q7WR3kXIwkKou6jK3zxnxw1l/B7uvKonKRMppnoYmzwwgu6Y6YJeV
QdQpO+X+ayiPLQL8w1iFXSVwh3tUNdjPfW0RIocf3K7KELJlZAv4T8+9ENc6Qv6MjUIH0TO6gV3g
1mYacwmEuhR6IWR4B84E798v+CAPM7LMOWXKgMHp/3qnER7x5rtlEtAy4yRfyzH7mz68bjbMcKNw
7W0zq9EvwSmbfU/aaFF5gDDY6QkvAPLZJK9SvbDYYaNZ0SdUVzLWTMO+d6tC7hg8wwzjh6dQRTMl
30nt1lUnKpbpZtO/DmWel8hBDKTpd2wkWqDLkYnqJzcaeEu42KiAS+VPkEbA03BVc1R5L6Ym2y21
fVmkVy8cSpIJUs39/MMecfPOyWTiOZhQ0J7TlLhvID0ROfVlwa4l3cRDABw9I3Bl+hUCHTZpY9aj
QE9JGEGMMRaPktI+OcUs3cNl0XKUlBlh1JlEL7l/z66x+CIZf9sz9+CeNFqwZS3wKzUooAZYC3Pe
6pEOu9WDrfQhCD2c9GaTIORo98pcKM/NFUlQZkvmBjxOZPI2HkIWMgsBucgKzpQv+6XPUR45slcZ
2hTrsXvDNd6bHd3xwg3Gq/xsA5wZk62oi+kqLxAHhoXM5eW1lGq2myKknXcCF15GFbHGAPhaCRk/
gil6b2j3/cqwasakbBPvICwZnLypFMtMEdw34Xj+9KbtD6bCKMWBPweYocA+M7NvmYX2cPZRNKjX
J40XBH5JZK3ltdbooo89sJGrWlgoHHLdjZQFPHinBupNEbqIPiFFHSJ7uzujAZSHn/7nk6sq9XsY
59TR3r4jh1DUKGhJDTYJValXxLmVmzdp2j7Y1GqlERF7m+raPY4gwQ3iLzF6DICDJqyjUH7oDYUP
+18+oFKtAJaU87plE6ybxTeZrlJcY1Est4V24IR/F/v5OIzf3YXETqaJik51eFsDZ/YWkmJ0WaXC
0gundLIrlQq5EHgkDQW42Mr9jDpbA4G6WBdiSFcunLf7kmRqNuHHrpcIbxmyl4tkvdmNMAURfbBJ
sG/DBAN/xssuPJzdan2/096DWy9AaqEMz056T/S9/Wuwem+agBTJzLmFjSAtAWxyyCT3nLWl8glO
o72USecj/DalG3+woNy3Etyd/msLlUFyWQspt7Kwmzz3evdaaR/jeYIaUg5YnFd66uRkQ/Sl9TCv
eCtGgoOzHwmSxcbMMhXjUB0pNH0p7ZwotO2ddVs6hwiRpCAJE1DgUudEtMtdB8i4uT9iQrGtDvxT
L5/WXDFX1kIOIh/dzn/+/XC+J3lH6+KxZIh/IsQTICYA23YFsAmWQ65diacX2RQBimd6x0XkyXbB
VKBkKqPPgMu3nOBvZjpn+nTTVEAH00NAOTvGahQPbLW6S6aWz5mBseYWP7u/R5XCqT1cBNQnAK2f
c19xx7FUg1mIu3cf2mjWSdwYfpbKu4R+BOz3uvO5vWu9NhOnMM4um3QVmU1Pl7MeoXGr1D85aPoE
fJgIw3Qd8/D3EIqP6ajyz+QwjKASo8pYLdCivOY6cuy708/NOt9ytBGjjZeTyTdlc2bDNDdEqyKm
4n3ugMsmCD+cdvXEM6ZyL0hDf7HXKT/43bj3UqaJG5vrJ+pmo20/iCSqTo5TKcGbMBp1wuDFYQ3a
TW2D1NarANyHn7pGO62RlmQBlXEbTejMEFsF91ia6AXSgglhSJR4BJNhXHH9J8TPNUPQc1qVSnnb
PeGlNO95e79SWV59ofBbZOncPDuWFslJ0Csu2AXlio3Ctm4nVwTcS6r+R98YAekOpShwNCpsLAQX
WcmSTCE69XpPMVm6M+LP788efwsEPBBx6emi5Z3ymVuW0wrJLQdQ6DHmhTiUB0EXl/UbAPXQP/FR
lUXDU9F/81mV5CHcJTjLiQBeazkGF+S59c3i26xWTnRsYjfj0i94if0zs1sp3oiLqUJaz2SMbNQQ
J/20aUPtwOAB6O404D5C31eEJ3wyOd/0t6A4fC+RuqNpiKlitPvyuPdA2AuxuVDBNbQy82yTB5Oz
M3nhJvr+23DRPYSW2j+D78PkWFny/wf9IbtOfQOMNh/I8SHewfpELa2/MTu/+Zw9eOJS7Ky1fjLo
3dv4P1FaU4vyM/wXYtxqJRiuDXKyOzby6gOsHOuyH0hVm6Mh5Z2JsSvC1nOlneXJqPXlBco3Znlu
EW8aq5DaArBJPdSspj79VNSSSVausDT+/4WG5JjUbF8qsedpeITo4CfT7ogRO3K8dOCyJzbmlzm/
JGQfJ3uuuHoEM96Q4sgxB+ehFljnQXzS9d0zO27MeznxSX5iqA2aiBrxUTVVoQCsSV4wpA/GS6gW
4vSvV8Cg9ovySUcD88UyMdkQHTCkj3Ynsso8B75reUyuPKA63kpa6/YBNZhwBkvEsyfip0Cb6TqF
c6COYpF9I1zdNruMV1mQ8VJfVIvIXWYdYpZRMgcscqdc1JJBMD8uoKQPcD88cPJP/TgrrsfoyZ4Y
MKiwnB7oz3jMxoXqJqA8qls8LJbF6YRu2+mDtQvd4lZZQH0IFqG5V7sxnaqkg0ApnFWNiDHA7/LH
YNWJbKLogOlK6s2dtl8haY/+2ZyqPJamx/6AfvALmNOkjQJnaPT8a+u/xCiH4m0EZAxlDAR6garG
abj50WDc4NitS4/5eb/eJe2nd10gNZd8kZnkDUribDz+3HI4T/uML9jZL+LWoRnAr3lxMfb/08Vk
RPpeUJVfemuAwABDHQfunobTmhGLFyF0021UaQlgJjRNbkV3yVNrrRd3/4XS1cdhw9RN5hKaS+y5
Y8nmIOXiPCTiReaX8zvhXylI+oLWqClW/YQrZnsbON1jxvU7qflN9FBYvSTnM4mtlqUXHnOngX9y
UJeGcLSAP8ZS7Pe5351Osmjr2kk0dyH8x2CGmf543ixGeh/Pp9Fqjy/UJ/Wh3/5wuNLNHUWSxz1+
q1zcJNzvsHlSixuKxa7YWNHVnt9ddIayyA1Ug4Bq1Ei5W/jnNwQWyuOlVK6RGUoqAe/vdQJjODFX
d3Ry1XZcr9+Vg8MFpIii5/uvm180CZ0wO/L1SWGQPRhWlR8eoobILs3vxzepVwFiyMuj0Rg/pi7o
C1JVnhSA/JNp/n6KzDqrjBBVW26Z6o6Np5dD1ErV4q1NywFFD1juFONWiji9FmoR/cfvt3SCORv8
R6pc4Sr1MgeJEv2cRARUCAMkN+nkYm+nb64w7x+z6KjyC1CLMSsnntKDlXJOSwso2XsbHo/Al1qk
dsZ98oMR0X0ODDKOFClmbmTPTorqTjwBDdZDn85zGj2LPB/HFAHKcx19o0f039pnocO+CN2JM7ax
HkJbVwwEL05BhkJIsQX0PNWMGVAbvDB3e467dWKhsnBPhdZqIaKIBt/WWTDjol56RdeqRlodatVJ
x9N/3D/KTZqqJywVh6DYMfeiWaVCUBcp0uKYv61YQN5ueUgm4FO+e3esu9sh8359r+kra3Zw7XWm
1NEa5Ns373l4LhEwjnLHgsgxkWcbb1DSEqppf7X/TddfrldM5EJGhGRdiiidf1K8SZppKlG3nkUM
QbMejMNE/1wNHRrNPFAmhl8AdDZ78xgtMvs4eK1TsRoHkgIkwiyMDsiVDFm/2o1UzhsbZWWw7Ya8
kW3/DNxfft+FnEa6Pnkiv2DD8E9PFVt6OHhtV+V7xuKoAzwtgvxowjECjkYhCWuLl+UPjR4HCShb
KPilFe240SaZsamtDtdXvD7ROgTgMoxWQ1dSKx+A5bEtoHfhQxHCMYFKgUVWZ0zAXT4jiM5u/l9P
WIoSiOiOA/cGOXISMs+luBFygQL5eUup7YaFCMTDxU38tZW9+kDPgcUQyfa9fPag1csqV47fxEkV
ZZwd0/qetfflSu0PPi54ZTE5H/gmbhR8TKNxIjt/irzjry3kvF532hDRon9QpLvmSYvEKIEH+KjJ
Ay5pI+DKmQLhozA8Km/Q0E1Va3n+nGlZ4rpwOn9e3zET1tXPuWPZO1Bp5ovRKe5ucwVo/niJ4tAL
8XCt8Ne99Pxd/l1qx/NJmOZnZsX9noXjThL/e6h7NuVFMsIU3Y4toIHZNjAu5EYQyehd+aH0CM23
U71Lu/q7D06btS5pn8xq4Wwydeo7yTlTTsq01T3QiElIvBiVStN7TBrNc84Ym1VVvWPblfY8mP3N
XpjiQi/RatojQCEelyrSD4M58Nwi+HaD8b6xzZjct85LSuHQvSRkpTe2R5IKw2FKGOyzJEAsPF2g
pdTO2dvpE9KN5hqF2zW4M8eHBK1lCGLI2H7pxo/ji9RnQTjZTX/0IqVUPMCqUf1KE3l6RAqU+jSM
fhkO845O/e6w/XPkN6KFwuqJDTy5Zodfq6Sd6y7Y8dEzqi24k7/c48hmmGJDv7p9IxMOM0PFDJoo
wGtUIXe4OFVvNh/gb0sdKTFKvlaNpTMB6xX6bNKT1920/Wohukq0JN0rPPP6WaTBxoKiKg+yweaP
2LQbKiDgMVV055RD4tEE1NGY45qvdAUqeVZkOFmtHsjYz2LNuhFoZFufTTNK313Fy6GRI2NVPd+e
Ls7L95nFCkUXf+R6U5fPAM/su+uONXky4nFmtf7jYpJ4IYJ7cv6j4gC7Z7o93t4xfiAyhRtnEFzr
wOxEZ0jWqFTnRMP1SWuN9jc0lPRqhQXhg28Bpkhjs2rY3zSh22XWZ9DmLniOqKdf4dntvJIwWcrW
XqJ/6GRbLUbxVyKL0wMP9saD1TmwfQ1rMQVQVLcudlLY3tzZnToSQ+sDcni13UttXm3n20fO4csU
1+amtvokmEnx41PT1Jy8QyUu2Yhh/uRoHhkM9/sAzKX1f0JmQjO3+jkTUva84xzqv2k9tQ+9gzpt
cVEvzUJ/jQIqn9E+h8AAI1TxJ9htIMO4CqbvJPdV5BRxBtZeP94O4Jdg0euSTEbWp0CkeXr0iNGt
Y/g06HG2qMrDQ+H0aNMVoN/pFgvLYVud45rjnZeenFI3udji/SwQLfM3xidBcEHErIJydWL2O66r
ct5OPN9B1ELxA/983wV3pU9jTCyhcctzc/vi4id2ngde1osNkWGoLdYgMo/9uMLjR2Yc/8rovdEP
dCJ3TpNL970VXLLo9DPr5DrTC0a3r4n+9KRPXMHc0w39FPRdrAcATXqDWpFdFkxk7Jcy0BY5zZn0
xnBW5NnesUw9o7Fv1A67tvh6HnG5YDrJiy7bC2kV94SkavEyeVvcchtuyzO08tfg4B3xngzJlXaQ
8PA9hfAFS0jb+6nxaso7ea1/A9CiHbGRKGBwHkMayZXiwxZDxuWu78UttVoxtaJNHTnM1X8vOjKg
aL9Jqx5cg1n6D+fynlsp45NWCnqMSJzMp+NGyUqX+XYThAAtHEWVtNxK0wTTba6YjoSwEAIWheXq
Me4doOQHS3oCnyDUkrOVcYWl9k9I6z4IcwBtM5gGnJmg4ui+2VrvDYaRTKM6lzM6EKSviJAIiv1T
GWOeV7gGVB6qx1uCCRic92WkS0js7FVW0+ZSmIIxwz27wc/6MPZ8mNYF8yRwvv77EgAkFhlju6fN
wiiCWVQ8kee+gVQFkD6QpDuyZX8u11A70gDKCCnMkhMWcTRgXp6XAz60W48anyKvf2c/zxLx+C0f
oTHGjPFGoePNfRpSjiSkRj9h9bV/sI2gvW9dfMx+bDS2p5kCR8ktSe5y11exscSME7PqjXlx48eM
vt7ETqLMFptLJFCGpAR3gfOCnx+OfJMZ4qLpW+8buKs4DjUyLpkPufRjMD7szXL+3kJT7sQakil9
PZfLqRm3Y2XbAwQCbXZYlaf1+9lgXSf10eFhrLR41x5NQtdixgTXLXk5Lptu8QQUleLWnT/gmKvn
sY3SgOEG6OlKwQJSueWDoJdVNUN9sCvmuKVphJR4hg3lPNqkR32jRj2VVO8Vo+X8nwlu+5rkPWtU
b1oxYJuI4RUiVoeOwkIFMb8NiSttNOuPVh9o+LsjaqmLvLRgfkPIif2jC2QdRrGU1tVjD9IkZKij
WwyAomKMbxDrkxqkpYbdo0csB2lF6ogS02JWPuWRBTI5/wgUeNW30X30HaEt6FNiwrg5Rvh054OS
rT1FSmFV6FKvJXPZdVDW0jNnyycZX2R7qSYJOxui9Bd9ru8LLVg72nfwQa0TPcGHoqkpT7xzje3T
ysS0MgGe2eCeXDs36ikMtbYqbusGSrNi+VRSYgyrn2MlG3/Zw6YTeW4XpmPdgQJEYu7YajIgruFp
i8VvvGb/pgIJJWn+JxQCbvKWG/OH4lNlGaChrlEN5GfY5MJBnFGPxJVJykQ6LrsBQrgLHWWlrrFn
5/cOC6rYZ47Q5kS47lQnEuVLBlLTtCPreYDH6s7rOfGQiFvVS9sogSSXxeVLFF473n3OBDRLCzL0
jsSchAcifNT6RtbPAgL15qVpdDyFXL0SjstGwoIt9C8XrYdO798WkfU2UkwLs6rFL9yTlOhl29S4
lJoI4FVkNgxj8o6KodZOP80nLFaLhwxwqboHL4li49qJmMn34gfe+r9eMsSsjkZOnMNoAytUWow1
ZSXA+JUCguQEvtBuqCFC135cj+EdVDUYgMDPsNTyferr5YV/dqUOkrB9eSsyaAzGnFDnTPQREHmh
2zRl4UV+LvvdCcnTt1Gxtto1PE8u2Ib1cz5cqLo4pzSZogcRfEcH4DCv0EveBpMcmPbd2pL5UtKV
EgBzrusaFOkEorI6xi/xKqQEff+Dv67O8BO+7sNg0vGGkguECpxX3g+lxtt89ZCtSJeN/REoH4RB
w6iOGlkxQW/A5bIXxODKcd+nAC2/OluwDfhMh85M/MWcGiz/5O9mI97U5WjQBJ6Biq1UWvztfd0R
1QgAzq7Km8BpV9dxZllPxWIUZjNYF3DgvsP0evxN5HtBRbOkniOBWw8sWCjT71HzA8XMFt21tQn6
Xtz/ggUeWcdd3Hx6e3uMlVl2CjbqeFaOcP06IICtsthekhxR7bTZy9J6PSFZ5WmQ6QeFPtawGglx
qHf8Ewou3HeWNrZNxE9dWSC6KdfakALA/TKtfIpnl5UULKTtN/5DRFOaNAuH7RXN8ifk3VCcWD2j
/6JNJiqSJaUt2HdaiFFOShXwwQYmu1ifEL+/2LTs35syYIgl44pVdKJM9uHGbvS9iGo9HE5xV43f
xrOzUM5ao9t4ATgRHCFdRoXVC4AWLNSFUiK5l1hwXdu28S4bLyeg7CsU4rUcmkHCj05u8RKyQHHJ
BqsDEnhFIm9v8H5iOPx4Q8INR/pL9DmsJ/tIVRfGYvIZhdsbb0KGdBwsxpAwh0qfU0VHkrghG74M
wBdvZYqvYivXllfM1u40YU+sX7jUqDUFRbK+o9V11KNoiHYexBGt3VcE1uk/OitCCu0ChwP1EhR9
ks98XLHgW61JltjYkhNy5HSypCn+XNnIcEOyHr13yARF1ag28e7Wg9iIrAEm1sxK/mEIVEJqc2Ph
xnerlo5GiNqZ4Sfr0WpvYEIu8W3xanxye7Ar8o6qJeVlCD81gq7JOMqKtNAQeIxWHLthWz1HSpgd
Mcct4IorwOm2xQRN4/nsygUOhiRyXdhPvT73nsI1p9dTlpHQJKaUNU0W/6I4VumyzJwL0mSipW7U
NjXURXe9r+fNbS2Q7M5FIBxyYp9OiDp/F14oJFaBOKbN404dk/eSAV7pa0F88hy9+T5TTbuLwmvj
e7Ll7E4fU1bKJrbMY6fC/qskgfnCcIwonH56CT9SFYD9s8NV9QfZGhFWyxjBXw4yu4IsbeCaE1xn
hMCYBUtg/F6TliPcSzrzG7z9j115nA31mQ9/Dpd7tK4qj/kSrYolUYH8j63Xz0l9XHasqRijkXNF
70NY6WmU/jdcjD1rGhUxvVwIV7BdJy7GSA8tC1fhpEORiHR6WEns0ajaFliJZif3JBynYO9CjKga
K0ws4sGoW1bzV2rs+hTq/ak6OHaPGO9sO2ntJbXNoxOfKYBu4mtpflFS/itiB/qOdjFF6FPvvvR8
Fjpyo/13eRniyhQZ3f4pWSwXiqwk3opGO19TPDVPMzBT+P/vzk5/4Ke5NMMk6ryFKyirWzSN/Wbz
+sYZGlVIXNqb2NKTRQzf/gDqdCvlqtAV6UWyWnGBTDX0Gej/tb/WvcC0jYvWqzzwI828WIHyXdDa
r3HkSjjOlCGCUfCDjhFd1lAhSquUy2giPxe+/brpol443UJeUg9PO8yYSEMcD/EOXfS6hCjQbcGA
sTu/CkRZ+8nCN4E0LGRtsd07sBg+dxVICWBJHbBywjJYxqNLhYr9peCVASj/Hvo8w/yuqAZRPJVY
ZIhRztN+4f2PV0JL75ADlzK7ZgTwwDMxUeT3HgZkZKkzigdEhp33eHW2tbGGpNO6a4gsrazQwYXN
RZGnyyB8UbcV4k754qfzsKcuN7yoFmg6p6D2ZusUN0fNKzT/qNLuAI0kzsdm5li9svBGE4pSFItH
YPFdlekylZmWHSzhvBtZSxFYgNi5VlhFcGBKbVPr2R8Xuqhy6g65iiUd7kJCGHfVoPo3puNIMKng
M7We93inw6+us0dIsariw6MXR3qYVEJzxT/CFcvqgi98To76KEajngz4CldAD3GxJdAsGch1nbfq
C+Ypm2BtO6ZsrKemvsJfG7CY/U9QqaqCggsqxCi4myn4LUlrUSHfGfx/YybPLC+FoByqPd8MLMl6
2mBKlOZYh6LcEPRpmy47oh5Fr7pmkdfXFQfpENiGgekLe2u6s6AfgPF+cH1JcQRYXxOSxpcDi1R0
Uibt65GUQiRgT9qPv12/TEp3Ss/RF47w88qpSKOotAFbw9FjT2gFh88tV39w0cP8UMJl4ROW4kTY
MulMW/KzYVF9e+T78HIu+pobcVDs7NFPhKF6CWc4I7dUWlp3BvJsgMGkTUEoQEcgJ23gP9i9365I
YF4Re0RTXfoxTVjvayqnI3Omd/7/wPFvm5SQZtsNp9H6rZIDtXHLRxdQLGyNmdmyijYwnR8ErsB7
C1u8vFQCq4dxj0MJBCbGhOLFrORyiHCTsNGxfaGTJ1vOWWWycCk65Zwqio8DE5d/YAD0batI1ffM
/FqUbNCCZmZDThN11mFZvyXfUqkNtJ6BadyaRZ8R1O5Vu/0xOTBRURGz/iSQkvYDaEEr7sqm+kcQ
h3H0TiJQZJBRjLhBKyNG4ss9Mqq6Et7m+dDtyl1HnHYn6aDftJdV7D1okNenoA9uafmE3di2K5ib
cUwwTF/MW6bXhJdXS3RI+UBYGZcaTB6346clON4hSJKX14usScMT9dMJmiMYT1JN8RwY5dd2rgW7
nFrNKAZfUas7RWSLbBoyBOYqUlJiunImEVcrw+o3pfH94oc2DjWmVIMwtRLHNmRGKC7Dlyn90aZZ
+uVvQBz5soz0YD2uQEhnY0AuQVgzZNGiOYYagj6cqMVToTPAwRixt3jtDJLHE2U/YFwQRgLotuIO
0DZYuCoQw3Nz/Qwpd7nXwv+gAmdn/CF2XDJpeFnM1YHuZr41zkg8Df1XJnVRgYx3ifQ/QwQbRi5/
bWUWnqyipqgPTIf6vho/Jl2KMRD58wd3HRKw3O7B10KJxus5dEhTOVjhjKZhSnXCjUsolo5yk6ef
WyQvBQ5UuiVDw3QP+XtRUcDhhdQ4RSSx0Mo0gw2ADmXMKgLPrIEGqU2oqcFpIZdOt6uHL6Tx2fuv
1ocdsvp/6MMi192Bnn5Sl23HiBVYh4ghWadD0aak0gQS3VCkoS/tRBcHzd/2jNHbXb0EP9BjHalr
aQXrpGw29Crge4ChepWuqhoUIhJc1JerB4nVM0wbH0UZ4eMZlBzWqnHicn3OyQ5rmXBdIZrR9s7F
fQ+7CRirj0g2VJn1SF01t00Fh+DAzzkDFfuKkHpMbR9pcwe1Q5xnblDPE3cyo0oj/atIYstUjrdZ
+EkLs7IPgkV174FwVZUvGD4DDZsruN+yreKh/fjTxxS1c4H0FS/vxRRNL7O9cvk4scOvrSEMkMGd
kwgmNuTkFsjgJ35G9ERVxv/1JclknlKQsiGFfXh5ZG+EqwQ4sFVdkTQISUCm4/Wh2Gfcfx5f/IcH
iOIAmmzzji+8o8opUEA+w+s/j86tAT7l07gxAIzZTM8nzQOV71dpdCAG2alfZMdGsSrakZJraf3e
iMrCh5123uXlNKhT8kTvdCdJWxyHD+x07dg8U+6GB7NRI2T0cgOb1eHohBO0FYspKwxBzXWOGbGo
0zgyC/fZHcpHtKAl+SRHFXs30YcDa7koqSXuxPr9t3r0A+0BDcGEkWJ6Qa60y+hZ/WeZa6pBlroV
arb5VhsK8G8RlMf9pTC95ogjqZIZJc/K3gEqmePNcYyDEb3dvK2/u5rNIVv1JRroEi3HCuMbM5Mu
glQlzaaCNN8XYHYIE+4yj5EXYDkbIVt6jU2+8Nw+v23CrV4jxElCeejUEmNfBCSxHtEPSnxt3HZL
Nxi6HDe50BpTFqBrP7X4GEJRZ8URrw0JfRRcNCpf0NVLgj2kZOND4O84T2nRDEAgIl1PDYbVNOxC
5E5SHGN0uQlHIQGr8+wILaSYBrtMsBbphATTJJxPfF6j+8yn/KWkVOFd0JFbH6+0/VUdnOQMuOBZ
wHv+A92aVw1xRIAcIXrcCQcfKAGXCDjMKA6pucuR88VKKezYa32hS9Gm16w03QkQPGBbx7fNlB9L
IaF8SGmU56xuAmuu+FQctp4/cUka3wKs3MkD+uAc2ZFyanHq+eJdIViQvoSWvWqhbwJdhuoKIaVZ
CnpaEv0lce3gGoFPdCrVSDAYiMnC+tj/r14ye565yQRTeavn/h8kOs2KTWOr+nIr1r4pIpVEpbFr
mO8NRxx99B8VPZemu/qJmS13ioUXPYxFehzcUqFinvwfpAxoT6jZ5lq31YgkObOAMVoLMV6Kfugq
Aqz6RnzxFMBo45W8KM7K0H1MlFHjxqngSC7ZNcDnG24lNvJgogzOqpQpupH7u8w+VtCPcR1JX/YH
Tzw446CQ/vsboVm7LxR/pXb2Ex1cUxaU5o2ttvOx30EXL1vEjD+5PArHDsP7qNhyruZHT1fk9FPV
/ow9irknj6ip8tZC2tbPyapePneAMxJv5sMfuXqo5aI1jAIu25iEkagN5gb3wtLPD1hsNme88QCA
4vxD/l/4BjNOUnPoiPK7+KGnjyr+PY6S8UcUDSFqD47AarLcS8yUi/Ms4bgnB6/lVEgsIJt+jy0P
2rytbPBABJBDboPU5GuSW9nhceZ3HeoRHywPQuYeAxRyAh3lgBCBc9tvHBon0NqFfUKqfGbPCzEs
TNVcsTURSZbAckP3NwjvLlRFDUlNQyUJF55kbqr5ufYEOwjoCsMpNW9IhN44kbV2dYBM9a7fnWHj
rD4KvSwAJijBZnVKzy1zcliFsSrW5aJtpT22hgLVcTVGsgKcsrPSlMMRV24F7KAuW0oA0KIFsSt2
FxU7N/aSHJv7n6wT6uBwBotuLA9L0ilPRjNkev9vMA+WuRbgF8lJtnYB98YUqxoudOYSQADI8v6f
zNnE3XyawJwU8luhtYN7vP2NAnBuYte9mwRdaYgs579d8ygVDGg1gt36ckmwgvh0lT24JI6DG8vX
NkdaGzqrKzHRpt0jD+pboXBS6O+fQE41VrUsoVBJS+8I7RUx18Sa7Cz8SNBmLby2Z+lAypkmVp9m
MfKPCmAj0rfyE4yrLemVrzH3KJeXsmvf+LYy4mKYOKKD3epPk7UOclxUhHQkZPz8+0NPzmWLCrVN
3fbe2O/0H1EYJH+X1tiWdSMf1++0CPYJznnmArLSGZUC9QwZTJOXSICxPphnMrLV9caNEQrANkZ7
IXZpEpM3uZnqq9nFh7cRvBcXn+IElPi+P629KQtfzW+pje/9fm0M943PowWXZ1dufYq5/jiD369j
nuoB2H3w4QvTAKRdAYCUc/bajqiKwTHeDMKqXh8Fy7d8s6VaHYI4gCTv49DzNa+55nSmk8/K2XeP
YjLJf7nED/Qf03OUKijwhcLXAhtjInxJSif5TArYSv8x+AQuBRiNeA5GdUjbF/gQoyzfr+tPscmS
y8lhp627I0YSiLli3eBsopHntECv9TR+TOO+pPTdFUpZ4M4HqzZKMqow67Ulx0dgKJzllUdNRzRB
JVIciY2ZDSpviPclcPyn4GSlJKvQiIbdtRL5eaS8OBQYsTVrod6KYGh6HG9rzZ3dUn8HzC8TrUDQ
NuXnSyOjXiTpLCDYdnOELEuSkKLXfEOsqsOGyFw5km6q7+RbW8DV65qXg42JPE2znjYOak6df/yq
Tjcq+P93aMaDXRfXaHLkd4rD2PpgJEaY+HJdxCl+t4sNV0G5cg1aib/8sHlo+eiMYz1nuW7tsKrl
jv4S2z9tTHuZ24eONzq8pAY5nJh+QQf01JdO56gGpETjSaDDSC+2cu7h+8HuJyByVCAQ+S0Lu53v
yUt9xQ0NRkM4ixZQYGWTMKh/vU+kzczsAOn/yDAoxpMTcEboB6wsmpLMSHcUwGR7il+PBY96Kw17
SXn67k5vN2/Yn4kpkYHykj5QWW5LHjMT6NBsQ4JQeUx1kvP96Hkbrm/ZApAuys0FQL+aby8ywCOQ
YPHWCXJyuHYyIpXrqXvNaAyC+FVfmAu2M5jHKa7c3VfBC/8yOQZvlS2l7VGDtgZo11QKRA8kiYuy
VueS9xBZNJBxXjXm+SrxxgLYfVRNphw4hPxkx/fNV5gyYOTtNqqUnY1u/QumaIyha794jo4pXb6G
m5rcM0uEDve3lmAUdL8m+7M1bEHS41aKPtRes60m0aqR0iYDerdMULqOR2QZK4xZFOapV6hn7AQ3
cwznyFaTSKvDeEpx929njWlAnQqtA/z7m93Yb9GotTCS+iLxXkJzGx28k0Wmi1eu9IuKR/J3lJva
HOUGJN5AcUWDPUqDbbZE2OHKrSumDr8MoEpLJStTQsQOXOeb3IZI8yJGwaVioZGlxusgvrddDD++
4buiTYw3IRth08doAoWxZsJoihxSE7QUh4bGxiqB9aEST3y/RGj5WqM0zjexPBCncrx7lPV9MUs/
1TDlLGbNauG2S8wS92nh3w3UjMkDUje6lSIzInvSnavZsMYL4sylqmbWI5GHSGURmAnNbU6rG7QN
13ZAS195Ykm1YTv1sMJcOGngLRrRktzxw6J8ayO3QqAi2+Zs5hw3XI7Bydk93txWp7Zop0izAtW6
wF5mUhvMpMeFrF3YIZQ92hG6twTyBmzetkYazjIIbOgf+VIOfHL1de2Byg02IBUC+2MZ9bR8aLEc
YhmFS6oGWOJoPv7NjMZqhAlv54pLrKuPbPxLdCes8VMidJ3T8LgvA6W6VO659x5WUrUTchhrj8nT
jUm3xRIpBoCDEjrdNyqnOsXLpVSQ39Y+nWOIoQK80u7YlOZvHgN4aHICpazonkLGqLypeyvCIW16
Pp77wsLVkGV2xhtfKtsREgnfVPrdAW/1rNBbVJxe0IA0MzY9HPyNJ1SMWKRbtyvOV3/y85OAlVrU
XQL/M6FP9pSH/9XZ1oXjqVpOa/BLLqdWAfV5oEsqVd6bqoB8WrlN6byZ5oGd2ymrOFpH8miFoSl3
tSNjtzsWYjJHpEfIhrWiq5ymrqlIX4ofWM9D3G0ztFAoXQZ1bByTaJjSfCTe7Hje7XDkpVUSyKQV
W56e/zdTGLxmTSj2rwXwDWZ4QdU4xOI72QjqkTtVWXp9gaTqksG0LHwNzWWIjWlH9j2bWmHLpw3x
p+WU60NSPvbuuOn5/zyhMjfoBFW7v4RNrpmQoW7KhfB3ITIbaKnDr3CuhVF0VX/8hRXBsc20ry7t
MG+mBI8lCbbUIoID/1auNL1PGjhmi6IDG3OobT4gTEfhfRKVCdbIlpXkGG7TaGgQv/QYVzgMsgbm
6aQsyjltlzYLdnXXn2dfeJ67GB0WSb677EjygNAvXk5ZyU7MewhbZPPKbq6n7QdqqT8bLsLRiSHA
lshB2MqhcS1GBFYGU6nUXhpBT7jFfuX8QWC1RRhXDO2efeoh7KKtcGgFCRJ5fcm975YzoELSkicH
AeVlf/2vHSw2ZtvG7vqeIQvugbGQi9/mjmQqkgwhnXb+qUklCtiyol4ySzQjpuxuUgywJ1x0TzAd
YZJ4pmTWwTWQ1GZCR6ji8iG0/iWaUfh0y7cG5RRqnFtgwxJiuAoDDQZX8rldXxoJmF2krEJnuCjD
273xihJkx3nXCuRdtp2aAXuzy8ti5iYiCn2zAeWA10gr5XzzMz0uY5AJoWDE27GgSMuzwfeWBdB+
quM6xVZq95pKDBOpaVw5M+hQ6McsVYqCBUW2q2724lolAtmLwUcBfniHETids0KFOfeKOcs+CPSr
BorDmmbESIjZTrlska7r8TjqF8XZ+q3S29Fq77CpW+BDI59AdjCIYIAUfKk+oHSNHpaezDIKA3I1
3Gv05Hmz77bQYBbssAEctCnqFYTIsRNHmmHE4MFfI23I7dlzVkaCa014bidPrfaMBnGKCPooNMvX
ddoh4RuVkqVqoh1VWtz349cDn3Du8+OGnZ0unbISxZ4i4NPcA6kW/QfcJ0d7OHnb+wFIklgaCSnn
+0iFAUw5zcKc8bZLGAXTbLo7Nl7MlR01gl53xCADXOJaXR3tS0+6IKLT9Jqj1sBW/2bzE9/MYwfW
F3gfSOAV3nuzl3q4GIolUz/7RM3/WX+yjSpQEe6xnVf10SKUWceI0GUe3gWYXOKFOv5ep1nRcmpZ
x3UkNTXUNeIXHNqThmgTxW8MkgkmNstkkOsig/3Zf0Nfe9OOarEcBZqxLwD+TuvxUUW02wyOHtkN
+iLgcSPJ5l1rEm2HkNWEgIbv6ZnWOOgsVx99y0AU1jKCywvIrDStBKiS8GAxXM5/kfpmiE0mmBUR
FICWVFH6Bet2adnV/KqK5VHOJjMBAdLupUv9hRQErJPACpdZNRjCoAnV8JDqTLz/7mF5vlGtgunl
DfdJzcgOgN3oS5JpIKMTepYvOX337/vtRSN3z1NA8/l81w3CILhdtEvzj2vHrVRABv9KDS2BhIe/
IJUDEmI7L96VWub8uzau6lUMbJLX1z1an0ItzYdfUpB0la00+ARGl5GPhJYeejoBpf1BhipkaRrr
dTJ85BX7+UodU2O32KzxWla0yl2vj2RKFe8UqM/mbrQr9qQfTOVMNbonFco37dtFuO/WyaltssgG
l7GDwfKtp0wMp2DKoTrwVbvm1WB0TpFJ/LqOxWLYsf7bWbRJYjB0zZsvU+YQ1Bk9HE2nRF1X6hzv
K4GQx8SHUtpI3EGooBVkixNuRHygAYc9aFTIhqyg23p4A57f6C0s8pnPsJwmTfymHr6fTWWCz+ZT
qOqgQpTJ7UA5aQeXRIj+DH3cXaGT2VTMdKzyCDQvPyEFjFSbobAvQ0BdIn0QZ3pQVOw5WaXpdEOj
xMY8pEW0q4mcS0QR5hChLl2XJ3bjS39guScSD7wH3zHqGXy314s4t2JVJMglv365DIBKD+6YMcWM
dywMe574q8gLRHIXA4mC1VRwHUZYlB8SreQwX54rXGVF1/l9Of4Wl+tYhbJhLeodjOUEuwAI9CCb
TPRX7hrnB0I7q9TFQ3oeHzSCCR/E8v8gQwxW1U1HWBKOy6F7vaSi5PzW2Iv9bZJhByEUymyetco4
u+foM6Ydog76hNSTJYyygUehjWgc8jBLyr0LONPCtYV7o5ykh48Hfsx9+yrd5MljytEm9/jOwQf2
4wXbJbm+1kogBd01CXabj/ho5s1n6FsbG2Jwu9LFHht4IWxCcnD8DCnIenlUIw8HEt78q0lpciXw
dBvgRharwNfKq8OQ1L3CON4zrKbqOnkwpI8hKnnPYUPabvUeFOl7iHBl8RPCawyiaWK2zczF+gfr
Dr5pqoth9l2T9XmCbf96eWPgrh3xzTZvn9j01k4Yljg8AYbI7ONSXI61OHmIazocyvj8X7nO/l0H
IfWRtnRBqRIFq6xf/TYIGoZxd7v40Gq+d1mSoq7Kjbi8Tkavh4rU+GXDcOkBux9POhFWsCsgq59W
tpswiuchSuRUwqbqKWNJ7qY95wBl5j/9Xe8g41z/f1SU/0+WM69HNllavyOr6zHfpEqI585QTIdy
IjH6t/fLNC3sjmTmEOXl/XC399Rg8hpAcqWz7RccUAJzh8EAvM4sxrzG3rOZq7ckkaDZlwYmMU3M
3fngnU9GD8DybZm+WQz8FlDci6Q3xb9FpbsF+lrL0ze2Tq4/amXHt4uAuOPFCdUCka4kbUkvAUWd
3SqVXejTCXHQLrs4bzuKBCdSTGKJdmFFfskrruPcxnwCR9iCg+/TUVuskCi39kAPUM4blvwGHuZH
4jUZrG4SwhNgbVUnHGcrqkSozQoFsDE4LcgClNmlG7sfAsnTPXf5L7PzY9QNfH3BN1aPbrnXZxVk
v8EP/UNiIyiZ+wzSHy6yXVGzUREQeebZ9MthDAqsZsrHYwpFIogLSg2aK3nS8SZmp99IghFEQKFd
QY+ksJ7JnkcaiDwHZfEIT4BhNg83f3xGqZZE9MXRNi3fW5wqiul8OuKAu+IC2zYGczzYB0BpSOnP
Xzz61zgXGE/7FXv6S8aNxYZdn8ilSnWV1P63U1Dg42rkGNiIAFThcSgaD2KYFw0j8okO1lBvYbgn
NduX1F5sB0RYgx8mNg0Z8AXovBBPhzgwwMu+hHIcSV8yO1Y7ahYfit1IxYQURv5aTTsg+tyQOKyt
96OMCiKd7XTGoVVvglkafOBgxxLy3cBZI3yoAjDh2S/0tHD8+E76r4k78rzi/yAtujIVDUE6TMwR
nHVRsogJ3rxoW0kiPoLNHpVu7mOodhtC5j72369Qo7g9HbFJjK3Cbw83J9uLAWekHnmvrWbPlbIQ
QPKABEsIs5s3mVbR4mnfeS5bjLp20kKVIIBV3v9rIIYNpzLHILJEaPXd2X6+kxJRABhJUUk/zxQq
yYcFNa1PXoV+3gIb4pf9z4AtdMhuBIwiF3It/hd9aABnK2BUa9SNs9HtqhGMVBP7DYkrjluVUj1E
RstfHApBbW/CiQh3/IwExNwA8vDocuukqWGsuKHf3FbHD16xy9mcNj3qdQfcC2JkJmk8qe+SiTWG
TvPekXnZYp5/SgWwnkQLlBwYswXa4t9MdDLAhP7Pf6y+U+zVbYoeuiXZRI0CUwassop514+u3DQh
aFf6p3nhkaLvVc069NYWBTaAbnCtoKcfcHOFaFmAVMQ1okd1VCPAHfxW1N3xolO4Q45mJpAKJRHm
+QhsDziuKKrSX5friZ9SbMP7HXnswQWUMBl351Qax28rUhbS/aUHjnkm0lL4pXcwbgXtfSN5vxWp
uhawtHDcLd5k6CHMBHZrbVs2mrDdu+NjEYuOllUCDHfTXPvlYdFFUzTJH4rDm1CPUf9wejfv6QRS
LkyVJCrpiR5PIPUhHs/S7S3Wm9eW7qLuMAg2bTpZmK57KPNsJvMcrukPjxRatGGjkoZGGSSdQQdL
O8M9L4VaNlUme7yobcca2oa378JkWz4HpLa9tLvVRmPG91iNomFU2VaGfX2JumwPEkbiirdGYyIf
gkl81BLh3F9MuBTkNzGNcCL0QgbTHcTKwMYgnhzEwMB6I7CEm4HFDykEvR0kFZ/iMJ3cZ10A99R+
0RlcFuHQqMR8Vy/KAGxKpSYVSYbGE7CmZWL4xjD+7HiixRERqRlQTLlMrNg4LirpqjVXSXTGtE/5
kn7cH7snQ7P+f6Gjl7wncmlX+BmJtkczryeJG+SOaPLYRdEU7ELXP+nJWKgDOxqdlX8qyfrrbE+4
CRw6Z2HJHyLtaTxOojrOLrIds9SfNB1SFb2RLjrZMyOJPukU9J7FXTfrQ/rKf+QZ449LOl1YrNSE
bxsYy1fxgqaLjz06z30psj1yNZ2xDO0I97+3ExgR0bLYl16dpSGqTNdBxEbs5HxR0piFPn149BSS
CnDahAogkpoODtB08VPzfO2AVcS09t1AGHoQ6sEnkeZpASxZ1q4K+v5z5hdlgc33glvJG94stxXm
wRh+4FRE3bq9eUE8uxPuUuRT3WwKBnRK4qm8IKVSwAM0EZk/YvkQtIRNvmyznq1u2/jXzAAAWsIW
0qW7cIVrZnyRRLqtjbHkYoIrFR8z9tayLIgfEzcxMpAnTNioWF0nudomdb5HM6N4SQv/tQntIJst
elbFw4amQPHALFVM9+Kcdins0Chpi6dbOmqfmW1NmYftWOGFGBGl4EU3BmIHTTHYEbTVQ0M6EDi4
cstemEUXZn700jXTk3+mzfhCZoJxLdx/fYbla5ehrAY7Yg+kGz1uH7YIpd4TBgb32NK3tVZIFbFj
1pxrPrxKBANVsAuFR+1koJ8VJVf8FwzjmX6BxuLju0Az9wt092DvAYJlrTeVydzWKPPAlM69HOry
LEmWEKNh2VTacqfaHydqpRThUsHtMzS2DT6zs5TIiMage9VcBbew4eNoQN0ldD6+zwZ6WScK+M10
GwYJcp4TSEQhJL/NHVglWx7IE1xxcDQoWBmOEEPAKNC/nOWrbuHa7s97dCtgMvzrLlb7DGqT5ZaD
EoAtoKOHlnZItjMcatii6FN8h4T3AkUwvgh2bAxZiQ1GMBpj6LCHQOxvcSq/6ilqOl4i3d/gb6hg
9XD/w3MWS6g0YJ0g+RGXAbEqWxj/Ajtad+v+rdjvjTiBEzPpnCp5PFvDep0IWZKjiUQdjKhkq4BP
Q7YbBbtmfPaYZWXWieDVd2zKF+ww+RXCKcS8BJuXHfFs+wnsFrMXS6rEFnoY0P5GfRzE81jTpHvW
12iAdjacZXfm7kozZehHy4D8FO4ftNS66adPeoIZCgAre04Lb8eUqStKbtGIUcMviSoN0yKF+I/l
9HbskLv2p3h/perzB36Gqxljnkmgx/qeXtd7ro0kkSzgeVARCcKc/UemZ1kW2q9Dj7OQK3rvfHB+
Q0McGwUxC+rkMQUcph2Uz3YJysjbVbyxFG+YeMLBz4L58Pzvbx8B2DHw1HVVRl0tb46emXbV75t1
xDDnWR2ilG6URERsRSRfPsESSNybiOn6STO2kvIUzYC9MpH8JpbC7HZuvKGP6/bpTBs9GLOOTU4r
JE6N952CGtb5OQgd/DZit4OIUwZosfyo6j/BemlQOJ4zfRZerQkeBwu/wKcru7YuG1sAguLzEYw2
fHaW5HkNs4f7aQ0KzngUsZO1JFPi9DNzDuS6JYlXrFMnQ1YVrg/E5gBykK7+A+auXIogxgntybts
nBbdess+5gbjEllAuRW5RitQyliaUBF6iTv0/Cnu7zxlwlj32RX5eZAG99Sh0ahVt8V+M8NupXHl
sklrY9emRAV8nAn24sTj/1aKyCzR3m3EXIB0h3CX7EyXRSwUjt1cSuJ2IWBUoQgAjCrcS+Hi/nDy
85tyMjg/BQCpznLYZxaeAnslbeIfCXFX5LaPoH5mCuY9DXhsWrN++r9tYZw592k8RhiW56VlAZKB
3X3y85Pr7lhkWojSJfdmvFsc6Omb0PY35vtyyvpx0GNZu5Y6HDkcu52YPXVdsPxo4IT71Auqmhht
q8vRpkp0HNKPWGLjfmHa3mdzE6NykbF86jj2uZSZrGGuRl2yVn8xmweWP4r2476csdZdUl31NmpX
pR/gr9mzpYZ/ykmqO3xDypfs7xKpXzJnKlc7aJBrp7rzs6THfl4og2hNazbT0ttKqSOBJrJaAH3b
J0ukUmj3s9svpyW7Mkt7N/IpGG5DYNewDeO2FzLK0cUx1NA1YhS12fYIxziYi3GU8Ndqq6ca96Zy
3EYS0mSbFcLjA7QZ+jG/0muVMioESFi7Hpr3QnNX9dpjpaV3FihyoBSvXn6xFgNb44xHcQKA8yf4
zSmevH5sGBC+iZtk9ihx9R1WDrdmDeKCrsknSyazgQgugnYcbzLxk4bbQP95NY249eiPYVne8uc3
mTrdwq8lIl+KCMq1Z/4ELPlvq7jw58NcnPWicAWfyRNMdFrNCBFJ7jUnYodaMlPs47jliTVOtVei
fiDzuDY6GSGn+42lDJPG6KXYS2iBfIoi4d90qqbe7p9lUoumB/x44M/0dd5Mv1xoT03A1v9oyG7l
vXnMXNk9h3KjFZeGnC7NLSRJmD2WDncwuTzmFqwM7pvM87uP12JwmOwJkBecNyk94Ib2NglwjSpl
Nksgi5Ns+XWDoM+hnxhvpePROfdCuL4qZhvbdky5FmqARm/wVM0ObGVa7WeHqHswkScDGD5aNF+9
jDMF83+CnBds7pSXMc6CxWDi2TqlexQFhFGq5ClAOdDD/hEI2BeEatmXYiTnvYdVLa6RP2mo/nx0
2P9WwfiZOX3tvjtmUsXfkmulU5E0UXTJVf8eIrJRqxCsfaCP7+r+45Z5VAItnlcWk1TQ9nwA6rHS
DUfCC/4bIcEAHFU1F0YZl+5yI24S85SngTvSLRxrTzJAq47WlfuKgq5KYFtvONC2oVM2HfIIL2JP
/YdLYK2+YvH/wNaTCHlkCd7yp1e5l3aD3EF47mpculCfQHTxzYr0sfxFYC+ozS77jMx/cR7qhO41
07WEToX6cbbhMCJqDnaN0V63FVICooq5aSnJHDqkiAQ9SiFPHsiQiUwUBU25GYgeXzAG9xKzpOXO
XAb//2W1a3/oeC6kDt5ji/IjGtcCxTSFtuL3y1ai+3Y6/nVKXg+JIxak/0zMWHD0z9Ga1p/ldd74
Rc5DVf2YsBXGgC7aZLpeF/EKcNXEMK+0fohYFO4StYYYRp+dCV2XCbIt8WiNCvOc4tUx92Kl2ChW
WReEXnu5x64rPeDVqVX8gLKRTDKLF/PkBRUJozRwJX/rrkGJbeb/LRpErbK0cUzC9AwZoqKtibG+
/ko7c9hkaCDgu2AqAI4qTQLUmN8iBa3eHMOHApCtP+Jf+ayvAeX0Uo3HsXKUG3pjWs+XZMKkrjPM
IH+KssthTqFIJb2IO1guBb2A8pcQlmPKXkIRQlh18wUy4+cLK6Hup+c92urA+bMekwEj2ppefe8K
/aBpyKblL/TuADJv4oIs290tfhD6nVwfLs9S1GWWgS+mV5QrxMzUQL5O7cg/k0eg/4yCRFTBZ8Xm
UtyQSlmEJ53gJxczloBKC+uWx+x5fIRMvX8xVMmOPz9DLOKdQVtfxDLEU/8nSNauFFYrwVeFwYr9
qSC0kJtIUoCUGqOFtiJo/1mDiWn1e4ENdjMqQf8xHi1Rg5mjQNJUlOhusIN2vU1fvtWDDXE1lKO3
vWCrnu5I21z61saLV7RkFRWeS7j1BHAGSsKzRsIDZEjqPP5QZrrY4FII1MN+D0+GPQdUWPi7L+Sn
lOrpjuYnf3dRo0Z4lPVKNgoCAcuKRF6Oj8tmIVCUzCfsQRC8PVx230H/kDCDrZPgd68DO68xYtZd
E4NN6ILZ6K4SJSuoLeGiThQP536iI1txmbJwUaMN5I7HpdY2/jHGt+SkA9vVdBwA9R6ThrTXP6gm
fd/y8dzEmX3jFbk70AUbA+tbnZ4xXWN626xSBVmF0xa3RGu0rB0qrGr0bCSgKKJZbqxc/6l97bzn
+K910u1iCexxtYea7Gs5mWvgpIEnTxP4eLJPkyUmoK/7cSo0qPKvLlUJgrPrZaafCbTuRmwur67d
lk3vFQdFLH67xsX5DDlTtCkCXyrH8/GnpEyHopl3g5BDd1iNTuzpzUBgoLTq83cE69YGubB288mP
c3+eu25y12Jusu2fapXwoI5Huut5O4bUjwvecPeCd1zw4ZArQo3ltksjd+Y2ebbU94iuayPhveuy
nevfykJabsvqjAxLF9W7vz4NBp5XkXw7ipOvdlF6yxSpCtuMhRP5ZQvQXSbFBiYva9LmIlmO0DiV
b4FJxmsYr15DITYRYfMzf2giIYIuG5Cf9/VoqbXwehrBMtXFVjyJ0xs0N+BNtuPtys8zdz6P9sla
Sf2czOInG9KdhTywISufOKGeXaztNZ4XRjgR4WhpeaSSNWUEAg0iJWxisEggqWDYzynF+8Vkr7O1
OLX3XBwtF1MWQLXM7McsKxeYRg0AR8svK2wEJ2J1sXrleBruSfdqh840l3JS5hplnfHTncr+Riyc
V7E4YMeI0sLpZoDqtZoNFNj4sTpcD8r/dlB0kNJGt9C36jVImLWPGak+jFTwdJ7JTB95cuoLkCrr
fqkfqY9HwOwWO7x6sGh2to7tvVNX3UVPaX5m3s/DDdrD0kfricjxNywgMm/9p0CARlSvj7eb7OzJ
4VJbS/P760VGBPuMlbjLyThbMiZPvrodyhfVHAoLwzMq64ssE3mVYf4GeP8B8Sp+C4PeNop/h69J
aJSh0fB881NrYWAGnERdr/amiGO/AKSpSChJGZA1+VZ2W5hLS2HBtYr1J9jyiX/dlp7MxtqcWaFb
dRcy5rbTMwnnjNjAWz0yFzamOR7kOFmWhpBioblJIVaVHsOIYIsbRqmP3fcBsPf7RjqsgSSu8mHO
I952fEtkDgv3M+Vj9MvAuODZLQUi0xTMSe1mw/86N7OeN5dIA90IrhuaNgk0tmsIEUtRFmuqdcb5
sH6nFBql7RvYojI+CKQWeOXIhvDfGpBYDvQpqRQ8Z9SDfJodU8FjQhpSfvZLqK+0JCJ2pIZVGolT
0XxmMWlIzFWXLEO4fyevpsliAM6l9cvCYNJldo1SvruStwPJG81+eE6U+tWHjso/zeydK3qX3nRE
vOeWEA2TtPmd6FBMRYDOudEbTceTmK6Asjf+QOBLWoD5DHIdwoTcP1ZisGOe7w0IFEaPtSw5nf5X
XXjwTptulsHe/q+n8lhfu9LR6LLkkwIHoIeX6tQP0X2AoQamC7OTZ7LtWUvcfKfP/Kw/4WsXPSHB
5ip+5tCR7kIdk41Y1orOCFOQCTjOvJo+fVYGl34Pk0WXr+bzO9UIrSent2u9GcYakQ1RWaJHSXgl
dQfrRzRetj2m0vezDnrchPcXtgI7HkjGv0rKe0hl5uRkeX/uUc6UnoScW6KtbPnQT+vziG2xqfrz
1+coon/etje5RIY7zhW8i2bUcPt6PmKfvZpVici7DShr7rleMUi6EECPp2lc0xhStoR1GGZubbsz
gmBPmntkqfGXidhyu0f9NRQkdLOrXigihxlOozmy4kJlZazzw4mC6JB6b9hMImWeJLS/gEZk9D/5
np7Je6bVJ91uHEDLOl7Fz4V62b03heosBOsT+1eHxn7QMR7CRbx+5CLaidrJTCfw4lxCCF+oezrS
5hnk1diNMV3646C41EKARCwiIo9Hw7hRyLGwQwJmqYUQ/nQ6Jx9vNFUmk0HGEnplEtwECKvw5h8s
iwTxkzAfYrY1qAU5NbvNg9beBc/cvnfTKG+IPpMcZ7JIDrMSipzCZFLGGCQYd1lVPSvyJBAxc7CW
t7ZvVIe98Tu9U9HDhgq+H7kVMCgP3BV1gbV30SFqymvC9Ng6udoxG49sKBBsuqnP/EtQ3dTiaZGn
UIalz/YbZdfuHWLC/uLNCYXMPx2I3Uqf/9TxPn/6h5x2iSiiYf9dSpY6jcd5JG+j/heLPlWdgiAZ
n366X2aTQSeTtPrKxdUgcxSxRnDokMdlHWpPezX8Mat1ncEANcbGDzMn7JCzAjVeyNFrMl1/nBKi
DYyuObwg00LaZy434vaQlARobhnh0mDTyjPiKcjKkOX/uQpuPsBELbRbQvv52MaSUjPMLtGYZCWC
sNS/GdaFj9h+xfvMigAD2u5bbSFaoCfL6iqREXSxHo7YqjDU4wO0x6L3A46zznoePhWM4NFmACk+
28ibB38RrKdAH1EPJOGHmSkHnLp23+SEk/OTXcONvNwiTYLZ6vAtUFEjvCgDP1lccBtKBMjAnARM
eXT9h9g39qF6kviunAN3J612tw6hUOM+ErY/tsSZlsJasMMKR0ppbv7dQ+G9ZalIYEbjr31k+AMn
kqRyWNu+sRW45sxodhgQ48McOQAs2WPpzolUlPiFniDjQFrGuQ/VNm1PSwbm6ZeZx4EyG3jNDwM+
9iKzUYi2fTboMKtnZ6VKlWPZBNZRjKY2dI93nnZslY7ApspQh/Y9B7d8i3LZPo9hjx+xSGdWHzmj
EoehPvT238RyYf+4IJT19KkNcpiOBZihBvv/wRgmEMgnCnrGMerLQNqEBJjLe4VLoPJC10zrIuK9
zS1NSZ8dwuUixoB5jv5AYNlwkkajPty3XmZAblc4gPq+kzL9K/VAEcF+V5306Jsz0qWwVeTfwDII
lAsD5rJBMr/VOX5cEUQKcqfWtrnoHY6kZRgSxcQp/Fm3LDwnnZcB4yMca/LHUefWZi41dKNTukOd
dPNUsddMxOGO5lXeR0vQoCt7A3kUPnEXiSL85Jhb3q5sRQQJGL3eSP5H2cnC3NQ0d6DPZ65aKCys
IQapDjLSmisPQ3vsuq0mHMZeHKFB7fTRCGFH0WLhbHif/ds1WJ5BeJpqelQRyCR9/eKmq4XnyCjo
ieR1mlMlwlRE8bY8R2NALRulelyqJesjLVYAc1wvIEhOZKofLBnzNyTZ8Cf06jxYwhL1UCAUiSTn
5vr/2u5sA1kpU567j7MwMwInmGv9Dh9Drm1p7HhJiNdnvSezW0//TF98Rs0FGWCBiQ03hz9+/IEA
IWLRM4zK8YeHD7KGlZ46dJDxtrmvR35Tw2D5muEezm7+Kw5Z1ibaMBpmdM9RDl3MxmE41/V9XiFA
i5DGAkb3hkL+iib34xCBjkIIykEDvroXncBNRhMVByBp68Hr2+TpWWE5TgK5/EXLLsLMAv2UY3EF
OdmxCnp3pYlDXH4llFnNxB2AwbgaE1MiTcmXz++EIvnJbg/mPjo4p0PkIbKfasBTcKk2AbF4VXn2
Mf0gF38YaAtLePJz1tK59pN1ezASjMq/P0YLkkejxm1NpuO4lKFe4/aXaw7t0o26s3gnsGZlCsy+
d/kx3AoL+a8+nh8Xq0IF6iOLdun9a2lPIgYVMjvhVcmTLvFQLMj/NoJHLkWQ+BAVCBiXWVNBDcXa
ut+YmlEcTbQMvLx9SAZ2KyI8uexgIjmjEqPsxMn0KHQzwtPwp0vLTfph+2MY+QYCmZuWxIECVi00
Z9CGjRxF4EAqX2LzLF8b0d+Sky95Wv1OUF6g4P7fBSeNeRBMsQsmDh2EeD5zMAMGeOgb+sxxOSc+
9kmJFHH/U52MH1b2lgUJRLCR0QPqD69f+G3sewdCBm6DX80JuP0CTu2/ldJM9xGNr6twFOctlG8F
qlP+YtRpuk9ADa92/WEffnxIWk7Xk/+I5Cys6me+oEqYV50GEcfAliOqrfZZ/lT/HvThiMMmh8I4
hUGMAqEEhhMSbItyXEFbmkHQSgW30FkxpjovdTCyGnDPP9arDZAHtWjubtGcjcaAXP8GiUWVVpd9
YxXw2zjUhiiNTJEAIm3RwozfIHaXJPJsLTuJSkUpzllsYeWHhyU59Y7tRSiA1XRwf9X65LOtfAJi
Dwqv0RzvjmUyKbS0Y+y4/3GXI+tzii8eymeBuSceAUBgz0a5p0r4fIeQKHcMHHWyqLMBBGXAaYYF
wjQQdZOJZ3KfS+lrMgMc4buFdM1s/qc3pOIuEjHiVUQC+JRuTnHj0q+04OZpDTSi2u1FRwrQJkr2
ob8nDsIxXU7egNzwEJgtaZ1e/tgUBDUNfuCAkr9mtRh1bBHoAZAHfmbBf7NwFRHyJrgDx3DCAN5L
Pp5n0VXKpD5aYLcaX+OVR7gzUiC3359U6OJ6JVdVs1Xl9oNCWJcLwy3E58w3SvznPIcdmLnWC4IA
5tTSHIRbws5+F2TQUlfFPr8gCADEkxE2yfO/IT9KI/z1GCJcYRKoo+oy5I4MNWXPD4VukcT+zTMt
3WB/li8JPJJ9gWLYfTJuGlTG4of+qINmTiJglDhJdpF4NEvHMiBgV7VlPqlW/XFs61ASlp0FhaVy
WWSqmUhqwKEtlOY10fjYAb6twiKcCLcb5oYeea/sc/2FG84PmJTkOldC5uIjNNP+JdP64e1yixUW
eJ220kgTd4ZYg6nV219QZnEaB/qfiXN35a7JEhCsRMIfMnAnAXnu5m324rxQnbjrmAKTOCcbTyPI
ZObuTUrXBrebU30X5tewMtgBcu0Ec5xFGXQZMU8FGlXefOYGpTPfZXZff/Eh8J7HJoXFIlOWtVP7
14mBSxFyNuydyjA2rof/ID8Sc1/9iWPFL+GtgbczDKd03kqglYHyFufUo0aNQMPXsXRwo3E5imiY
f6vHnMZwLMSJ1PfS2gCgVCVElTSJwtAiDQm7hmMHPF9p6OKYsdFIm4hB4A9yn2TzXDRccT8kU+T3
u3ZG6difBs9dQ4QJU2kznW9T0ZylYb9fHsLf0S8sTLuDvg8rBQLjKrigTdIlxcZ+vhgcaqeQoZh1
VCCDh9yL5sAbIe/ZWZ86ZPinhWK+Vx9MGu/9hmKFMNYaDXJhoq72BAOKU8Fc7txbontlZb2TyRb5
fPAqvBclNigYxSeXHwhgm/0eowjOSTMPdj0DVeiHczao72/lOrJ2nC4nKw5svR50KlkOmS95Jt+k
xTq7YVWAbE1ttOQHyS/x++ja4sqSdtQ/BHcL1e4kI2Nb4eWCCONC5qQRS9FiCihMSV3DpX6klwK3
OgosOwm2RPZSZPxNRQv3T7JFP1I7xpBLcxjpZyIN3fYLvwCjSWydC+CeVijFIrwvuaFNTb6vSPL4
nWVzQo3YPqeRBX2ZstA8nPUkQmDFfJKBTA0ceUAx7iGZzLO1DseL4fFBXvGP18Nf8elUyEah37WA
/inop+S9EQ7XhBuB0YvI4PFt2yIwmYwSk16Sni0COVPXGPjN9NFyoG0UeRQb8VPIB3wFv7hEu1To
HxZqPlE8mk9U0ib1AVfHtIohjFjgmgJPoWD3/gBLOE6iBYBlkeE8jv8LtOB4hqXA6iTXXuD33iQT
RFcAgBXnSKJLnYPmmiPnqyIPGmEnXVImZx2V37cWGwlZkDfpQVZvdjWdlmchV82mz/Uqh5Ic55Rc
pkzqjO0iPfsy++eR7s7SsNbr82XdKBXUqk/d0V97DeiFoGQnJ+ZyuhfvU2usPIhId3x6UyJ8cORl
tTkWRlq9WquDBq4M+aJN74oJX7jMGbtGY1pV5JWgy1zRjbXxMjIWwL4qJef3TSvj4miBr0/mdqlE
Rjo9WyFxpWkl6+GPOXxxWHX9hGOhtEF3xafsPp16dtOCYrtxAiFg/noM4kvCZJEprlwXqQNMP0cT
/tyu0R3nrL+Iz3ko/JiC6w/FG5wcVqDIYZm2WnljlQzjkI42D17EgI/+zvYcwDNfYsCTHp2PtyQd
n6PBAgMHCJBrRJ/gTtU97FnvYmFCuck3zBhiC9mpJon8HShzjpMAtNoy7/hmn4n3aq47M9DenjmB
vxiqPJz+RN4Ui8xIAc+Y7GwwwdcPgco0M1Fk7d8BZsHRbYF+Pk9CTNhnOmeY5iDOFLm7hol8Fw5m
aa23Yt9wXnybC8fGZtFO5qVBDtphcQ2DILzPcHI07/O+G4v2IbMDL74r2ACU/p6SMWLn4Il9Zi2K
VFpHT0mHSzIj5okkQ6r8mAgeTCKtGLzo8yNtImrEDW4TyHMHpssbnILdKE3CbsjCILiI/sDigDmO
HOUshRE3H7XCj60HAGck7NUBKlP8W476/HVFYkVz4uluI31i65Q9PYT431j7YI/dZ5zj5Ma/11kK
UTgp8A08zT4uCO2c3YzTNKWVWh3zCqtL2U049hpbx9AXB6pHppM2QoM8hqqr+z9+414VmMWntHEw
Y2nzkm2jG8y6MlKs5QiyMhM6vJgXKGxNV106/XqyXPX2sTl/2UmoPTgonf7O8FIs99jaiG7KmlIk
XpCI0QF4waqczQwCfnN2p4LMqYuNe15KoL1G5hBLY0X7I+Siyh7IMv1oNNbwWcTGvR8s6VPKR1WJ
Pvski17zUcYvhAcoLU6TBY7Cw01ckP7fJLelUzRgMHQBq4s298OobZHVmBX5RZi0NMZaFP6MVBJU
+nFb2oKa/UWv5Eamt+IBeYbr6KHA1UNpvPl1nSP+K5/y0HVrsB8reLxcfD214Xcs+gO4Kt+C8BYf
eFEpGc2bGEaoh2tlmwqW5EYyum64sorh+Wn0kZ/e1K4lHOTCQvYVa35delviTK6FP9upNDzHOUnn
g6Sld+bsyY/ya3HrLqX+PFItu2caKfaECLI5zhYtgdowT667O2/Ez++awJld9x+iNFPJ6zJMa9JR
pj/gKohh2QHhnJFdeePyPXV1/BFk0fvmLIsYcxkUjzgKp7wToanKf/eWkYVN+vhzhr+bsM/a/8SY
3g3W3KRrKHJQQAdm47z6dTEfv2aYvJNVo4WXhfOZ014eVQd7RreI0+7wnZWgdvBz/MZK8cVUe8K8
wMWPENStxH7Om96268IJ8Mr+Ppw6Jx8mA7kn3A5V9jzVYh1WkIHcKG+H62XJ5nG6Jl5rfbXBaaU2
zkTOX306lMMRpOkOXo3Yr/ZPxagWLCnhWg91dd2+xDQXcnKVl8NTaBQVOG78ybj60JPFpK4638YA
6tTCrMxDTtJnUGYqw2ESHEJjBFn2oZ/xqgQ0dUM9md2O+6fxaOYqw98p1jMk7C22eUH8Qmar7Via
QjiWfYHJstzT1CpEeH5hz4yO8qoGM9inLnNcBW8sIQipBbScOA3swDg29JXvWXjQSziVAFS954Yo
h3469BKZn6isXb4HKBEq1ogDraSo3hqW8QZPPUpNYKtGu3e+XlCLTOVu8WWPzCLJK+2Ma9E0fKXT
JZq9s1oxdJHFblH+By96Y9XC3FhB2S2v8OfZ++S0v6kmWeuf0t9m/C7/rSNrBUSdMDD9GZbsEWbL
u1sYdY5QVaGFBIWFNWSmJaUDfUSh97Rse+NvUNEG29VnKb2iBUCdxgDRs4P5j0jz4/kkXxR2MX6L
HlO0X4IEQE3ItHlESLc44qS4DeS4fUaYXzBXIdjY9978sTEify2lSOOsbRd9u5Bg2WM7q4HjTiAa
qBMtzIWF7E3v9cO9Nc/3VYOX1arNI0wJYEHR0Ra5/CyxRjrXYmoXUFCZznRv8icYgSC1oHJzbK7R
efEYvioGkoa9KlQhFCAaOm2PprFpR0So7xDV7nW7PC/OSgpIdpCZMTnEfHAZAwijQImCbw9aUEWo
9wWQ3oIi6oWoivJxClLzueMTrJ2YxEeNjILWgn/ywR57sSFTCSIGuaWgmKINIOPg1/ftR3kV9XYr
vOL9QwySYPlLeVpXgcUiXPehr5Pus2l/nzODjHcL5Q1tkovIOlu58AryvJxIlk+ZSSwvh47S2g0w
jptFjRb8L5zi1DvTEmWDs3LY7QnKQGheqZVw2lA2yLGZp4kqUYyOOV5WXBrm2PUll7uISRv4ycpG
4rndXb1TQB6mRVlY+sVkl3MeiISKWL+ENzDQqDUZG0AtASf1hACbEak+PvNUP0CNfP/ucvRk2u7c
LmF0DRsmv2F0+maZZ423Wbyzk3HzzAVyjIOgkQD0NJtV3YCR6lA2jfTt5vGhvWQhgAYpsEk0wgrF
XZk5rh0MiVjm3NZ6EUQkCL+T6PE3+4RQK15drWgNsJxH5ynyhGCrrl/jaax9LpKVH370IYGQKjpr
vKvU76Xe/NJUIyR/C6bwWl5ovv6O8c5IIyPpg8+FoZmv/3gKe1NYKCw0M87LpUb3NJMmueDrYenu
8g783CLtZxMkr04RY2eGFi5hmPwHbwD0MoWq2Sz/BEvJYgg3HEDSiGfLgjV8p48SIizR1kvZISLT
zgCyF1fcSUoPxCUHBd7MafxJ3E68l+5lvr+tDQWvqu8BandT2f7g4tKo5a7HYDRvELUdbN2ajPw3
2J4y5M17f2vMNUSTLucn8qKjwFULr0AvPMrHbLff5osREkzYEu7W0XNDvpPPvMHh05GZM9H0a9d5
4g+ROwhAMFL8qHYARC5twH9wJHjIOuSc0Kdo1Oysym9XNOdvmkXef5IJiNg07oAOTE3bTIh/i5le
38QiivHHrPug5t2Dpj39W7UV+uHO2j6TBA2dr3jNO7KxtbjUOnLmpg91Vkg8bgZ2EvUxT0bGQtSU
DIDBEsDwp4lyGItZ2u5ej2ebvRbomyUYZuVoQ6IdzrEOElYturN2oadGGVjoG2ud7WANf9LLc8t4
4ugZ+81PulMcEvfm4ggFcy9ofgqKJ9CoB2B4QGwBQTdpqvZIjFLR7aIXapB30CEkAkQA8CNg9XHY
j+ZT1aqk/L1SRLTVaEnpKiH0gdA+DWP2EWswZ2QdBs0bS94otIg320dg2kzyN2Ts/4yYnrprZeVk
nYK1NIAjACpV1mseqzuYB09sdy0sTatw3IxwJj2c0I0eXsMcx8GiRXAQ52iIzO/JgO4fhvwjtQHV
RIEeqTlZGAGqvqNK3tXCdCu5nkKxWKBh6IzjgpQnrtX0hKA98fWQAnWCM5gw9lQFHjt+InE7kCHv
FsuVRYNpq7kK9yMdqP1AmkmiPGOgXlSSbaATegP4pL2z5VwaXPFsf6PmW9MIh/fSnBiSWDQyJtCD
PQfDkjhnVUWtHSI8Fv4PE1TrM4G2UPXRUf+dcZ1f3syG3zkxjqXV04QDsAZyIXCZ3cJwMFA52nV+
Px4ATG4HCSwxtiLoOY18DwXIVRL5Xi5KuHQgdI4cnsJft7Nzrn/ExNWrIgYKa8O5KWZO9G/LfnKV
1t4bTdEMQ7e3v/2CXbphL/WQx7JFoWG+xKDEM7OGSLygYxsBJxqDe0g+Kptq/Q6PhD9NfRadeesn
WxDiATx0ifuYf6BYmCkePDC4mxezfvsEuQ2uheniVGGULFRuUZTONSzPdWxiie2Nh6shBoIO/Fpd
4Kf/Dp95ZDd7Gpc2xODWQvKmBSrxzr94/887Bhq7u9l95N+3RvOC40PFQTROrk2v+uxdgi5hRxm3
33XpRKDBSlKnGqRdtkObgA3z5ZIq0F4jQQxJuahH4DTgYIg5kipSgyxY0DqbMocatYljrbKG9Wp8
CiXemuRy607l8tk9iIKC5fAe6DupLDVKP4OnUMeGp0029DQ0gMASv+U2SeCNq9FFOR62msbZj+qR
Bubu6bCM1EbbTtcMc7mC6dyFgtH3MeLFTU/ZU0l9TgIDMmP4phAIL+AN52TlWjbW958OMetEoDuu
IDTsGi8sMymf8hCYDOHiUe998wE2MOIf4l36ngEF2qBt1wpceFMmpcbNZVdsKaybxraBl9isNVro
493C3Z4P8AhcB1Jeh8uUknzQOHvvRToqZ1MrRv/Ubm13rPLZf3wGC88u2iMnNo/CRel4/hjCW+bU
JJoalb1vqMQHTBmOFubsM9e5Ti42RvEtr/zosHpdISLcucGmyi7Se4JoIy+Nno5jJoVHzL8vabNd
9XorZ9nXHMolFM3DvkYv7pMIigO54N4ayomdPaWQJ9mgD9d1qjdAYdQTYW3+Xj0N8EwldBU3Aglu
T7HMKyl2jucW867RfrHJP20AxBhO0LeOA8KleRSYkaVs5HgRUGd9NYoZXM7EiyOW0aph5xsJd7VB
unlwVOBDilAlhN1G4fqhWPH97kjWFX/2oILCCtHfrtRk8vTL2wp+OSKkY84aYmlYmRj9stw5MIja
aB9Nq1VHDlO5qZ8lCvC/EnTpEwtJGQPcrjGGLKioBRn44SRF00CAL1aoPOc67UhYggpzoj+KAVEj
92WL8E/iNKXgL7J1PeyBN2qJ8e55RA/Ud1+2uw8HOeyRMxI6+22LCNRmuTopPOrivPpsfUJHHVB1
2iYVOroFkAcPxfEqo6jxWwVQSV8hf5WN89GFF6rS2f3yRNnFR0Pqnt+vn88GAEPNAbQs72I4o09M
4eknvWSUV6Wl4V67DD+uySMTvY1NlkiCk0sA24t/Ci/CzkBq3GtsaK5mOuBJOdCpJvdQdWE4bAdm
lGuaTsIIJNscU1ZfFjJrN/g4MRQV2xYkglHryExS913cLI/FHnLq15XoiH2MyMRb3msheYGGbVUw
B+SeNptrsOpv2xvFLS4zK1dKFXqTy1kEgfd3Df3hgpngXRgJ8kW5VubwGuhuoiFob1jViKGfvZTp
15nLdSIoeVPBX0MtewGoa90q7zlRN8/ukQpArxaTv8l+jwmPQSBT8f9YowJFGEtvd70R+2f8JeZm
D61x/RjK0gLnxH1SzwdEJ/RjElVRM/G7ANvWgNQZli3ZXoywNhZ3BoWgOmeEp1C2t8pubc9XpQkF
fjGKyTxAqLoXEX2YY5ZZuPcgrJxB5k/C+wpPxIgy/v9uyWg+FmyEwnXkbkJRjLXHy1c5N+jQwkXj
2NfgTNWdiFLzqdVAp6pwwcqJpxVStnRwmkqg0yt81m3xM+hbbXl0AM9aqDaJtJ+6s0xKZ426DwCS
xvL7oxw1TkVgXHAXRU5nUi/Dxej+Ms8gD4lUrLqhTaf5y7M0n5y658qK8yzXzL52EWLxRRfVUsE/
LXib6rB5OEhvvW+E6jSl5gUbP3zkigSJM/EvKcbM9xOLgmtLGDfbF+xuej2zRSzc+tpGlkPvUGpw
VV2dun8Z1iKoN9cjdRn5RaCYktoPqY7h5jT0E/H/SKdiPqF/PY3VFOzxisJdX+rRemXUmHEx7lQp
AKKlp+XkYbXeULNEbCj8G/itnSjYfCkrqG5tFdtONKIbn3uqN+kh8G/5dBpqJp3ubr9vFTdApwml
M8ApCm4RBd2tgfQfR2VxyIOCMP8vIaXgeR0BcGdxDr3jSc2uMfzKYQ0kd/TAOfN6BSLvekPvjS01
oDQr8Obxdr++EFcKZKim5hV+WwQgQBhisXFWiGJbLxnDzEZonWZk2VZ1QlIg/plam+mRSgHfuhRr
4kbitAWEpDWdhFziDAK56ZqdenUf1aIh57etJKGj6n8LnK6CIu8d+2zsi1hiwNvIb6wALThe/Y8U
XoRd9+bGPGBOlEw6WDGGf5FzvVFWmHU+gjatDNR09c0aeo5cDQKVqXm1q9MIw3rV8DQjCdDzQEEZ
z1FZD34cPr6Wg5faSkDPdrVt5xDjilfODDxAKWBVhkF7uhqxQv/EksgurUAeGnT4NpmedDzWfi8E
jTAQJHpJpykh6zEV6iwJMpN4WKWvUT2stikvyi/yfY5RuIPi5OUbtW1OIeCIwHYzpz/p4QTZMn57
aFY4X506BY8dOKL5f6Jfs0Q6JW6Ctqdd9dxPJyjYBSKmzXbcyWCHwzy/MS7ujqCPxaygnMhYiZ/4
8dmdM77NYNC8va2dOyNJ7xRsH2kzPbsvoDxBcgRL/rEfGja9lOn5FRvBj7NFDYiXeo7VBXoySldj
a3AHrD+wSNReFTCyw5lEPpwEUfyNjy6/ccfNDvwa3trAXkrU51V/ZI+VJPOyOTvTE7Ww1H+q1vLO
HxxniuU20s7RRWrcu+fZVxoOJI/dB92PDr9Soou8NbhlHba2QJyyEsf1/hxq0HRqZ0n9g2pJhel2
9D0d7Nr/biLrHyFKFPAufXX6UJmY3EWGwHdS3iWUekicX0oj3fRrjhUrrhmOlX3k8J5vtywyNNPx
GxzFtepM1m3YpVP1AcmzB1FF1AnEL7vABja5RXCsJldN7JDgEpmw2jDixiS2PA12wD0bsKDFhMz+
oOrevSHjx2+E2aXhoNLr742yCiAXKDrVBK+bdu2tQ2nHi9N8s94RDyXFc7DgygCCkSpcVQTQzu31
RegUTNzRr7n0/q0JrwWLZdw705lvMMygkgYUViHD2mIidRPN+05Hc9Yr+Svw9W8kXTY+V4Y2OEmX
09oqGPpNLT7vINgbJCyVLOZki0QSHy+liReRFFTez7Uud5Fa2/PadF96btPAJuP68lhfaDw6e3Pr
7EnMXjHloy4mQisnHOpn/icjD/RJo+tRFsJyyJ+WTnM9Z2NjvxE7CgvnqtbLqkAai9JAjvBg2LqB
TTgYlnMVsYxntKLxoeYggkljSl/bJKJsVIi08aCYrU7lowWyTy0rAjxmA94DMYEVM7jzW2S4YAXA
rV99E161NlbPKc12hbjMUhU+WN/jzWgnDeo24LP2B9JEisKmvaRCTH3DpcP5GlkT3zsTDaSfdnKt
ZyqDa7IjSQrQ6lSO938NZXIZCalbBob+xJrDyP/2gO1Re8c99BhiQ4QIJhVxkjPQJZ/NOIJFc4Ee
3JHxUVa9LKa9qNp5XiNuXexethB404uHTTKi3MsnvpYdhCUqMG+19m3wKsNrNeFUMGM4TKfUNADR
vjrUxTTjjYfQUpU8yjAwevGbs5fkGRTWOoxP0ai7vFrFwH2Hd39HmO+UGx7Te0dyymMX4nkH3Wll
tQszehMDPDbQkonv5OAs/Uq2OveRO6cuoqjSwwxaId6G07qGJlAFs2I/Hj381JaUwpfT2dA58EbO
bXJEypy3eCs0k3tfD7x1dqv6nJQnAplaSS7B9mISK99OFUkFzd/Q9faOS/SRdO7gO3xyqD0big4B
1O7CtNxkOp5JxE/21QN4ufp3Yl2M8XTD1nO/O5xmM7nnccyYvPE847XEEDBhPRxlUTjzRHal1RNX
QAqvzOIi18gIgURXY1GvhHXkapuValwPfghCJzUbsnBYmdBTn0WWccIvdqGG6eyOyzv+r1/5CGh0
POxm/7KCL7ZFhSeAp2AHG7Ecb9vAwM5H9apW6zFDiPDXWIDLWfGBiT1Ph64MJKDi6tQ0pOK2jHa0
rwH2AVsL9JVYw5K6VWH37kMuKOhMWVrpCbR2MFDToEgVnfYgY3VKbWyKGuCpBsW2ATJz1DCi8vnf
f9uBpixYG71FeYfBV4ol8WClOWHTbGEh/T6rn7rKJQZeIvZhFbRg0kPDKRLWblq9Kz897QLvjFMC
PVvWC0/vBkKPIh3yDCb6vdwQxMBKhB6ZoA9WKkJvRv6ldvJdpIcue9mRaFYqlYTPiLCtqoqQ8zGf
KeCglBIXYMa5EjyDa0ORgtfsWiBv5RN/V47C9Fvp3BMXSYsc5BrH6afdSoQTOEJ+jPN8GuEZSeSP
6wHB4lBknkS9gGEve65jhhUrAo8KEVGNQmFm5UYRv1S38r29nO9Zk75iw1VeEsazmF1uzfwk5Mqi
vw72YSB7VPXLfWam8aXpMxCpzmQ5qcsWCrg984gozBva906AbdbkFk7+rvjd8CS3r0Bqa9OldQkU
K4FmJgOx7wJyNzX2pdHDaX+xZ5H22ay6ZJPpAonRckqvbBSBLW2IZDTi8PkuqBHQi25qSXSMoN5M
HE2lKvu0ejBqfXZE3NP3YRXTlHJIMaoyyOU11U+jlFJ5wAQsOi1TmGHp9+LlcALeLZcdOLckTUZB
0egAP3xJphlGh1guqs/jnF9l5Ve+BSXAcDbqQBj3PzdKZ1nOeplhaoeqIMrLxz50SY2/45wKyHN2
MH5tJSt+TDK29zDZesLRCCnCwW8vzyyZAIldcTFhPmTaq66GjY0CJ3ECcb0RLUlM1nDrt9KQ9q0t
ZOcOGxMhkp6c7ew0NFiBRCpNOFobVuUeMWmlTaWfktVxZWbuv3be1F47p+WaOwZkibOID2+1xpUF
MZIc1+dEIwK/9efbulbWKqhOpszs06DZLz4t89trihGOt82RXcu0QotUTAjilYm7LDhW2QN7MSrP
QRx6aXhoG/w+eec6essRsij+XkaEph3kQO3mnc3b00eykohX5CgXJFpkTwXZ3sYn5uhXWxrhn+Xo
8l1QM3XX81lRqFjb14SEbgBIx+OlP3orJO89dZAFtnwzUO8HcjW1E6gxXru/A9IazOJDkDQ/apvd
EW+T/L+Dz6vUAzbY5jS9NUPpP8M6obqDLQkcljNo2W7o1im+XrrJ96Yj3T4Pd0Q9gbXuCyg7ON2q
DR36NJcRNJ96fHgXovMsg3u5Eaie710BHcwsf331g0GEiLFM/hPFN9lNKatvYYg6GM2+JdolPPHH
xEC6GLPqR7r5cAO8U6oCgt9OSmwVYF2efFEZ6VRRyRYbKs68549KVxcJpQVK+xoR00ClFqIijGdu
fKwizo7OFYZcVEkEcCkAH+xxx9l/TlpnwjrVoMp69OgCwap6ebINlcY5zaabUsafhNZwWvpzCDZ5
YcZ2+B7nDTQo4b2Rj7RKaFzWvGC/id89+iIvVg1E2dJT3uVsVzPng04GHSbzCGMtno1OR30McLtl
15mbQj8nEnUsugo+rA6jIx6LzULqj2eid5zJoGjwHsQEjewtC0BsJDr0kColBmvdC4hYJIwoeO8B
4s4cgFtGmwJAidEwbBr48kFAbL0ksapUnykwK8E7m7bfahgfVO09bbeWPfCGgvgrCzdiB0nOtyEI
ayV2z8JOgGJAT/ZbzleRoo6LYcub5aBuez3CNPsLsoImwrncXMvefouhb7ZUx8hK+pExBQWYjYS8
JqdZSJ5wsOqaNPIQYhJj5wrpRRsdmS6+GhuAvxYu+Q/gEcz2sG8GYeIx9u+3b4vYzeex7hIk+aqK
uDF+jDdzaTYnVX1PEdwDnqJVNRXmff+pgeIcdvfWql+lYIRFMVsHtUL2HjArztBTbSxz9XZbw17p
c2XrRczQ3JsKkqYizjAbBpuVWDv1mDznknM/XWMvDMCgF1nHj3kdWfjE66C8NjhTeX/4dGU1suLr
mp/YIQaupapVGRlEQjFFOSx5nFusNSLgS40wKsNKBuYGHsqXpBoJoAovxgBfWjF/IuwxzN0roJdA
JFCcaquWhe3EQeobIX4G7gETbpZJsETrbBYuOLi60pM97mldGa2utrnB2ekR48IEZnepMDmzh2H2
Q0K3tulQvkgnA/Mbk+IrWDfoWplxlGjxQVbNJVX2Tg4mLCGHlHNZNtHl7E1fztYdn/Jdq3iaqBAZ
vnXykkuLjWm8LQYdohLLkVEQ77vb2TZYi3Bo67aSDFwJ2XOUrAKRrgVv7lUv8VQQPgNFKlvTA0/4
hCGB/EmDrIgo0ASllBzqsDAoGVv+umRD5P/4wladDHcx6+vLLjDxupQtD+Xtqv7EqiiFvO0AFhT9
fLAnvQPM+/Y3gGIXbUmH6Gme11NJctd18fl1hGtVRkWgFemAh3uvIMZrxmZgDV7JDOGF9mFdO0Yn
UWd98DceaZUvHtj4gr220p3hBdoMi2Cb9UoybD9OLRX2AcL92RY+iwa9LHO34Vmgy1QiIaBbO3q9
rX1oj3FhhZTiqMwcB3ZqSqZqXvwf9nfWQRACBQodNnYJ8w/rnmYtIzyvsi6SH/nYRLajoQrqd2AR
20GmpWDfaBy4tFR0X2mipAXaZIntuhUIaWrpJ0jJnqpTNeQ6foAI+VRcrAvHsHQDuSZMoHRI6QxE
qUDtZGWYuAAaUnaVtzsIIS/pXXIkAtggv0JYE3R96WKE3Wo22b20RGkrCILhb9wJg4KP5szpVoPQ
/eudozhUq4NvCVFYkij3EV83Lz++fEkrTO7alX0/oX/xGAP9acQZVG9q0Wmj/YWeHtPz6Q8o33Af
0jdUNAmUsccSQKowo8/iqPRF3DqxzMJDIL+3TSfi9GL0CsxI1Z47+naW4qxgKexuski3Z65nuHIh
uH4Jo7gYElUCeVkD4gW4c3FruiqAxjBHSKc05/J8dNdvPPQvTwlAoj+h34UaJCak2vP7T3Y4hXzC
5fX4GDD294K+siUnc+jHMf1/YnjzGZEFg0oIkjrAVpRVBq+lQXHe9fXXhe/WBrXPuz+Ga9b6G2e7
/GkdAwQ6Ha+zlFwB8jJ0DRpFTw+nOlTKhUsc2SFgENtgBg9AdRRvqEZput34bcp6k+lVHj+TTwZL
gF1AA2W59b2WBvQLCIT2HuVTFVH2Cye5odD0mckoV17b6afIAJMTwL1ZORTXGbyD1H2QEB33v++4
+tlE/LX2/IQw2TWBlXH+UFuxSQMLUjVEga0R5jwjeUGMozcOGamHMbNOySAvX7VoXxfWd4XEjBCA
o3Cysb4ZUxA93PlxpeII0eWuGu0Dwe2nPY4k8rn/d4nPJ5LvusgPSj84Xxu+GZG9bUubBjKa2xaD
beYbJ/k8pLkY/+t9TtcsU1Hm1nt0NQTWyhHQkHuaIV1AdnMrpY0Ffo2ApA0jkNbCMikN2fXp//Ly
Zl3ejf0CGN2bLpwa0i7rcE6iK8wsmKF2H4MX2xAZNjX0uzwWgmMBMP1jlqPASunACxsBuOHQd7Vl
q667o3314Dpzr8+jS51JuYDMYzaXbWadDOhnlo8AO8PFVQLP2VMJPeWzTNVK5qquEYRhGT6yrFmi
SHv4rpESDOkUCuwtTPBRFiJJlHi5AioXxhXhzncnB9vrAmtV+UWwZCzdqfAyD61Tvog+F6uJw16v
p01Yt19LFfWFoaZ5fNptm2YVL+g+GZPIT862M+kqDGCwkffwXg6YlF22On0pFm/OL8VHuy+w2qMZ
E50DUzBv+3HSnl+v0qI8QG80LkeW6z4s2tF9Qgk7ABiMZBdidYqVVves5EWsBpN8FYfShJwEIJ2t
d++pQF1tdNdZ3LYCShkO7Xoh0feBTYrai1OY3jmyIZrE8/2cqxxK4Wm8qAoCeXHX6xu5W485F7Ri
A9biClKdemp0g8lkGNTKWLn93eRFIqlkWuDtgDnKcNO9NqDuUXG3eDKIxs1caAMj7JrS1Q4zKVV4
Fke8mRtzQhNXc7i4PKisYO7KU32CEUK8QDquFqGTbToGNpLplURnDgbzFNuM6H8v0LaVqiZYX6jT
ktejQ4z17SrO7vomjwiKyKa0sAUQfrvvEz3Mupo+gsYsZjqo/iBP4AWnhVobSTAbTfv+ujD/rLJ7
FgRrD7Tc0cI4YtZfCHCBQ7N4hiTp1Ee6NqUf281IrS/TGlI8bcCa1LL7FTqYTDmlmtJKjnGdsuOe
7ZFT/EqwexqSLCb++/pgU0kDqdVfRK22++x6usGBDiwO5nLHUTSp9BG5HTCmuWxYFG2LtpwEYHfG
5+HgqvJX9oCZSQCQSOSMDl1rmD++hpw6pC6vulcRYTS5eIynaatq4UcTgD/+WZqltXDE/ujoM9gG
BB6DmZi9wmJtaUXxxehDXpAwxwQMcQ9k48hsSZe5UiwrGGtVDipv3zgTNkPOAevdwLc3YH7gGyyS
rl+7FPh3/pAAZeqAZlfNZhyRY+vGDlyXxK6NLXy3PBpI1yyJmIOdsjzgHV9MXTmI9g1+R9k6g4bW
a26LC0NwxpYn3KQ7fT6KBc4yh6/yw+AP841fByUIQY5XKKq8P6ZijuWMUxsjDUWj9Jfy/cXRnsTZ
cfqIEGOPrp7REAaBpiHKi7m3L0qkWnxmvNWCa4rgjMunjP3c70P7TzCs9/spy5UhHhJnaStLN3pP
soliquuZsPXzwTjPnR7e4vfOVobOH7i6kwvyD87HT0sVSC3Hh0gu+iEnxZF4iR1ad+dh6OY6wDzt
PoBiU6n7qgI8NFeHrKbMITFHn3anVrQ3VoBa/cYcC2ZUIGmYpIflYuBNPkNcy5cVA6lNRLHlvMG+
h14uq94vykpHBow3dJGCwqbN4y74fLjGVTcAdt+VpI+WLE8nbsdfYzl3Lw7riIfwiUO/XzPqJlGY
vNEIjmRJDcfuUv2e3FRYP6bqkDD9LlhFY0yZPknK5zr75skjzDCR2nMkrf39XfIzTGSlVd0U+RKP
guHOAS65yBvSS25lFg2TvOHX5wOCcE7E10iiCjxwVHkOmoLnbpc8CPzgB1gtc9S/2R08yS80/VJZ
DKNBZs0QKNDlmzSC0WxFtI8EjszLbaFnksMU2D0oGsFRz7BynlrrrmfxTmAJglG2gsvLJkJXtdST
twr+S+qZp+gZ4L08sRrLGpieBwmipkdDKABTKLUEhMwL2NCJ3me4STp/gsTCxoZDI2UgkqP1+jw4
6bZnYnVYsBNwVyALS3D61l0E82lgkxEsE0aKQOraV7U2jj4w1FVJHn+a9n5aWdewXERJf+PQMS8a
kGMmoaSE971LYWHdGHucTvAKUTOyVFmwNQgsxXMYjYlzwpYi/EDapyw6EJ7wcVBwgCLf3ERFVn5X
RDGg0dTFfwzGntfwtg+wVHd4+4yx+TeTDIFvHBqGOdWVPfkJSFWJonEma1pYBPsm+q5jgQwPH5Qj
JJzp9dOSuNTEeXEXHPGyc7ZEbyPPRnN4pQmnWSrpYnQ+0urnUnteCd2KNOUSsaln6rtKzFg+V0LV
voSU4WONwJUEwsVKmEsniSpHtU5KqH33MYTR35Okhgi39xnbgmRjZ5MsqnJ4bEixdLKX8ZrVlFS+
fG6DURAtCu1iymIFlGHcifrkRf0kBCyGNJE72GG+980p2uFEt3URbbjftBOpHG7X7Y97U2e/mWK+
yrixB43Ette1yN7XMzSLf+70qV7QjFar0g7vjdBd2RKGUjLwgZijVh1ZEB16jgJzcZVYADFIFn34
gjXcwEVTRgDYPagPZ8kHZlB8zUG8EM/CvpYLkhw+DkkcTrf0jvY6AvTLw31aLS4Az+uWQtH5VWVP
l7c+TXDpSyBvA/5BU47vg5yI7YPg1d8kiEKCqM3vbCIHUGTmiPWrFPr0XbbJm8vypzgTw984+Z4C
FgjSCQ+kWDnDlhYlOfhu9gXqaUppCvKCRzo1a9p68mLcv0GY6A0OPF0m480qAet383Q6+sCSepzE
4AYAtv3ORDW1LN7yTCOe9T4pepFBMgY2f0lCDK9So1UrkfD71gFVW6rJnd/Ix1cqUWbjrEybCO+m
idovX11qv6a8+YXSiXbDl/U3IWOuwQCBn01BU9vlzHRSd6uKsmVQpBAWlKmls3qBkB67MjEaNbl5
Fn5YfnPc8UXobqsqsebXbGDWxD1bvq2x4QF8LXI6GQAtgyaP9w4sUFvJvTdZ4m1w4m9MeFdXobQa
d0McN1mLqsPaD21S89fRI3gBQ57CkOx4Zud3OJV2kI1/rlsxV68XTRTuyQi9ayywxL6NJqQi5yXy
umWATcw0dJLqvYGVyod4/y66iGun9ACtNBDiVBbvBkukxYDwOXFpAt2gexC8ERDJcI0H5iPp32+A
H3ToWxfILg2vMFATECsXksdg6wVZYks5TQUQMaziRM+ZumXBKB2+3krvDQa9E/d6DFQ9NzdRQ3Ii
I95twJsEfj6fcz2J79/SUQCwQCcOCDpIVSxeses4RXE0yKZLXOv+ROAL0Y2/P7thyD3F4dq3em+7
N5fjZSA5KugLlDckhMUjCdHGpBksTDLoFpyd72vGiX0KS0bybB4/v7B6UWFS/VeacOU100JI4Tt+
Kimoyi9dhUywrECwG79FxS14TqVxicUfMTiYo5CkFxtt8LikJme1oYXW79LkKJXV/bsr4yK53jee
cJ0VOA2Di8SsAtyt/6RFX4C81hBxXaxpxPyrvuOFq/WVEVh4d5a7gVOevHbut+eV671hoImT4MAW
Oq/y+XIM4d4PNY04etni92SMGHhDXF9pYc4dPIvUdhDSmh3NO0Q8S41jPsVgYkhWGH2YbqXDZAbG
EpRPB4lhio6GZOz25AD/ikWtZO2cMpr/VXafUlQezWyqMIr6WsuTl47bs9fIGHbXMnRnCp7ouvmv
7WRAkCyMf7rLie60kU8cIYRupMtBigeRluj/dIoOxl620HZHMjuI8LrDnKHxLPU3tACPtQhfKaAO
BisVUVqcJQshSd9H1t5C+4aq2LlSbBavXetqjIEPR9z/IUTnayOVR3IdOd5zp6zVlQ5GzBL5YdxO
VGy/yICRBAhSXDxpHWV/ifE0hcAWHIOqWK6UBElib97b6GonU0oX0+Aj+qQpXOl1HQUQOBj7kQpJ
mR4vLD5WCrRhctPKMRcjQcY2G/THy2EmI8JbXtyW/7+clM6FKytOLYYzoSHvB3oH73YaFXhccZEb
Ka/nekucYhz//hqRcTgp2qlPL60EtJ9ISeaxNd84Hhpixum/m569nHq0hLz7xJhYvkwk/eP45/Q7
vf/0PAQI+QRl+B8liGAtBz1ccC+fSH4ex1ci5GntoFEUc0mS/dZXICAK7wc+/YHtBN8ilCwmEScM
o2oi/6Kow6LhB0tWAb2WQZMnwkPtOKtSxsRlCQ9xlz8cF9dpjKAYMEi+YoeCIGDuXthB+AJxQZYo
fwkyC+JQgVQyr5KFmB/cVKdp745j7DCPHFc3+bV+/IF0iULhFOycsQclB9KbfqAGj2dQp7q//3z4
4PA5PjYl5SPyPgdsfFqZLrjzBFXQ4rDhm/I2GiUMQGKr/eeHPT+g5WAUrfi7bsbqnK64arQe/VC3
jLsfLih5Z2WGg7rJyKZHkofBdrG0qllHGXXeZR03KQFKzVVj/et9ZgGN2dpyq90eM9HGBiZ69VJ1
ksBjpNmAO/nYNMd7aIcs3f3rONu4h2L0VI0mhaXTX7Bq6bLiHpMlpnD+P72sczpQxYvqAy+7QHOW
UD+KmF52NrtzPhtWbesgFRao5jBEN9UXu9rK/DkXD3AP8J8xBe65fxjscwx9Qi6NU1n9sWcooDeI
B+e7oxaSpwvDkdolXETYVM/LYQ7BarYVe0BTxlGF3ogy2M+J5T3EuY/GfakqOKBRnFrDBARooQ/8
cSnxMUoPITLcZW62HdF9ymzEBpUuxlPQECWaOWW/LsOaP9H27btTpxzV1KDQ794/ijT0guRZKVX3
M+PKxo5pGR2kvlRFpuouSD7pwAw/WvwsrMma1wpdZcHhD9ppn1hX5VD+/j3MK6ucC1FAocJhWLOx
5njxfd0E3t82FbGvHe2R/gnXbik9mTRVbFI14PQE8DnGHJu6pf5Q/6gZiocxnOj0MrgGRuepfJg0
jhSrHADfIs6cmuW4Ty3LaI3rTusCIWGxYvh+1vDrE+GwsNVzAnlJ7NQHOgFLhT0DhRoSBamJhKPU
22ble1W7j8eZWeOlzxHJL9VSMzqDEPOc2kndZSs+PYFibpwrDi8VMhkOAL/1X8j4jrv/mg0CBG6c
Sfwr0JvbJlDXhg8XSdOQaA12Ukd5kAW0+Dlb3Eg2HkEwbiUo3kDU3ePfzIpmLb/YO87BQDrWDH/z
hcUuyE9sxJKWlgjARrM1PfRJjxrBchVoGJ8mwtedfB6uE8jigM29+Sbk9BQKbxFlYVwzrpnWB7pO
j3nqqgNTK0BgRTHgmXybBNCd7MhmNSasPiEHwBT7BpwP9U4FjbbMVJzx2bSVcWw3iHSqRGdqgiau
cFncmd7IfCzmqNh5Jpe5ffVAwVr2gF1qflrzdvvR/elQXPxppyAyAMHjDeNA9NkjR/h7JARcVPKp
Yk9fFR1PA6TyxRjBoLbqiol219b61vO96j0a5EwQvovphjF+nhycvd639A84CSa7NMIyK9l2bpSI
Oo6wx8Jjnn7ao9eu4KxvRVP27c9xHAZ8zBnSiiloog28fjAvGlGyvfwSYUN7GVoPk47F0EEWED7i
MAum8GKPcQYFcWQXEwO97Vm3GEBVINP1GcfB3f3rYQ9Ukwd6qnh3g3ymg+7yt5JLKeJdDKOiV1l+
KGX8pTcSbOSeNqX+JfH/yBGAR3yJE10vuC4ZuNM0WCqEDEOufZRHy0+U4JNiCpuVlpbg27KNTmdm
TYCyMhUOm+dTF78AXuWyYD1CNOKDP8XC8Awupg7Ueiztzosdkgplwc98x+yiKMJcdnUr25ff2loA
pIzGZek76pxmS6QsJuTE6szINke7WW0MS2Ka1tQMi7dEwrXqZ2g8Sg6W2LK4IsQuvWs4T0CbfyfW
IuNCF8QoS5TnH5C4dR9zKjphv7aoUxXWrFUWpkWVd1JpPlfjh5r+xPPFPYl2ZQoBIXxmmuKO5Du6
dTH2eOVcZUPnImVAoe10L61yGS1YJJ0xf2L2xVonyYXMi4bN++Jwd+lTPCqddYlFHhS6ozZUjh8z
PKHz+vmihvtwB0s6wkyQ0SCF8nBmw7IvT/iXdbJjn29oj3bB2EgQcsi+0gXiw4h8ywtSFESSXiU2
z3aYCwX6DxM+6+5CiQGXOCt6HnqTR/R5BZ8rUcZ73GPr5r9OhQOp6etTV7vBS0LX1DlwspJRTyV0
woAl5h7l+SRrn4T77g9KesXE8tB6f6C+fTuXaKeYPyMwMkGc2BYY8pXyuCOGBmpih2Som8ABOmoM
OniO0us11DvgBfhv5acOJMP9D6q2BfGJLe3XhY9a8275nqB9fJLR5ohLQ7dvCLLp9iUa00gGzAEc
K7u9y7Yf7rsleh6xGZ4WmryDoZwuXibQxkHgmS5a8hIQbyH8m5tD0+xDaj50+vp7P44LM5/gfw/V
LVUKYaoFH+u18sdKMz6Ll7qoAyAnjNVO7i04PDvTUR7X5VROjifavYG6m6o71g1NGB4YwtKa4nBC
UK8dFGbhEdGOheGm7JnPlPnMGKnlBXUwiF6LW7DYS0gsRRyglYAokcIPooboAqJwtryiv7U5A6sX
TVD8v5xR8xC1feHPo5NBXJmAWs70RoPYgRgiCZ5sLo+9mlkecq9qUHsiBjgsxXEIzZLHfmZ7xA0O
DFs62stULe6fsT5nkl/BJtJMlMskk2CY4xpQkt9gRfePERu93ja56q56jmNqfFlr3CGTGhl+VWVI
L8Y+r5G+D0O4WwVExDi1l12CKxeJGV3qBKIecuCIZRJMUP11cC4HaoR5WUQgocWWmHTCBS4aZd+A
0zyHv460VJ/ALTVkyZ1e+KFEMv/XjZ7CAYWBOGM2eN/MQ75TGvGbsrUm5gZT90VTKC62AOeCUNEB
CM7IYvSI3n2irR+4sSH24jqFmgSTEHoEWdYNJhEIEpKojjRNHZTvspwOZc2HjvWK2rAFZJiKyTr6
lqt1+VL0JBki0ox1no24FgAVEwerF1NNaP9cw6LzForgimYwV3SSQBckUjWa5nLRMBpK4F3bfIkl
x11bDRGZ8D8NKNv3XOZnxixZtbMegxP4GPJCwSB6Y4Eek9D70v7T7F4rouSk3USbSxIhYeo2XMe+
ArZvcQ5yASZWx8NtNOkvokWBTzuX0b9qYxRR6kS+XBp61DrEy6RrVGocHNSPAjykpNH57kSFcU3p
2aUICnl7yyFogXuLmlbELP6C3iQHA3pdwMQkj8iE+iSFrIuK7bJpVEg9SmlFt6O5eGm+MemMxkmG
xxUhbODF5W2spIEYhIQ53rjMrtsPkirUFHbRN/FYvaYlhpNsdFF1nQ3Aa1gPtLdILGGfi10zlbos
iHMkLgYAXK2yun+hrn9SUCWMluXY3rAh76k5AhvK3foORN0IakSRyDmKg7PmNzzznhCAGFccvbca
GZny0zFbm8uyOJCLO2T/DXBqXvm9WH1df7guFwoJe0j+qofXnkxdXmV+kZ5JmUBCdWWoYYRJatzB
TLII4CL4ctya+fRlQZ4XG8DIEXdGqfFOjS0d1LwQ5hXe8yWm1oAVfErqbJU/4g2+uRxtUh3hF3Qz
i2QDCWEnModfmcGc9k9dl+QjZO9fQfiLtoGY0JI732lOEW+FxhdMXynEswEtZq8ASnj4/yw/b/ed
FE/urfAu5XcWp3knqJE4tqI9zzHEFWHStop/IIhfi2LW06IVT2tMd2RoPOxwh0MI5KPNeG6J6sk3
7wk4ZkTB2Os5yP/VDWcwWfI4dpg3/M8sPJJAU5bpi/f1jDfKeMEHx00s9vjSkEMCykZUj1M87z+O
L1pAiIIlEiWoilIX5sZAyW13zKqDufVE8wBZ0wFpA8ldnoW7WYD4Ujx+QPx7oS/RSd5FQ9NkJaH7
tYypxEuNbueph+1M6zHz9zeascSD2oFD+Z1M200cvfB3fm9pUv6usnrxkGHpAgSnkXQDI3/wCHRK
WCWKVRcq/tcmkoXz8dAD+yoXa0I2kZLSqHQA0DY9FHaoXUo245R3QqLI24vhElC0nnT70JqpU13u
WN2ElFj22lHwdz/NKdI7NTb0yyVTR5W0iIDSWDwBLGbxyWgFGhx3PdPj4UyPO1+ZoAxD/pMwqH08
5vwRlSqZKv0KBpQ4MH/QchPH8DOt0kxjHOnkd3BtHQ/+ULL3X7qK8dpo3aPjid/QYbqaNGTbDfGx
VBpe9ss173W9C+yN5OfXSUpvKT3l8E7ggdu3wPzt8Pn7NbziGWYTexD4DTReYA3QuQjirTo79Ym8
HGvLTA7+IXTnFLpDvCK5qhJvO/oc6BgzczB0Ko12QRXReNwuSnU2gTv8uxCXWNCkLD/8t8lxjKFt
qgWuY9S8prbaaLKHq6XSxHMwJMM6Meb7EIt6A9pACmXEG/eUNPBldng7zN0/y+ZE1d83YOKe+GbQ
6674nW/MIF6LlA3LaE/DVJcFu9knlSEfTPTa7E8ktqtbps6vUd8okfA9oHX0ARbK3yNrf8mWJZKg
gRVVe0DbCqmVNWGP/tq4KsfJqHftTDnLfNu+Uh7I2w+zBhdI2FHcNq4dAY67QFT13KX6Qk8c5bfR
9ewCm19ICQaF8Yx3pzoebCHwbj2Cme6/kt0z0nz7+MFG/KsTKHIa+3J3qQVQ3btmLqylHv2uHbiW
D2och1ux9ZlqjrI9O2EboDJhZpZtkYgra9DO20xICWXQDEMfAglvUnXekFLbDJ5wQoxMSiSqRMHS
E1lP4Ql8lDgsaur1dUhNnGRle0tkCWXrzBay2dq6WDbJ/jKt9hshuOTWaVoLwYJjtFTeOpbekhMo
9g3vRSYfj9tZjxtnvICSx/RqwGKHEfmE/Ok27EvEplHkxcpgiP6z7R2O13kw/FG28mj+lp96NY4i
pBOX3AOgt0CE7hLfwjNO8G/ZhufKm/exkgGFSkelWQ0QwIqVFUVjyhqH8w/bB18s6n5t8NlGh0I8
jt5bGjUOM+tUFAo5hX5cFTwNo+l67esUARUBnz6M02IBqj1tRkaTqP06fLZrFE08yivNOXZ1uK6o
pnC6Sr+s/WLy8W3rmif9ERTQPwcMqPwmPQa34IxFJPbTAvuIHigHhapZWh90zZJOPtkuopzUhfai
HpvXqQEAcNcPjs1k16Hmr0CYYnbCcVEpnqynSjLBiBchdydykKWZV+uiUSV4nO/y1P5AkKfV4adD
gAnU+XTGlpyUM0QpIIht0FwEJ4PvgUXAnxB5VEHfkPouxBySYMzIs8bqAhJ2OetXZ1DMRhF1f295
M9SAa3sO6YlAiNUQUEPDpm95aI34V5HlpGt+B3G6OosWD8c3EpQv1hZWY54JIG+11qoS9qrMrdIv
xhgemCGIhztU76JYDdtw4cav9pTf3q37Eq+5pS8SORVb1iRavvhpGTzQcaMErrwXPz2+JifxVHKl
cLJwzeLkIg/MLtjsVMijn9c6o6fx9H6Di7Xtleb1DnLZIwrGV+TZ+w1IlzKyjwxY/z5xCRiyeqLb
cXA0Koo2N9V89xsRGGZjJkeSZW7UMzqbaKnKLaXXWqYoqnEFZNiFX3BsUAzkjJkdFRoONjofhC15
7N66E8lUUYz6xIQSAWAlE+YMJaYJDZXXG2onZEFPT1jp0fQKh5lRr34VHuVR5Xf1hRbxwqLATFO/
ZEWlhNoDEMZHYWkm/y4u1kqgoFtfujcsA9jO0pmi5bocEfPrQyT8noX4gNtFshpu5K/wOKr3ZfSj
w4w3dzXnD9Uz6Ih/YvrUQyMWdT/sAiVhi2d4pCZYwzAvuIA5/rhejg5WkbUrC4D3svIQ90cFTD/6
y5x6AWXYdR5/VY1O0sO5o3TosKQbtjd73Kj46cxX89wVF+XesyKm0vORa7xG2xBwRQAEBA2mHEUr
hE1SwmtP2N5I4VSlO0RNudD/WBIIWeDSXwHdHYYVE9iUnk+rMcZ9UxjiUZ4ZEHUSse+eCBsLH69f
qWL1p4GiGZZANwEDHcP09Nh83T2IPJp2o+O6Ol5HUeYypYiNT7aQS3xhV8Acfisv7ezeWGKUxB8n
IWLN4O3kQakdnFtYIMUDrruON0/BFReXPZzzXTrUeCMW6/6n2HKZ1P82D7QAZiJ6eAaZ0kywKTOr
3L7QARI7LjF55f/nbzIKPQtmz2bzpUXwCZp7k5P9P46nSX47jctwhNG1x2lxUgxuF0m9hOvt4VY6
I1PI/DesraJwMdy6Rd1TBJKBKEtj6Y4FUkWJRTiYxHGJP5JYRt4U3Ng+LNpWMgKeL/GspPJYGNAu
3kBtXSczwxs/8kc4C77I0n53KQXK2+FQOC8WsyBJMTzo6hOzskt/Glssdlei3GT19ZHmZ3/L2ym9
mD03VuDl0BQKjCw2E/YiDsS+aFrcT6C1pONmH29dxIdqV5bPLxX8qwKGxat0Xe3tW5hPC7wSXE4Z
XcLXzMFUbriaYWFMYR6enXWZsrRlWCwXG2sc/8y/2bw9sBi9kD2OP3nbWgL6348lf9MAK+cnSeP+
JuY1azdodG0978KouV2M31DDpozcNIrtNOP51HZ2C1W+SD6TkBIc1eNsbh9t/saXDQYx6+yN1mtS
lBFodt8HLoVHd4ic3OhhSb/Z4jgfm7tX8FLnlo3EcpS8dqXmUBmnfgpm8xCOoqElM4lt0DKejePw
W37OtgFqAXLvQAvPGADwlK+gujXEl08af0iCUBDEB2TROzRDY/HtXEpa+yEO8H6qM5UN/tDYjiwu
FBQ49JUVpascBZneXcGoO0ImqSTz6wMSxuaGfP4q2zklw2vBvMgAV2KZ/DTVk/JZmbBOuWTa82hH
SY7jvUHVlHsJ+GeBpvWwU8e2gMNDmpj0IKGT7zPe+GFpa5GfGUfaEsXF8NdJCblvMfi0D1GYVCbr
xcOYmhTrpdYCbUbxGh8xK4LeFALo/qEAok/oBHC3PskFEaWwsgZSGAE1piklFcmI6tROM1YxrdPj
tgaVzslihJndQnSzQjD+qZWZeZWlz0kyqX98jhaF6MFkLBHAZ4lSO4xLN5HwOrfr52iGxn1h0d5M
POOGGsLP6Yx8AFDoUJK2fx27UGaCMN7GUsU33x9m+VNjg/zl0jN0KMCPRteaZMCLSRbJH6/0IQDY
FIp6pnDFQk0PyoAlJ3lbinOrxJi/LAiPFUI2AO9on+7+biiEwMQ2rWXyrCBJMHgWPQAg9TaGF9EE
aqqf8R1avui3nkVQBOkxnTUA33CHCMRJMjOfgOUeZoONEKgBD1BuS7B5rpSg82ccnvhSTgmGagw0
xHfPETEvmwXwsyu9usKHuNb/CxNqC07cIx1jZpL4HOicjzqGnLl7/pD1QSZa8Qq4sTOyq3jdYnzs
ZSMs3C5hKkn17fo5UnHuKEvDfSHJ8kHBHV7YGedI7N8XgCHmy4cJNDGK3T29bSD7FQAIkyIUS9jF
sRAQm4ldxhDJj4+EHS/XQpYG/EeCzzcSz7Z3KwhN6WRDWTNr/AeNK5LzEalg0iIElE/y3gVpBJ+q
uitNGnci1VHjfdlvjezEBtxAKw8w7q9fZz+jKrC5QHbjfdUksMcuubWaajMQlock8eAymiFxKzMa
MkGVdmbDpspx0Jb6WiTODTBIEaBMAmUGRjn8AH1XufXSjjOi9jAEodALdcSrPySntcZM6KtGGfMf
mwbTDtR9qGFEoMBEMSUj0FKzcZVFF51luCotQTPp5WIXewM12h1OTl45YrIpBWtH4LjvlhUb0DgZ
iUZyYN9aT9FNQUWVWz0gqTjfcstSKOZq6OmesTEoUI2tf5OYoczcccW/VHRNQ+Vi60HkeJhMRfVz
KcfWcSy5CcgmsrxcGIDM1JObN9K0fzQRDm9lnZttni05noUfWR82/BhM/v5073hLYMj2CIBrnokA
CRS2xFxamA2Mtk4vt08eqy46sCyoTIlW0JlM/zBbhvsQJP2IxizBMHgdv6yopy0yL81SyNDpuuy1
HMj8mJZspHWGypcegkbiffa1Ytp9Hn11XS+YBtTDpOv8gshLE/eEOrYoUDliMfqIvvT69YHAkN5L
twtS72Bjy269CLUAgKD3Vc6iOkxCVjCt7cjTs11TV4q9x/QYx6zCJ3rTNu6AudZAZIoP8z1sg/hl
BEDFircce9XP115Ksb4yGExAgvoLTwfKRVzF2Heth05NLb62TbBCcN2MoQgTrVdCA3WeUvh5FdV6
DbQe43Lrs7KWHGX0mfzaBI+dOcu810xBxB/fqXqcgDyySKjPp6aU5IhYwUHcF0cAvIkjmLJ4UcJ4
TuKFsqbh6EMSjqOpeY2NDMW43Db3BKA8FNgoSEr8I8ETzrIv5F873IfHesO2dGGzlk2z9xtbExu4
BEV4rdk8Msy9xD8EV9TPjntZEwi/LSjdj1+AGPdbVJavbXfIaV7bs1SnSCxLr/kepjLQzy28zc6g
Ui4IeJ7WgN/axf3ugtMrVCNsmuCV8zsk66CHK39Pbe1ABNzSuPHoeMJ2VEnWmjYzQROsSSMSYQ+9
hTO8vvX44W1Yy997I5kHssEwaaj68MXJtOMCdv8OTCTm1v8imIR7Pp5h6KXBd2aZNFGSgWFF5S74
UAKhZABdJpYCxUItR/TBugkdiYqa/qLjhgXDzNDTaWjIz6ePzN1VyqENm/CtQDVdY/J1pL6KcDaQ
kgHIarM0iTOKKmceUgNrE7rqzlyOKDFaruXRuD+42cBETSlUVQwsUZBw0x3XaRVhOllAhSU7djpY
Ktvl+iIhabpNdVhi3Uxf9o9PQrOSaqx8CwU1Rzs4yM59agmHBwNGGge05GI6T0WPchy+/YlneLeE
vcAg7Sn3qdXCthbWiTMGhkib6TRJ6k8iTwOPIjwyZaxaBWAfCMteW2MdLmVkWfmpvyAOvUqP+gov
b+xGxifxqPakDSgzPWi01neyLwVyE/u8eg4DEBIthUrNq2MaJrBDzKWMK79VNV2pauNxWW70nSuV
RcWC8jgVZaGiCgh5dMtiaQQcDZ+4sWzx87q4uqBSmRrbomQuSewzwDKsaNGhnv4PpoKF1PVpcL7I
aePorU6GZn0hHaKz9vz+z2sjbXo8sIgkAvdG/pRzskJJFpZvNBAFpK42Ju+ILoYMpOQYXRgxIKjM
UmMxgF3PZT5Ukt0shmA8pMTmHmrkSyK/0vl3/fpL5T+0KPvaXqxjQQ1YwM+UYqlcXY0V2Z8HcM23
Sov171OHL1izx22B8qyUvE1C5j5AC5nIJ/MxFt8EC4vQHTpI4Y+dIhKOqZM/DH5M+VRCmMLcpY1S
MMkHt2VkLuEDhvPaGDrfO+U6fjK+UMeryF9GT1a06/n9UmfxpMDfZMfZQU+c5eH145ulmNd+3BXI
2hjgqOrXvlGx2VGNObYTGEaiJEFqJzx7b0toRsE59iwbYj6vtQiAz4ph625QKiyJP4Hs/v+7ING/
z+xvDa1AIctIQoGzkMRUNPk4kP+UGzYquXDMnZiYHlCs4iivBCNeZZI3E7TiQ5jkAzcOdFFdwbEJ
eMSsxcazEDoyTMd719uNqCV2M9VFwBiqEJ7iJuKDRexgvMv6qbJMSsNpQ03Cjz/J3K4AK+xT5saG
s+AJxNaH5mSeNO2p3/WeLPyISEDz1iv+JkMQ6SJOL0/RnUfEG422vpF/6dL+hlkt6FrK2liA/2e6
WRjOh1vAaQ/i3DOkTdyA++RE16zh7n055TH1ClMPVBT7zgR41ZiLFVcBdle9+xouLrOE1rYnPbex
AATa/85G8KPmCC/urgV9rMM8CnQXE84Dpo9/G1pKoyaUtxrCDM2nT5ZzKFm4SifxA9FveugkUYTk
+cfHoI/fXr4RW4J10Ogy2aidhwRkAUUYq5hrsiQp5+YrLl1LBvnDCPp+Lv2h+LQ14B0kjL0gaoJI
lsWqlVoIe7mkJtnuWyerKmzC/EZ/F0BFii3gCYsTSOmu8NEDRRpbC4968j6Cel1Mc6dI++Fl3Ceh
NKwDUe59zJCGDXYDbqFEWDOzbLuGNi+xxOOVP5ePoJLmoVbkExcI1XN8sUpNdPKg7vt7EQ6mmYaW
pmO9Q3UUeoIG+UvzygzD3k7FNOg4R/Ld8nYL30b4gJ5vsjcWHhvlFuZ163IO//Ramo+vFjB0dyNB
oBl488u7GxRoYqmFYiYehgctNsFyvbJ+RQ6MQ4/66FaRIkWBdN/bnOcajMNt5arDzK+IMNFlyP7K
HNnkBKmJcsC6n41RYS1n9dv4ARUnINgMEvNfuMpJ/83Q6kqouqxXlRaTJxYIFPmxpFnuqRmcVRr9
zxCCwmYv9d5304oIkV08FPdEkU4gArEuMV04myJOGiiFCzgtH+MIoozFDTM9NVsOj0w16MlVvyHO
vqR7hRny44z1hZElD8jV5DtxcELceqHEpIx9n/95Mr53r65igTktKkHAwFWM/UZTtbNAsK0Za1pf
S+kR1TtZhH6DUvcAoMnOpRFAOsGufnfTBn9RYSnRtfcedm4Aykpmxl2ZsbQgB7rWXW0OXkNTpG24
00dukjoQpW2SYS66xSbMziU5rfJOzPwLsv/CVqbqPwDmxARkQ+Pm35r+ZfCKSguGGO8uKmAwhUwR
wCm6OYud1BRWkMSTJOjOqKIX9F4Gl6hKGg4reFdVdB01CK5mwAcd7cilbnW2DSlk3kcpGKlqsBSd
0/eIHKNa/B9sPTYC4tBrOKZPqdZGzSRmOcAcTowTZKfcHltmlKl1lf5Q1QOqw8lLyFvhXhKjn9n5
oQMKXytT9zuA5w7MHksL73XK5my5mPwi7G/ogTwJXHkbZ8Pn/Yh4Qb/x920yUD9iaA8jOiqa4ixw
V/PKM3ACxUJOewLSA8Py8cJtxXeEvqbaGlIJZOpTgXrnhDXthMQn4gFwhnwW1EgsHBZ7n95zAM16
UautKksicOhC0nUKRYD7uJ09L1fjGu0ubZBMQ4nMzp7oo7lp4JZGaCZtnuHgvpvOnkJjqutgzwKd
chi08bBDSJ38pvk3Ss4hIO/hsKYJfiENfgKmxsznNWkAmsTfv+jeVufjv0Er03MZqvNqmF6QLaJH
lpmvlaApnAKjNPJTGe7fYYhwpfpiPbWVPUwZSZGiu/Lb+l3g7yUjL+T23o9slWiOBnqD/z+VIKFS
mXeLgW0kyfH7Olb+43+PCUThVMLjyBxzeMJZ6FAZ+0Zqe0JayENWxNB4web+ovwNr0XY+/ACSmxJ
S9GBVXu1PRyBA5Y197Et5E9A1O40+FdEWjPKCFmJ5C7reeNtfAzlzu71Krb4P8fGJdVzipUDsoDP
LcFV3AoVIGCnQHA0w3MVkdqPC/ug8Rgm4sJTnpvWwmUimQeQEAiB4pvt+BhmJOLxCUlAPCvWhxJu
G0LbQYqt5TzwsNHDI9bgSoNf6whnxoZqTknGjh44J6XzbSZs54Wz1V/4zghEz7eGMu5qyAsA9pe6
1llfbg6ah8bRUfOW0lSRuTieylBhskEMvCvNtLnuLc/Vo2ynGQN5nYglTb3sKfwqtfoSXtSIw8R+
bkWyFxdGgVx/p4CZ5V6ESHlvDtosopRCBizzoh3Obtb9hB9MsXN/DtpPRc0ZJ2n2N9//P2Jkx9ah
DIrFnOcvXKQz+JCPgUMFvXfdjETwDBZ0XnbrWjWQkTBrQBmOgeFXyyGpsz0oH+jYryVeCZiBzPjy
PVW1KocBV2OuEy3YuoJxqULkquJ8YLWyVoDk/0xMcmojj7X9xs1YlkT9x3RZs8wCJ3ttwz5C5233
kHJXpIshJu7xAQgQhyEdzkrYlAaRz5atKbCGCxKywgcGGdngtxxlREp0CpR4mVmNo2weJHpcuvBl
yQGweh6pvko8fXX1qD48Ty7EVEJyxWhh0qmjOhe3+sQBbyTEhnFS+kgsmQdTBzOv+B/uo7D4jH/l
Ro28Sqt/xAi3c89fKyjn03ZB6D0+sTYsD39b9lTE8hcj8QHlevy9CkQ139GC/FrHSwqOhNAehfGm
xJUCPXU+LpoSby3Iad84rtup1Sys3URMG9JjDBSyj0B/KkBppo/0rhF1O10uAwEZ6OarH+Mn0H8L
x8uyQ8G+tU2aTJet18+ExDMQte5d/Z4+FfI+YBbx88MBxma14ydAl9G0gaLETjHIGdr4doDnSRoV
oNxSExs8BHJ2OIHnFCB5mSjZbY4/cImYKg+MqxNiOL5kn1JeulptNCvtfu+g8WzYlp03034zVWmz
Nie5mUeVF3JAJOGvMlTmw9JUUwfql/RIfxQ7uWblHwmjSBKz8xqh0XPP5ddI52DmyX4XnTbT4k6R
xwfZaFx2+0g9TkXH9m8ZCbvQt/ZlbuU+2j/4DpgydxwHWkHGZbfp3dDN+P/6TwavnaFG3xFtQYwn
+lo7k+ek3z2C7EDRXY3GjLDesW79tMLAfmbljdKQxnLVUP2/YxE4supNHm9B9OJn2lTnCNO7L8Iv
kg0zBUCBLLziIfOcd4/fKPQArlz89qvx8dcrRW+l+dwFTEKEfPocRakhcjJDNFcQSDwglWUG/w2u
6rLibwgIsYS8GUX6b5iii3P3YtfdE4fubE2qpsU0rItFNsJzEhI6B6yZZTF7L+roSvhhH5gljVJQ
i3X+CDoZ/9VDlm/jgHXjkTDtk/Rkx0P53wE0Cawme8AFpKfmzDrUkX8zNjnfBS9eMmCWwOW8kt1G
FL+P7Yn0KdzKprMYE4dzHlRnszqWBk3yGsSkHA9ndvJABt+89CkE2flvi7hAU0DtJIJnPfSHp8LR
MjSLYBoETEp5iC/B1IVa2kbgl5QSl+6H0psX1PGRr/f3ouYe1ViLsI/MuQ96+Uq1p/RswN1dWdvI
ZPgleOXZYfnNBiJ+a3w1cNPoDl+pc91/elqDZaBqPc9ESkOKgtKaL9q0Yyh15/G9WN4trDYcVZ/r
bLqgbOJtzCYVSF6cHCW4aCECnwgpZ2zSrHB/yf+mHyEeucwc2cQHTaeqWBs4T1b5ORzwUhvBLb2t
2wG4sHaWV69tJFn92uMw9UPm/73GuYkkaHQSkWUA8nD1ZzveNixoquUqZEBGujOiiLh3HZVe8qKi
y+zvm8uh8kGGTltweugfogtOT+Z8rPRTz0OdcV2zcv/8FwEWsZusdiF6b2zm4S486fhZt1v6z6oa
lWA6o0jRWOoHOpOut/JhldQ7Yn70DeWNocbaEckWBDqC/zPC7HqWKb9avw6ujHZnhZnMJ60QZCfB
T9OOrvuV4lQ2CsR6/pNywWGBQciDGxIc5Yx45ZtBEE4FoE79GyjKrkjjHwK55NQupQsEPBqyeMQn
pDo4ppf72LoK9GTRGtSKtrLLCkiUOlnKXFwVeYD6QJbQby30PIevXxAsgsmIn4fP7+hAIFGq7Emx
nDInDKJb2nFdgSLt1lRbEenDaD1hkBol/eCA7ifvvLytRLOakIGbZnlKxARD2VSrfaymOlPJfAJS
YVOmFNrhyykyiJ0KpsfiO6nePTeQEUtSAt0T4etdwwx4LP0Ye6GY9CTUT5ddUMqcUrV2iDA831NO
Z5xTMvpuKZbIjjOU1n/aIdlWCYvJtXJoySCAnIfgBtARksHstuWUKeJwb3zEpNtgFt+SksXEGoKV
2Ph7OA22PlEiC7xDT5pJXoWaRYfnJ2w083nE6Kzl+bd/zflwMNrHL6KUREJ07sIYhDRpG1C3sCH/
v8rqeax9sLMVORCMKbFARFbEu5JBHyxfez7f5Eh7nsnKmwQpWWL4VFQvdCozdKLL+WyWf05XFetu
yVFbplYZdoDbSvlpVfC/IwL9XPALqoumEIFBlfQ+jGyj0I+/ih5APqodGIPe7umnoOGQ63KpicDX
imbZ5mC+sr/02W9JtJc1uB0ZnL7rlyu3lGKIv55BgFaAwHRoRwvpBReBmHY0EPiFfdrdN2kg5+7A
+qXfkp4LdCNeDBZUgiE6mAWdA0Vj4fWOl3omGuz27HgHyFFQi+snUEKpLCNNLBawpBzs9gLgdTH7
lQhHpg8Ysnzxsou68tGjFUEkk8KxE1U+Vli7xg2IoWowk6NOEWQxKMfBhTpngR8wRxSsPlz5L23O
+pCuclAhcx7rNrOo56LczJihei7clp62qaCIBpKcFd8qw+/nlumJwCDETScVvpxQiPQdqYQ1kaAM
GPesRiTYZRtINAV5MIynh2l9+CLhT7qNyUHsnZXIQi9tJ6YzLnlRGn1BmB9QKPOOsidRi/Tphil+
uZLThD3V48VtgI1uZtxqBJix0fsT3GiT//lj0X4Tiwls1+IvXqkE3O8ztC9JSnknwtFm297z4Ynx
KT6arbhBYM5X9+bElMqb0ln2UR48bG7vmprGrzBr2NiIE+jylwP7hDlAqiynSX1u4OwVbXCBg5aa
ghub/Po6uQWOQpIA2YfcCVQRuzQFfsACAlb37rb3wS39ZiLdvUXnsku4rkwFCBoSWNf1UW2qn7vM
tSRmfLj++CLvWLqZw1iRlXwv8owwSt7rIxb9SvT2QglCJhPVVfACohHt3jfccIVt84+CvYXU8M9q
vfHUF/5TunPbJNYN2E/sEXQgSEYTFz0LkhoGf6bRboXjeCPcjHqLUPIeiuM9k3wc2Hvr6hRQW4Yw
ueDtyAonyc16i3whovZCwzHk0LWMPxhcU6nV3CNDc6b0H5W3yrHiPZMHxhsxzRuD3ha7ZHnZMprO
qkYTN939hpUwbrbXH83uXuLb7Nd/X8TvI6OhLhg2fVwv18KEQuOEC3Qk3fODR3vfb8+bYdECge2f
MM3wbfL52rukm3Roi78oqhgTRlU9z30wivUHkhfOyz77yDG+GDpDUo+vTFJV5xECZz+K5p8ciqw0
kKXmohAPiSmIE93pOcKeYeEAg5BFMekkd/Qd11S68E1RzAxY8xYsfBbQVmBX8+zaD29rwrONhnYF
IS+rZXzFKH43F7zsszr8iQyDprPHhz+EpJAEcAefnduhwrR+TjjChxc1A/uJSMEmOXyWkWh96TOP
vY3/PVPxZ38Quvy1gJzUCvOVNlJaoABqb5Pv7anZg1ud1d4MXQgLgWojuhTPqxTh9FIx4xsUiQH5
s5e8NxsiXD++EHDAK2cLkuHk9B6PlEoDtO1ZhTKNAThIChCYi3ds0gJlYtz2mRnppegq7WiGEoVs
gvOtSfcgq2Hi0UWqEddusOu7/rxe//IPUqsSVlU1yPlST61OODY54GxR938usC7k52A/TPk7jxDm
O+c+4/6ygOszBBzSkAIRvaNsILWz+Dj5FVRJiRuL4qXHCpeY0IxAxHoD/8kgqUouJ9QodyptZI/D
5KgX5VqJnmThMtuXH8TAYJCK3ymq9JCmTF9mC+daUF1XSbzQkjOSXhghi4jItloqT9ZCBwH8RdzN
1LhBK0MVPGL9IC9PkJ1X4CREQea7CeVW7KIcm+YdoZ3UsVyFECZnkDd7cy6q11dsDFlAp2dh0ibN
MYq/H2p+88LcK2njhQklVDMOneSextfiWjlEEC6hVbpB+bNZB0w/bdtQhNeO+i18urexf+PtaqIJ
wJQZj4Zex3Vki5z/CfjGnMNugJtKdxMKstgU6By7sYz6Y4jjvbpddcPHL/SldQ5tblk4EOy1k2lR
50KFFSR4m8MTleJ/TLtJ9OP3QNDbFd7EUeh7D2hSsU5oYmq2q5ZFFU13eFSEhDKXmTocKh0QPtrX
LUPrmAyeVQ/AQ7+UVXlln+7Si6+uPamj6Z1KsICKR58bDRx9tmwHlhawM65nQ/IeVqvNWnbcNmoL
oJ/7pwzE+77Noz2vWDRZil1WBCLwvNsKzchxFHANTF7Xon2LMAREaK/jX3lx4Ifc59dNuaDxS70D
BiSDwyiy1dTEk4tQ2ZcTJwFoSuX26m4HfArTat9XLuVUERO8eBaZDU6ESor0BLtcqZ6+BZGsHLC8
eYGjD77pTGcQpMdGESvmlo0ZYFa9ueznRVPeGt+uMzx/4ghW11gx7voqOe2ZBuFYS7cVBlHMnK10
GW/zDXdv6MWCPUOfu+9Eiwv6n/Fqsl66u+YH0P4xU/VbGOz5efEHzpx5dNwfgpHdiurtgHL53LbP
Bmianq/AzizSDg7gqwiqVngl0zoTInRyDMLPQR7aixOLr/LZxUeHSM2oPGcRZOn/oiBCnMK43uf2
2q4gDJlPPzmDgVGbm81+ZJbizH7Xo10zLQJTP+mPcPVsQB20GrIlm1IcicQaXSV3THtd598FPx8e
LUrXt7nHDZ+ELvq6e1UEBy9SD/JaLno6O67CSJ5V8ghgxx2r/U+v0+nsWb6OMJxsSqOzN1wJfu6v
NijPqAVrdkt2UscnBHw2uX2oI9XrEWKyqYXMZuH/RqJETegzYROTkX6dbefP9fugIlppUKdpKY/+
VeUTVeKs8ZYriVB5GiHniEh1tWZRpWhpzKjIMBxbKdpowXJKX654QgkthCpRTAKjB4LYRmLAI2dk
tD9uh7qV9dWk0rJzoxJcg8Gj+12M4Wrkfi3uj7h+cdzovcjyl3kSwxXhMkLcEK1JvWjXgT3nMQjJ
o+IWimGZ4RcX2Wb5HGzXxRt4UmJHcZqUlc30qTbkU7QZ7uLSv4dc95a68VQPXccJrpXU2Xg+KN37
eQdXmrfftxR4E7VyRKDn2HSeVolxiYVpUvo/N2+mzaf1P/8MlydqXxKqoqZNBKfflUVHUxLVig7x
K59vbOFroux0oIB4GXcEpMQHB0C+9S8rVwyFCBJmuXF6vyCm04euScrA/eD2Gh3OUhyKd+AHF6nO
ubsV6UR6Vti3b7oIpg17kVRRrfPO/B9MxDwgFeLn/TrO0xxI5E5nBJWK3z+CPtDG2ofF1L45Qg94
RjND3/ChEB9pEgt0yeBIpYb9RYiWaM8Yc4XZD/r78ID7iw0i4vOnzSCAVFShNoSIAeWfeZ/IcO7Q
YANMInkBo1bE7SpWdK9Iji24hJv1s87Hhtvm79DO+W5hhskyUmMuZSD5EGWQ5mfsSLfzzuQ3/R85
AJLZzBj9pHs2beTuXtdZvL5l7Nk1+4xSkhGDYHu02fTLAkuF0Mq6LEbMDyYmyVEcXaHdXxyWh4Zs
ilqmqhm0PAk0S0MWmiydFZ+sSLNmh6DLQOZ0ELxjYGHMsMRsIN5T0q+zZh6wUxujNZolJA1NKUup
Z0fhpNJEElGHxAfIYHYklDsgOPKdJNH6/twIKcs8VCIyaKZCLT+edHLdMZ8LSm0s08V+HjN2WRjh
dedy2r+d+4GhL+KI19mz3Etv8BUAuSsbiKIHnBu33I1hsr8of+9+8DD1vmNK7Yu0Nhb+aLY6sTTD
ew8glXPyv4ST6H3dufd/8bjolToCefDSkgX82AHZ9hdf714GNNtCfhqd4xZVflx4L3u4zwOwN9FQ
Li90CmKt6k8lTyMMkJL7gUAdbO/z2kGaDS35g4BM5PGaW13jX/hzHH2C9aG+1Gh5ymsA7k6b0cZz
a5MF9KRerbbtCd9sxKNtOoWHOyLDu4CwKM/tzvKbfeTaAoIRZ5ANHokopt3X8d24Gwew0RorFXJL
QdyD6iVSGYNkvBEKvlRabxKGndZNDfDL9SEdJss2SML8IJIuN6jjwTip+VRxPFYR4wG+pSrYPruH
D3HwzN9ZBpjH/wNohNgEc5Q5l4E0JnGY8iPUPVzfKRZtFJr5cFtVt+fbRr0gZLXtDPrcEzGLraJM
oWQ0+S6T+YGjK2qQcHD6cRlkD6LxEwO2iPsMhHnTKzUAWpFNB1eKOmVDjxmPxIGIfmlfslsRPp+a
0DOgNz2q/G9eo6BwUVxVSE+Eaq+zVAnWIcswJJRBaPeQGsEj6MwQ8D+sn4oPQUGfLpfqo59EdtaO
1A7TepFrE2rco/F51ZYdmtiEwrSJNLyR2HxL/YPY4yMmKr2WTI9sZLR+7mtPM6Ues0gyhD5l+USW
GZ+lU36pNextL9VyfMmbWgVpJaBTC2l54G2YqKbTC4b7NM49GPV9Xv8GvuIhSZ5gbynYBoE8IaWU
kJB9GbwzEpCp0rJbCFCsfYJEgZ8+4pk11l+BdYvgoBVbsu0A9gZiINDn/aKkyZ/lUZ+eTuJO3dtT
IGnGMx6Ozot+YnToKT89xlUi6SHZztvtoa45wdTWdDgKRE0+TCF6y3K8lMqjC4vSZNHV1wT8Nbw4
6tZMvMBvL1m84ckNRiTWxmj28nGXESkUSupnvLbAjOvDxVq7VqLyL40sEC6BDm+f6ArHJjv8xoj8
ia1jQwicztZMnCD/Tsn0b1UX4Z57h7FKfa8gDpx62owCzsfK+1gSUe5RTHL7ZNxaNqRum0QgXiu1
ZHzkJBJMcUTDetxgFG5AUxOBIOe87CAzdBr9YM6HrVGSDfcgAGTKsR3XZCLc/KzI8+yEzoY4/EQa
Lj+MmT7BDdSY7i0s+/3Qxz2IVduNbSMR9Ul75R4i8Mqtk+T+X4nZ6GcThUbdvJ/ee+NfrStf/l1z
8oeApq+Ocyjwy72j7y5trFehNYcUo7L2qI/FnKz+MtbAfdVA/U/erXJLT7qzcApCo7zJokF/4qQK
E/BCIleq7KA/dEc36pYXmSxXFUJmSyx0sEVTillljGvTrn5Evd30b2r4zou3qI3G0zC4Z1N+ftxK
Q8TB/AhjYXg483XAjaovMr89ttZH2jUSL/W+V7zzVYKZ9jpjwSeBKzEZgtQV8B64hiY+D+0rk8Oy
zHfBYGTk2VN0Eoqr8iPOPNMMLidTH5K2c+8R0r3abTbJi9okfJh8MUTRm/H3Ckk/Uxvb6/AuqXA8
nyS/Ys79r+3qHgbyxRbGdSBnHNupQGVYIvycbg72EuCGYU14PQAUVzhTuhIhyL/gDW4j04zFyH6e
ZQ+6qBTj55M3NgCnf+gJEsUrOp3vvGESOBeN+mekGdt5fj9De29b9csywFN5BPNRN5XLiFqsZOW1
3FsvQoFIxhfaukzWORG4dajkDQrGtR6caP6VwesrdxWlfnUce6DpGG8mPNE1OvG0rKpvnBtJiFzj
bq57pW/OOTUcvLERA7DEji6Rk2Do0XjINM55eP+4LNEHSEufGujGjbhpVxiyrurZOI9mFM6n88Ek
A5U1Dxy44MNXOLo8nUTxJq8UaxOQBCZ2UpqCn8aD/ckdIOhNahX/lNRseSc+aOJuUZhgL8CXlhbZ
k516gmUYLaCjbzcWFRU7uWEOSSoVxRduP7ygP4Q/VH28lI0IykwAIMbzlnQJxxfs0Qwe2v8Dwjga
DWxdy8UE2NWfeqNXc6uqx4bIM1VpP4H6saOVWdPJQury2SJY4Wac3eGmAFDGSOth3DFKJ56UA9+d
te7ZbvpX5xOTqNjzSQMTs/KbPKdrfQiaj3CO46SzYYnN/nCSI/jMZxym31sJN9I2lDwRyQ/rByyg
QC/h5Cp69ytHQVfBeGSO8D2AOSBvPlO1GnpICNTLd8qTC3byuN+zxTEhUfJE42bH3G46+2gIdbzF
B2qsJL4J4alPuRBTtXCXtH+WvAyyhqnGKJRCaitW3v+KrG/kvkslnRxfq77g/nr7+kqzzv01CGfd
Zgo/6kG2CSW2D9/kGaR6W10yd5JdXfwBiI91P5us7np/+Z4IskPJz7TSpMyQ+pnJ/cLqn+7+5CW3
4mjauIjJM8dtcZ/es2+rf3nL/YRUcJ1NfAKUnzt8+Pi5c7HJdtpgxxc9QvZ+raTnY6eA+zGe5GNx
iYi/8Jnp6mEe1OblOlnguQ+QlwDMAzeNkPiUrjmJoDehljWZGzujf2m2kGKz6Jp2V6b9g4fYjNk/
K0Bq8KRCXKxuXk2R0NTTkoCoahYmGBql4o/kYX9njO8IxkdE9/ICcJ8Pde113aax4/nSzEWLWl0y
uAi5SgK0zwY5A00mAsX34wQMVpbP6pk3JRq/2BavYgi0dkEMz5Q4qzXF5xcGQ4ObZIetu3Bee+LX
DLL9EdAGPFfrjCxaj9AlvVCO16udMkpeAqrJYkOveCiYqZxgZctPX2HVxzFbEMExKnXFblT0X17C
ZsSf7Xu88yzUlg+NkZaXs5WVPRhtzPaTZ62ZUGRS2VRXo5f2B+UMWOp7xFHRRpY+6rADvDG8dSTu
x4zxscBnw8TTnPO7qfOh5An4Iwve9k80+8XRMN2MVVriLdZ8CLOwArqDW2m1xWzEKi1LvH83Nn+2
HsT4Mgqf3E+nqq35VgnO2BzAkh9vagBrzfHLuCA8z/q9n17yBHyc+xdNsMk8By12CCua0xGkQU+i
W93sgAZfRJrA/pcmMnlp9wGk6RDCs37FHu9+F0pED1Hj3EYxNI5qaQkDUQLQmfUdqktDFaa2btd7
Ilk0eIfLHLkWMzchM5zpKl+GBcIauRMa3zOPv3GJq27hlTlWeChGPL7qBhkdFI9k5BQnFCMl3wwD
eGb7YG8c/kFpt7GpSJm71W3YtHDpRAtmxi/RBaArPV1nwU0OurJLYdbDbg5ocZMNIuO9VwGjh1C2
rXbT041w7bVfmI4Oo1wW3pwSJnZr43e043tb+jMJPWEIpFpFgbJfnbnagTQqH499BfFoYF4o4fJq
APruTzHkT+SxqCsZgAGlg46KRpVgyg7QtqMCD8Rq2FE0gtlNN7Kw9qezPSfui32MzRtMMPIcOfMh
2+RbM5evniIwo0tYKjA6PaJpnQ9UC/opCtOktua8RYnpi2yyPclYnalP4CavyvGYOIAieuxn86GY
DOJNu1OMaJxUjjlqiaKNOJ5BjQkjZZt2ET+SjJdsqtXIGhd5GpUW+0jK0ESu1ffNsFl+fy0x2cta
ygcJLEzLeP0mFbhpZKNhaY9g3FIHVtJiIKxz/20mdnXqEIWLj1sMZxNcLlm4yy7Od3WUZFtVD1EA
2mXwahaQK400RwOC4Q7+HHOyaTuAAGLX2OT6H5ONTCuJsz+bCWXnnpzTgelEylC6NN6IAfwGXP9D
UV2MXdcAx+jl/AYjzp51/fqrntPM54e3sILqYqGZ9QObDqHcL0FSWkIYg3OHG72iykqdZIQQBHRI
1L6VnPNoERLbx0TFlmxwLxA+YAqdk4ixWZlJ13Moz4dDhadsNtaG3sw7/7nGEeUCkkjvi2/wQWjh
izw2MWYD3vrW96K76aJV/UkcwXYamR1OxQ/z05FxtmDZFJCW3YcIBMhEefNASoJEUw2jwF5HhI05
VylpIbVbh34ljPJGfFSJGqOuieagNbFmuXFWoRDmFa41sKSzsYFYSOREkciZvV1VSTHoCORIQlsr
eDnARNh6ePOScqwO+XS+IB9gDMjX64zzrkmfNuPITc5DtunZmIgKc9fusulc0XbAEWjV7x0/SRzx
l99UXagjlO9S5HobjvyO3ZaCLh/+tE5BZQXOLM0LVvELMHNYCzQIjSclzw5JvsPre4SThfAM4jE1
I0vzqqUEsoF6wHSNe/okGpY/JO/yB1Mqqvwqdw2dyMMHvSIQIhIgjyHUWLZNcsS+u4rB4dnP77/u
96pEhIlrQDddr+7N7nf//xQvMXfEdDyF7v3wENy8mZy8eRUc+eX19Rs/VXPil8HtIWH9HffIe0r2
RonyZ7l+t2ZLQt0Phk4rGL0OGDDORAd9ieWZp4ZLSgC8/sVv/p/B/BuXSHtWXMEuH6wPhSqOjueN
pxyvLwccZ7QfDtJCExUMKlYK0OKzwY+w67IMI3mfKjQ2zdqQJlkgKH7lQL6vnoSB1xWRMeXEintt
TTYr6v6wG9vEagf2I5N2y+pB4HpGLdySaIi+hnDD5dk+PlyBON+nLppmnxDNiR2HFaPE4BCB+llA
v+NVZWM1DH/sbzKG38J6A20DK2Kj6ku2qO3ZTOHCzxyvu9Ui0GeStxMKLdJrSgaJgbgJS3ItA9tT
IOK+IBj3Te5hySJJU5T2ocCUrIKzSaHGNJ2yKn9OE4rnQFGpC1EhkeIRcy1L0oJayQZXQ5LHDaG3
5vxXyc0jF6sTBfrzO9VnbR1GDdWfEks59EVNWO1aqwRUjuhLqlKAp26rKIe/6+9F9lgqkJ5CSwCD
8kFAc2AWICdTnaFWQybFpApdXBf1ZXOQprAYP2pvplP/fare1gZTdzP0xZjcLGwjqK+X93DdvrMY
SAzB9IthvEQOdey97xgJIptz7OEkGEn+ghx2NuSnC7h54ePKTtMk1yt+CDYBTW7BUSNPKXMYFKvA
nreeWbb/dPkilPjXkKaB3A65P/72WtJ3KXq1nEYNIr/YtHFSkpdB7FVDCjNk8YcX5p+xBKXH5RvH
t15aTrXpAsahmq1ZZXMwydW89LpF83w2PFAJoYshBNAt2j/M9xqYqGulOgXd5jinWJVaVDcJRWtk
Gg/Rg9NQ7GqI06eJR8QPlzkj3p0k9FgIWIqOPlIY3JK7vf72MhO14ptwaciX4BFeEMWes/VOVlWB
Er0KfKE+HdBXShqT16MNG47yUe+lasg5/HQyPccC2fa4v3ale07n3m0qM2IZ8sALZAxahpkJJheU
jjYANHEVK3f4xGb6hnYZd/KWA7Ji3mnosImwevJCi1ZmRS3IfdiCRX5U966nsU9U6vZeyjTwNCac
2k0mwojtGCcnRxrvCfmTN2FRLngbuwdHLBslMgV6RZgHjxOpiHQDWNSPLShPVFU7+UlQHn8GCLzH
dqKMGytwzuA2w8GQUC52Z2fjADcHXmqQkTNV7L5DX/y1fFskQM1hcYU2ezL3mMlQUK/7Db/xJxRu
xxm6Rw9pPV1u7AHo4Do70VwJt6PaR8UxODPTMME6m16TBxMuohazwm1iZgL5u0Yb5/Hqwykp2J4I
gfA+GIY2GEblGqaMg3ciyLHAWBVa8WHA/01CVri94OGkqQoyCuNuounfQkSOdLgW0j3zRT5rAVQ4
uYFHC/HEvnlbym/shvLtZovsb1jREHXbFM7Oftu8lGtyygNmv/IchXlUWw4Iz4fgS4cDyvt8EEmW
OXqcwmq2nWMixaqIOhTq8cTWoMxUMSw8nT1db9SSdq6vuB9Kx81E+QxavkOZMsJ/LPQiyYR9Gcry
sVBpMLLypljhkVxzxvRoOlcyz13536MV4H02kl7LKjsuzH49MkzH+s9Sqox5Lq9Od9PLUUvy0PmQ
s9LbNFliBv3r43QdbrDXGG/7cU5KevEXkV5illJn/LdAaG60Ufy0LYa126zcpXbE+75DTiWP1XHc
kSRDFg7S18Vp6xPVyArfoanw2WFnAAoyu2J9wfnIYcC88bEJfpC8SvRO5tZ/ZlZxOjAslCkAKI0n
JG6X8GuKnxMVEWwSSjEOeFMeg80/cbBgZvXg4n2Wz7A5NpY0kFVntRefW4GUNxRy6HQPpikh/MyJ
in1CNMWWhtbgEbLtiNtk59d7v3KoxrMAFtLt9Qyn6wGtoLyxOvsPyGt6f3sQGlneGu5MNeS+0CzO
IU9I3aHoX5F+HfM/LG84UClMT5KIYgulO20sXmdtJ6hoUG01XWaEPDkPYj3LiQNKH+UPCZ/fTcDv
7KpJdWEiffq1GRl93uScnwTjjyHlVv09a8vAEVc9fNPHsGogu42O8UNTx7WkvW7zJ7xf9YdAngjz
BFdshewYAVEGzDHon0LUXm1yk04rsNk9owQOoUQhbe/Oqn8DzZialF+RIOo3RsugwmCmorM1jK2v
U+8+hNQA4jgaP2cOus9lEyeoWVJnAtcvXfDAuxTwswla1h0d2I+/J0HqMRPRzUW6yZtLI5kg7uC+
JHhXZQKETuu0QuccBgj0RboUCbkdo6vAb4qshFEIY/dnj4c5fSJP18ThJGYbA5wETTvbJntARltX
MBZ+3P/zYHbxk608QVb1K+gm8c86TIOBIkxiiDbCuESWLDrDlkBat4BZuKnepoDB3tJEfU21vM73
CzeS9pNELKT80YwNM+TqLB/4Vh7+3OdSYvcTOE2XQYAitPuFsOSAY24ZBNnKPlppefPNnVjBe0yY
1t/fOuyYk6ewaTW3KS4BXtE2KY6I4u22Bvj2jenvOw3lXxtu1WqI1Qqbc4SMwNYxY2mGDo7gMR5A
Ppvd/9ldbehmaajxCSiBg1ccdN7KT1KINm007Y3hEOvDncy9MtyJa6SS6U8L8Cs1qDPHSZ7+v3CY
nTP2hsrtBE7vtAoGn4IdzJYrK8V5lkVSibnuLbJxgdGAeE/wWm2Va2OQYw2qKcqtMrIwl0SM2P5S
LhD0KfancNtDtzwHA+3xcjvY+6I+hLF8QrOJO/OsH9UC3WsGtHMH3FLxdqs9tl3XeQ6OHUCbefeS
ytWo8/kU0TBoMKqjtQ5w2VizWwE9e0jFlZDAnqTUQccrl3c2W9BBifDIQEcq1Nlw9E1Fg286Obdq
TRVbzhvlAV/mHZirHqczWERF1s9r+T54EJEEXjlbiyke5wNmOA5k+p/Y071wfXSuigFSk5pC1MPD
tbl8aHVe227UWiv3kpp+RKmX4OGUTbvyPTSl4XHkwlazb5WdprWMsI8si6zHXcWo/qd9NJHgAn7J
8Vrh2MqrQxUsHdWShbVdIXWuoY0bagf0EHhWeAy//fzrJaDuDMrjrx4WHCbwwRSguklaChvVpPMT
1SpS22FT4Yjjaw33kvCpfoNa5hPz8cLp7QP62GNAm3Nelta+ahgvlEolkyMy58DpiqAhBxVZ82xP
Ngomwnio6zN+O29alib6Mi26TQHzek/q8BwMhlZCwO47FWILTcPoGeh3sCX3BRGvPrWJme8AGZsz
nH/oJ4ef3e+rbw7oGIX1pICnx0alACp/3GxbLSl12L1MIlZc40Wi9ua2k8iDyh9EFcwvNF6kvTiZ
2qdtJU1tiG4JLu/iR1B8ybo1gvY6xNSoC94gBQ8ghK9bo/MTOZTe2qLvuZuekO2424Di8Gmb28WB
NBc1O3sk4WetLFrm2E+zx7VIUKQPpF+XxvNFkReGxUDj1MPYV2j5Ngwud2n9XIr5/kG8802k3GTS
uOx77AKK7dPMnYeYgf5yrgFl3LZzMDMSof20OWL6YAo0boy/vdM6pk7OFSwWdP1tpDkY7Yp0ZXSj
lyRhpCeX1TY5B7xnkyxtNs8sHHMQXDshm8vKaiRVywxFILeAV2yc8JmXcc6ClA5LSBp0izTiLJS9
UgzM4Gwa4xpvu9IUXOdAfOd05R9LftoRlhPAK9/iOEZZI4kBT5OJESZOHssu4xysi459YFYzPZ6Y
3YlMsax9vJS0nmbc4gFrbrOU/CSUKr7hws+8R0d/8wCIET4EQM1wTUSElfx4e44f7PpUye3o9fLi
hGzsKYDnhVHx89pSFkMuFkIg4WAV1oNyVL8IamaKDzroyWQjKqk0u6yTNrT0A+hfUc/yfngEq1UU
10wkA8ZEBcVxVu1dooYwz7S+00AZZM8zsI/ws3KvZaaIrHzBY8q/Ycip4yPBThWhbJmQ3gZFON6g
WcYb7luEPWFK00paR3YMgPlywPRA6opUkGq0VxD70DoDzgy5SmxWmmh0gN8e0zcb7Byy+b/0CpwV
CVXEMW2GlmkjQ3s4XSX+oZjWI0O/4eKlQz9S5dNezwnTxahSa2oDjfsSBD5IkpqXkccD5VAByoWI
s19LISaoHt4ELPfA75/CRGgvqLqi+6mGRbPhU9FbgI3lYfTQPnYCIYT/MiD2MZ9u0xDGeqfMjQB4
dYnuxILkYy3zgw+SGsvmI8W6dtmyrBebUuiK3Km3hdJde5JU3A0n9WhVmm4eWY5WfbHMEuSaC0kT
6ZTdfmUyeSi9x/PaB1oxOBNUfYxmo37mXsHUK76ekY5yVAPdEgFVGIz4KFnyjNAqaQNZDaLC3ZeM
1zc5qAvp0XQk6DglVWjpPxwmUmxXHLM5h+b2n3qMY6zwWZqbHxWQ94u1894RYnTBCZJqf7C19IAm
sDp8Ba3rbr1A19nN0GPH1+qvBpXSg1h6nlfTJIn0WkFLGzlkKsiPJ+rSMCsH17T9Xcxz6VozHVpK
0skdDaFBdgLB2ifvb2iPGeBXnbb15JClmeUMdJIduwjFjv62i5jKwfVlABu0wUwB7VdPqeh/am5w
UXTJfNO5xWNYrXCsdIBM+IpCp9guaP/+Qmsp3AS+8+gBkago1FJjtCoXCz9TAApN9wiQtJYHqIgy
uVIiOyfulhET+mvdPTd79IJz2JwLA0tnX07ILKr9918jZ7xzs8Kq1UqFgy1KHf9ARcZHmD67XXYo
GRFZD7jpcbjjodfMzm1ZDzdQZvhg1a+jTMDRCGNwdB3VRpoK1Mco8U4r/Z2eBhoCn0ZCG3KwjDL8
I/99yBqWk/82heP74cQ4hDzcBcOIBBLq0jWp0PoUh4ERzLH0wGzlymlI2G4GR9aOqGHj33spzi0M
afaOIpy4yEf5nxrL126wwUPyxqKybeoHFTXwFarNIz1jHwSWcr4bYpEo3GDCpWYzO7RUG531xFWP
xZ1qqUlmRj+uthGaK5EmBi7Mxxr91/nrQElnE8Zvz54mu9O/Qvwe8o9gvR3E67HxaZBx+EY1/PGZ
IZtalhSdlMjv5bzB2tL++bBdx8T0NdF2ivyF9si8vxrNuzNl3LSWf5MzhopFdG9vWhdQ9ouYWEdZ
76xDxyABYo584zsQ8bH7U/zLxaqJGKEGigXeJc3fC0GIc3BCwlRp1x6UjRn9S23DLiK6TPulU6od
CfEe5SyW5SXeiOGK1dcXEMg466EIMQUN2peYAsfXfprV/HnKEIy354MxEurW9BxGDKYX/MY74DdI
/wz4vsDWw1RfQ7lvGaN9TSkHcy89nN5nAA+8VxoKzhRWAXChPUWaa1qNjaiLsQd+fcV/XbSX9K9V
vFTgqxUkrl7+hqsF9G1sSt1dbEOLCIdn/ixQpQG2HtJ1PFRg7KmBnapyiOConpfo4mX6UQlyBHxW
uAPfStda7jXo2jOWtZJc05k6cAg0LYWV7xv6UeyFXFfuddN/gBmrVumY4jE2UAyfL1Nb9kwMzyHs
L1inR0Hy3yJ2iKuR5wTmsDXX07x6dENiqznsjQGlampaCIavforXLcYXJ4BUWBNJGNfM0mTSIsSQ
4dHjsXPKzBTEibPJabYTCWds86feQNCSqe/vUuxYHddaW5Zx7vkLvAjl6+DcUeNWFCNB2wFPvUGd
mvwC9yNnoxowchmgPbzQ8N1hoaASfq+UAeryP/eRGbAjv3De6UymmnJooOVJjdz7eP41BHzaIaai
ZzZH4LTgRnnR40eUrXih8tRswlc8KmIV1pZBmpI7ISp3kkXCsxRUj1KcPom2ubUJciI5eI2ZZVNO
qBAQ/rXKKYcz9LxPsBDPBKHXA42zQPWFR7MToaczTD579pccqUDOnGD62BiNenKqswxRGbSSNb0Y
NEA9VgeO1ncEoz/aPyq3fpzQ+YTmAOSov0qqvAuJwJn+ROofr2YJ9uF6dMM72YRV2BxUe9S0TQz5
+0sAlV/vz5XQk+3fn/0yLOzG8++Si5nayyCNBYZY1dciGeUKd6Gq8nJsyxa3KFacN/GEQfwjnvi8
CZ0jiVzXLQB83bhJEFYstwIo5sNyRK8wIb/r1MDBxSmtV33Rg0BLDsWy/AaxCueGujVfnrtBhPEI
A/3fH3qys9zN+GVmWEkaJF3ux1aJNa25/c6qYa2tv8gCZTq9g6DLeBXB7KUjDoLqL+ZOQTXXxf0X
gmPBO5uQoSvFhJtSjMWwkxJk32Fi+grrppNQofLYL7+yvkN4S/lZ5LySAo2s3ht+PF+BhprhbyVC
zqEAwn+VQCStpKWOBH4B4ADydUTSfBaJUCNTWRXd/Lcll3SeJIfucUpXG3wn4dTqR46DI/CCUMRq
bebczFN1TjamJTdoI3MVCRr41ILbsMUfst17/ZAvSifcAS3RN6uAexVmHA7igegXYz/ZpOPoU5s5
97RxzNN3v0HMJWKMOkXSq4qvS+Yptxfa01gP0n3xrrnkbA7lBQpEBi5rXqRlHpWbOV8i8dc4KTQV
vWZwAMhDibhblGBohKgTuGOX2uh3y7+kbQwjLwABPK+Mw2GlLVYtBsvJqFPWaU/J3XSbQMVhQUSK
e6BdchFOFU/mv7Mq3kbraLGuX2xtWkqr5eEIN46UQYPI5X5I0eNrPRXn0Ae2D/3bRkb4kXTWS5Y7
LMTTO4E0qyWO9juN27Y5t64XJrEGLArn6UVvdtQTn5XP0cZyzK7prMkftlU9cvSE9ZpLlChRTpyN
hBKvgNRzdJri6fM3h8G7ka04KMfuw+3loIr/uAB9AunVayJM6K0x30OpXpVk6QA2vp/BSpiuSirP
djaB3pv2WINegHArqGYQ9vFSuqvqx94r07aApdsDZ58xMV3C1j4Q+nFghw19Ac3NGv0DOSFasx4E
5T5KliCvL+66BWe7I6eXrFeBW3zInZqDy4Ge0oS8DXIbgv4yDahvYtCZtVFwlTR57YuPiGrBme0D
u81q0nBMx8mDFwINlL7UDNtlshKl1lHNg6t8j/s40zJSozruGTmcIMShwvUpDz0aYeX/EzSueXCZ
nCEUSvD1osjNT1gFVKTP5RJq0e2qjPUvDuvcACWS4T/VyjgWdYPggC7NepqEgyrLNRQJ+y39sqyw
ABNLe4fo/m8ZF5CBqIAjIeXxCgON9w+YCDuXAJd/6t22IIigEV3k19XPjImkRRQMktgBfRUE7XdK
0cncOiIq0v1p4LfDj39FRXLFAq0gFHN/j5XEvHX/HFl1Of2CAzDhmmLVYSttrAF8l+EEZHCcK0pQ
oNpfhbkh+ynRlozvAWoSR0FxYMtT59cSA5B4VjkfQ03ZOYRhJrgO+tCVhaubnxwZ5uf8q0boAS9J
0UIW7xsx1Ahwm6uk/WeqOL/OhtTos4jGqudBAQFvFplvQMKhKet4dPbRyAyru2JHi1qHzpKhdPCS
LT23i698lPMbDHska/QQ3g78j0Jfdfimnl3QIKLnwKYi2fdGDvUoMavIh8U685ah7LlN4FiYGAmO
t60BT5++lL0CVCYGM57mPYNuM7PWvuaTcc+sE64cBTBOdPaIwwyefCvT1KlHxz3R0qMPekcO5WX8
8H1g1QwWoE3nSf+GbDQL8jCxHGg1G6UEz7n4lCZvSeiLM6VPkJV0171L5ZD2jRCh2nRdrkBon92k
A7Nm7cOGAgsHVFTdGB9Dv7yAWhiFzlcfpKwQTOTSsaxnrrJRRdDCtsbHrIPgwalgQrz0KWbnN0zI
vcZoLjkmPWIG5Oau1K0jqh9wd6yiXCO/uvPgEmFvdOHmGiLJdHB+VynlH7IXj2inIiS5XlcehSMf
qG4FDkR7MI8TONdKZlT11umn1F4eaoO4raUvnR/9IUGPlJ+SGFw1akMPHDpF2tRimd6RhyJnpHXX
4sSTqKz0L6INN5+mOdZPeIf0x9A9zEK6/MqbNdicQ6OCy93qkEO13bBGS8Hx1zuVIfmjD37ctb7W
oj4iDOuxiqvpWeTyavjzRBmDIHCjmSzIpO7j28z/csolS42OrTLUU6ZB0oDSb/10hrrapDyXsU0i
9EyNcKbEDIG3Et/b3S5+oywaeCaAqVOM1aVC/6oG33N7eq2bSXN2c+oKkOChWO8MtHMBEjh7Ut4J
QcYkyJhfJmkwAbGv4Y0nMZ3/+rtQmyCp3lPOZyfkrjFgQJ8TagTt59kc6ei2O1IvCDwHLx990p1G
X8yNijqi3Fq2wXQjXynASea33iDYxa0QreJuu634mwJBptp8JnrXPAo1Tw2JIfCoCl8Ng9JKty6C
2XJkxrklewJ34GTlktAUa8iHXyPgeIPKWOh13wpqzd1CLg+Rtn1yeG0uZJXM2c1dEh42JFZcwbit
VKqobsJFNwgzhsWQ/WqkvtSjnKJHZLCMfVX60lfgHSHxCDyQUqxv5PO6/u6ZrLbpSReNG07B4dHA
vMg+3ABLz8eWsE6NcwvejjpmDr8pHMynCqDm2IMBWT3gvOmLr9ptmlsE+H9SdfWrjF0r8d9sh2Ci
8KT0eO5Qt/+8kxTCAQf+mhUjmhUyxqw2B+TxniNUEtcsWNM5wUgbyR8icliDJcRgvSx2ZFA/fjos
lzP2QWgk5epp8kEanm4ZpU45GqvZ+sfLJssZIs2uOootr7obxzzr+tPwiami+GsPw/N0OrurO1VO
xTxtJ8nuU9Yd9nZFkRum7/NTVFKL1ihZeY74AtbncZWzC6YbFs1lAIxPI+rzkcEbnmmDqZJu9X7Z
hQcwiXgsUTcOsC1pJjy1U6gBTk6xMeBzyJmxz6cjgaQg4xk2+/xYmMmFaibg9ZPfZhndvTsVgWxy
HxJpyh8ocoExiv1fad7ZiFRynSFjj6rqWVb80dB1Ni3iqN83dzMO4EEYtGKp924rdIEwuqjaPkxu
6xXjV8m69/bZRyLudhm+Z7AWxtVQX7Xy0a18F604fG7CrAIGtlUYdjTsRqThWeH6PgtEBzvbtHap
1iP+RfJDQgMcJ5hEqqn/GQ3kxTT84bnvnoaxxyL0rw1hBFb4GRxr4T+1/sZ2FujopW09UKGQX/5x
TVPGgeJ9XCgSTFZjyvIHt3mgObzcgD/SvPETCA9bP8SDrjRxPIq1TkK4n+hpHtqMjP3p5PqVHcyO
oK/c9DBsEzc/pRDK5vpqFcJ0mJPgjHY+8E+sZ9Zb+2OMVgP3oF6fdqXsf6nURTp5bGzo9Kn02jJZ
6lVjVTFDohkutVMg85JZWg7PUYcy1A3q0X4FWf7vBJbP/mHnlajLKLWysKqDRYS+8N4HMMcm57vs
l5z3/4Xa+esfJ5BshO1C9uarrlAjOvsie8MlqAPFpd8houlPjwVLI42vfnrV3b+JeW7kxfWXmpZm
PAFaWJ3AJCRIcJd7nK2GVCGzzN/Es6QqDV7IVCpkhd7V+93laHUWPy8QWMU7+5/KIeS+kZ27+yNC
RHaAjfV3aUC+9XWe/0V1f+6+TEuoF4K2yYjpJEzgvfFYSgk1kWaO2MNE+8VBo8VZP/jj2+3BrHdy
76DdtiWE5CmLHvjtIcNzHv6tTML1t3wYBhLHDvjCAwWbNdyNmSEDpv1qdEAvV56AMdZSSQeZmF0c
owtSe/9VwzDBaMxpEbCoI8yB+BKbXmgtstTc0sclZsLNo5BH3LouGpTiTQxjD4gSu0afkEHuWPZA
iELuJ4z1TdNYAbjYqvGieMRLH+kgp4fRmtcwoo6IUGUbgFQdbQR12krt35ZytCkz1L2m8pdkhXGf
GrJOsTqYOjao5/LEKLJ/9WmiY+aADQHmVGGM02G/lLMWePVTJMtlSKzq8Hh13qAv9+SHNl4HaqYw
H1eMOyGI1YhFf5G0erULbLoOiGjDekUv8sBO0wUVMCFtfOsM/Wu9WHcHTu+RG7YXEBXf97TlEH1U
lXNQZX6Hw4i8qaXtYDJcYQ5WVuy0ChabJn2cAHKVDIITmP1VfwwwBCM0eKX/BR8S4cXx5ty+f7jg
nNTkS3HyvQl18FhW7Co6eSqlbN2x4Nbsbs1eTPnsRYyoDGlNj38lGNvw6woAtlDzFD4V+yFv+b7R
vqBTAUIf/jA46SVbm7HcIqti+/IqlEfY7kQJ33knPaLdSHRf/ya3Pyi6WuWIv+w+mq3GtVQS1OcK
/YIsTvgMZnfLYuAumDKhgwDHV/WyCZ6SLgB38KzwN1a9ZtC9GlVAUHV0jTfbl5Hsa7XRI/fpFbeS
VjQyPQFG7KN5Fj794QyfGj+Xq8gP7CG8hpMW5+YcOvGbRfzoByRjNCmK85eirVJGoq2dz3UW8FTs
Fek/tldpaBMsdGPyMRi3sMXDfRd3FHxX3ic5H1Nv3bbqhRjB/nNLtGFcgKGLVsBNueFFbjWfVxoI
x0ZkrvWcoIZbu0nKYocAgRCHgOqeBQ965r5RwACbjadBaQIENKbFXxGXVLCs+hMVZvg5dyHZInjA
X0cUhA1E/Hz+5u6wLttNlaIJX4Hp+8itRk6GGPe6og7CQKVN3iRiqiOkPZecJwxuUHnif5Fl0rRe
IYKxHFfTEg4vi8J9Cn/LzUU09tzmNxjcXmXkx6in2XcmndvbTKqESuqeYIWmJO+YcvHnk8qFEiDu
7UnF/yL+S9/MddOcLpRaJjJN5v36sQUPRex+4QTQWrIN+iGikS038j3QvuDxyL5yN9/yk0oyHpRH
+MCmWwXzFSAfmm8T+pTz2pdqlXK3GYLKGB1AAkITkrcjC1ufxoVr4q4D34sWzwS8K41LB3hf14dR
wGevENTiFCidDi7zA81FhJOlM4WCSX8osz75qjIVhNgxhsr8f5r+jK9STRQBejWryT0eSafYflr5
YechO39TWEYuABVDiRUW/kRaCjBBfyLLnVNd1zC/NV1Z8hrnMkaLWQTXIzl07o44SiScDpTS/iDi
ClLh74pIYfF9tJr59e4dNFeZeWk5mvDajwo4UgtFD7dFaRYpxGgqjuSJ4dgGH5oYjpzRjYA4qVbC
eR1LZrp3wp8w1bfFNE6R8PzNrI7xesSx1Y58tGRu8JMs6rwYy9//30c3yyUnigUsFCoCElakTlf5
jh9qOYA9CQBRa3HFtoDMkxcDi7mNoHMW+Bx2NTP8P2v2NQkfprQzHQM8Go1ZQdP4r7E8SUHcKGqV
qf9e87dZU2i/88tKtrkOQRflIdksR7LRXC4S+1IMNu6yf9RWN9tobAwUC6QUBiBMCY3xlQ/o12ts
MKIpTWtkBxm/9a5yMr+jcwDK8WSpULQDcnbgcJ+ZIuQybbCNU1HuEnn1RohrdnKqzHe4eQKL5ykb
o1FCzq8Gmwk9h581eRgAorgPv80s2uYA5CTWMwsAOTvQcZ7pRmagL38cfDRf+8FrB+mWJznpWE4H
OjDTf2eU9hldYW8suDD03nXZuHgPFJS2HGgIUBavN9XjlEiaiYZEN7rTAwn69mIvYcZrDjCVHBRs
8kj5mBDYdjc8J6ivHuu+xlnjuzBhs0VRFx2V5ujbPY1zEXMuYN/Aog2F3KwNjDXWnAj0e5q2wD/S
pOQSmOd4dR+/wJ41vt20nS34dzxRXihG7GJ/qgJzfcBuXfgdzdJSbOmFrHLuHahTxiTpEnB8+KrO
SNhKqm1uD/RJFRhEKwLQEoU5GN2BP1zG33zcU5eqS7e/i+LKt5MN1NHVqf3+KUWRvkSPUvo8Inqr
IxXOF9yzEhSD6Brx+kINldZx2O+kluXVhLzqybC2UZqJcUUjmsHghrnTLCfyCzGqyzYyVDierwbw
TuMbtQVoAhuvVvqHCRJzhVa+TUODeB2RaY5xGSvTR4TGdFY1Vyl8ppNYo6QY5egjhWTklKJY6YWf
58TEvKdUa9pvK2wKG3dIJH/EoB7NXCZIns6ZGYWt0SMhFI6qO1xHsCLiZxxYawkuP/jrCk6aY2ET
V4H7tOaQr3DT9cO3lHTyx0SMY0XSSZX5QiuFnnANh5noFYgAFrpGI1ALlNcQx6568OCvgTCkRKaj
dZVDbGuU/yFfKQ69bkMf0NOYMurznxaQeRD9Rm7uuX2b5fUMpqVtPMd3tJupw888PRcznxCeeMj9
WWXshOOWTaT93lLuzgk1cINOUeTmgB1fhp1CoEANkm6EK1dEedn1Mcwzuup+9TV8EpHkmQIpOytz
0QT+Mq4FgpX/f9r3bFNabCTwe9nZNfjHPztVO3aFdJSjrSvNjnv8sxkxnDBfMzIRTSezijDIlGHH
1NKk2Fttj1PkqNsW4GQ4og6ZKSB0OoKSMbLAUuPFH5U2hfkXXzUGdDNmTvk+YZBWGeLrQmniFR36
rFrLGS3zn/tnE+66rDc2eg9kL2zUkN+rtHQjqCfBuJpNvUxxeKCXi9oEjxTup+fPHtG6OgGoRils
sbWPhJod3fVR82pvyDUOOL7h5xYLFnHVBrDd4dUCX1fnBzyAP25jsw0dbPxkp/dgRjJ/z9Htlgys
swXig8wYrVCXeAwliZtvzqh/h18/Tf6dWFfSe+Xl6MODoIToUDmm3jJS4lmqzpkIAv0yAadEfili
JwcrVEX1BTL3nRQviMLf/UODh1fGGKbn9+Lv2fmS+2Plfzf/vUlB4fRbFjdTZlRZYE9i61UpPYFu
Hvw/KHdWPcASNU0o3xj/BPoTP9ehDzKa1o3ozqPJnKN6zx1HLU31pzKTLSwCO8njGwV5qB1APDM7
vRTwfjKl0/q/eY7K/KJRE4UqtL/megNEMw8PWK2/dh6elLEREw0WGAQ4Yx1VjrodVPg87Gnw1Na9
WljegcPMiyh/9x7zk0jtA+ll2pXY/fa4S6l8h1LKxR1vXa4E79+yPVShUhnjCGv9wpmZZ2ZMFw4F
ouSFP8IReQRqQsP2Lq/SrAP3xXlnx43ieC4P9nlapFRYbC5sz5IuRjkWEuTe6tD8tT7xGvfPfVqh
5Xe07h2+NqEItC65UMDMbaBHLTj+oTyp2PgIYWstuWqUNtwCowz5KXBjSQmQEqbrPdGzlsUmsV42
AehrkvdasJOxC/2BbGVqrMaTlDT2hjjUWYun4hsuIgH9BILBSts4qiwe5sPnK+6KzE+yXzrYAi0B
kk+z8Gly0r54eKPERCZsaMYlN6KQNskQRPnNZ3+YThWgvqPIRCwKH8k+Ono7gzmaXjzvZ8T8ylN3
cPmwQYnvb4t3zEFKUVkXuCBIsYtiCAmLxsZVM/w7FpOleSNx6toUb5Q3J5b+A8yilhrrwQ0UEm46
NS/VIaW3zNkCKpAfF3AToB8Z6toB87BtAqHhUW1Al1jc6iZBnGpNHwjjCP5F3Xy+jRQ0GI1pyqRZ
HL79CguwAjWJY3k9jh/mrxQCJwapsBoQD4Ssp3Mn2X4vFE9/oe1bho3wqpuLJ19oPIh+Fa5BNZfG
8KRwp7hchL4gw+FHuhbVt+OzAWyDV9l11dc27SkKMwgLQUSCtAh+eSytsWVz2Rd5D9zcSXhW1hP0
EZ/HWW/LOrvyqF9QWYwFiwkp0QAuBJneyJ+ukk96X+omw5AOokScS1SJ125JiAT/AFKGvb1zSEqj
rZlCfLfbumOruyCnvzi1jlFlivXFZYt9o72t8xMj+o5vm91wEryL3TAKkfVJTdcn3QvUQWK8R7XW
yJ/5QZfZHW0/BvaDHfRTBAc6QxoreaweFVJCsPHKPjhEodkoMb9q+XFNCTbOV4cgBLfmBZCZcZ+W
l1QAYleh7ny0FUFrdqDiFPHuTXEMV0Hp54rFGcNQ67zlklQYQxKT9d7zaB/3fAIjZrtzLQhxq6h8
Tqd3hoB59d5xvAK3CoIWOIBYB+u8DkQH24PNX7/D9MY4BaVpaSo2PrX+ssl+yxRfdDtKGNYKkgGt
n7w+giTzKFfmmYu2Qs/NeXWEHpNkb/1y/qfZC6jehF0oEBMtWcYMZsVWhkNyldE2kuH9SMtCcbXm
WZV1R6q8ddoocCyRZAHTobg+a41ra6RsRfI1N+6jXL5B6+dGqmWBB6NNfRnAB+XFT71ECvmImbec
vGUTuDsgjWAw5MoRiJe9bXcEzOGN7Cj3VCJ9cvOmxGxpEI353A4Oc3aI2eh+vDvqDTppFrLHIyYS
gETjjIL2VGC9rFNzdXoqljExkIwVXr4rMIsEFqOmtZkbo3yWJngHccUF0oM8w6FUlXp0hXks5tsk
NylIRfqecySVXFJESTx2O7Usuu/D9Hz4wh/f9hBqBpU0uL6/WcmdE1YznOrHlX1PKrbE3578x2xl
FDNDgyFnrpfLhgJicIYLDA1aJxulWibvhxxRXnmwl6ET9PV3P2ShjBtGwqeFHqtOm5UJ8rKmWg/W
lyYDwRvKkuFNn6BL4ecfRonUXuhr41nHeMWF9iBefi98K/E+ofBOw9nAe9BTxqVotjtKX7W3VLt+
zYV1VKr6rYDtH/TD3nIvJQfR2ARThWuGGcdM2ZBC/DghMfZpvUsOxtRBK30sg1ePnO5OKu8rQfqt
pvSMK56Zui2Cfh3x4jpfQiQNiRoaDPuDxoTS5cxc2Qb5EwSo6TawIZHsQGC4obqDbEx4hbHUFTFO
AUdJkDrVX2d/ceQEUk1KpfO7OJTxnc6r0SHs23lbhmOXBymUa0z2UgImxdnks/+7dom7aKoplrXN
jjgFtZohC96OP4oYB1bfNnSjbf+D6Foj7taD4HdVWTgwNe+fcQxFImhqt+PZwQuaG7/vU6QFFsxM
6YjuBEngXoT9lAXZyD51uNaRFPDxyyyU2L7bjbCtRm4PHdQCmkT9RBKdnz7hDIC9WPFxxnm0Ufyk
pXDzdERmmHK7D/mv4SL2KwD4hfzpr1VYSOSPzscbe6MbRc7o8eoV2V3mIXLaUFKw8gNar1I3Ixnf
742Ev6oZzq4ZGPYhbEis3TYFPXqzSFsbfenXDtDbTtld8hK/on1b1r+9HH0oebl8YEgXdltFb9tX
T5veeX59gHD9EjY4n64FesGXl7+FUTz1MWMCKEqRjFtsWxqUuP1oifUA+riCPnsGuHObD2Mtt5EX
60AxORfgqUGVfU5G/zHQ5zgRcDxbNCHEMOX5yb+rX7jHE1ErllS5E3B9Rkx+LFyjdojtNUXmCx3O
X3ITFjmZDiFRHpQG9pUFFxSIUvzSg5Aaw4nMlKBhoHWQHWVz/Zq6BVuUgEfK0MsgscUsnKlybcPX
E6uQQGFuYMRfK7ogOt89SoQ7zFh5+dteofqJgPfDhFoZokNVDavcdpVVlZQb/PgsKsmIIsUtkQk4
sMXYtgL+4w9zRCXMxjxx0Eyt0aiNBnkvx8qjcoRTOwATmCJXFDzuudjKBOW/5hPhB7wbzKMww7LF
Mct5k3OvbE57tKHx5P+s/RvC3u1xd9dgaC+FZrrC/JrwmnjMXKe1BWbalS5BS2i2NGerDwgJn+zq
wwRoC1h7/FnQx+QqJ2GKoDOYtrk1tcBUXA+wy3G4/Bcezonh0NGfZNLNTgHZ1FzvuJGXJ2k6BE4Y
SAoudr29hxSwJMoNUbH/Wxw6TiDYiPnNqmosTK8g5U3DtjdGbQJfmuWpxzdblg5fr9BfyG2y6N3v
FUdFOscm7goknonPNAMUSKFBlwX95BYBEMaSmk3n0fvCPWP4X1VzWuguRv7ns9xwjfYrerd6mjYR
ebTT3wyGLYAs9wAe//p5OrZsm3DZg5HGtO0RJpu5kzIYzCQz8L4EjL55gcS5e0H8v2o9FYHHsBE3
auobYKF2YukQPj0JC9bPlZYQ2RuqdITxfL7xN8IaPGQ7gRXDlt1pRbUdYMvmmRatkueFTMn3gJBm
JeqI2alwpzAipHPWKCjn8+hGDccd0k3KN3vx+DvDDNM6KM+9s4yut9iSAU+qR3KJ1sLnfZc33oI2
XODt42+ULwKzEwFAvyAYg1El9GS6Ry52X98cMi4q2RAkMQKm9UVjmp6PCUNG6IfIEn6zheW8AHOz
aLu/O/GeDcxj+Dat4HlfTOV0lmpevYs+IPEjJzZ0meDWIchugkgONdGdgdKvOghyAUvf1Id5ir9i
H8wq8i7LKIW2F7ldwZjvB4V4A1F2Zxi9wH04XvJVvf62uFyMWPGmajdKnthhSjvxJJvAIwmRoUZK
gB5EaFwx6sw4a/YKjN1qMtfICA+UsmNlfvYBVi0qkHQNvisDByJkmcxHhH6mEkYnONua3L56qY85
BQbA/I6bLD5Uw7KgZDvOi/yUPejnAPN0nzGd2/Cc3/6ErjewLS1wsjwtg/DXOgH5qALJfs1XbVFa
rA9TjRItKa/C66fN37Ip2VtwmTmu3F3rx2mb/C3dEX99RRH9y0eX0q7feSX8HI+EtcYM+0NHdfvI
T3PKEJHagsIc1Kz+qcYjmM1uVSSEW0b3QU3f6kT1a8ODq+i+1ul4Z0gcq3kH/bPppSVZTDHq0UtM
mM/XH/YnDa2Oxg8eWQrICltaAes/694vukt/tQuuiqEbVvsphZqYg/J6ncNK3MtThc8k3Jd4cTir
oB7pCe9Sg1VDDrmKJulkzI5gTCEipv+l9sYgBTR4JC9ARUFuDvSV78fxZuzplrnw5lesb+s3dZnT
/AdQyQ2KaQenzArVxQbSsh44WMsGTVmW32/YwwpshvBNyrQn5pnhw2GwL/2QXoETdgvoe7WdPn05
UqlLBfzpnn0lGwjN/nz6YhS8X/71McfiCabAnSl5DxL1Bisn9hA6RBEwxwTgOTvFk1Jo/wyx5b6h
YR9zEWQ7tZLXISdlTxn2hTfVf0S31lOmTmoXrp5Oj0CT9J4JIAQlhuOepzDtRK2nu89amIBIkDyK
3W4/yYUH061DFIO8KAOGx0aUkUEIl6KWgNvWXopGFW7VCv4DdtgwqEVue/ybzRhE18ur94eEgt6n
pOyushZDbFwTahCLtswNRjWImvy2l4IYopvEjjSsRxdecJwlofMBHSlh3CwzqTJH5ONHsZFKBDk3
6VQwrv5hNnbkQ0adcHzV6UAhImJlV7xk97yqzfQY5CpuoWnx8drctWL9eOYWQ/l9Xd+byBAC2aLO
S9BQEJ02bUbItifcaqJmvkwGKTWiC7v9oN2wezz2eb4pUm7MpDrZ1JDhllIKrvZzj32JvVSLFY2v
AGiFCV0gdVB+GqKLC52dRcM+Ze1YYK5WbS7g1X6owpOCe/TFyurAPmkQTjSA2jGbTi20vJkAqwQ7
ifooXf6cVI2RQqeaRRC46YbnniEKDDpXhmwkDgl7+5WtshQo4JgudPFTSy0IB42YIpCkuPbiGWvj
yJ5Sdr6e/jpp3uGlSWFQdhvEEBRUKOHptxH6fP/Ak3yYZ4iqyFpaRq7vVYRwflc+mr4KhWZcHiWP
Tr9/d4TvCqLxqvMlv4EAa06OckdgH3opj+IfX50Z7jVKHTowA3s4UbJ8u5yYzrFxdWBTm+mQFWtG
Mjzlor/0Z+lzSSfQRBOHI8KF6B+SIu3Wh/4bKF8poOsimI9mDAhDTSM3IIOvZuBkU+r0X3BYSD3H
E2UuVWQm5FGWJecDy3RzIOKFczdyDYW+Z/iOjfLl9bzliuabGFkuwzpxqkZnQwf47j5Bg3JCXLSW
qtoswCGwv11Ho/pnjJtIlq3IfDkwtUtOyySg3gB+ENpBAim1knbzxFPiPusXCoKDPEUD+MtjFGzC
6IYfbcCzB/bk2DkVb+JOOc2n3sWfXkNXILkI8C8O5XzDWlI6N43ccPzhwji6X2tQ6gX6AP7ggGue
HyIT6gKRWJxDxnAApj+zb5qONI+LG6lOuev/ap6FXBVCz5A4Mmg+uXfMIRkWWZbvsCwFkiKcKjG4
uQHU7KVwmH6YJZxOIXgR1LDUySBlsi5KBEp6dYMZSRbkjf7Mdk/fpT9cxnV6n2jLOHWIZ44Ic7e7
pqDKihGyaI6XsL7y8HBFZ3XG1ZekV6SxiBM+CvUtJPVfIGsfkaRZaQHjmzYduhP+Mi/FEAn3wYPy
5+aBoyjavoj7fA6gmrKy1MBbaSo8MSOLPdtkrYS6jPsd9XKG886qiu2/m5MdWPva0xT6ix/CL4bI
/TMb4aHllmtgD/RIUy9czN+B/5FpmrB5gXSRUIaJiTIZCqHrNpiJvlCDrjogJwbF2V/ds+A9033E
9qkbo3mSnUaDtXT9abNCRcEtlU20Om1eV29E/QnGPpJi9t2oOE7mKTFQ30FPVDHKzko1IzrH2hU9
ueL19x0mrvnPnjqxJunK/VpFvXnVhCm9ypxRkqWl5V1mdlSgEjk10Nx9EQf6cxZejEWvcltlWKO5
agTGvvc75YQQvbV2SBQFa4wsG+pg5FPPlLzpaAbhM2hM+HPh9bDz9/zh2K+LORkKw19UthzcopSn
h3UvLxP1TZtfi5BlWaN2ZDCCtlZ5wLarUYSiTwv1dsJmNGckq/KScQ0dpSOXnJGoh8UMvxSVZY3h
MkAsMQD3GDzqy1XaiOMUw8ZXMSWIL58sJ2oQqBexjx1EDLxls+HZ9EfLO0l2fCL3GfP/7cugfMG8
j4K2DIso1aZzHqLqC62HJaR06cl3X2SK44GASBYGZI6XXwsxE0N9fPoJ7JunPGaov3rBstquss+9
6mhZ8/4VvvkMyv5XEXfS5FIupB6COsvTGq6PMG1fQb9i1OaE3kWGlniQnxXx8gmII+qcLyANoNX9
RCHTjRLWpyRBlXocVMmd0SXiBNyU70Le0No3PNdmlr2UyofyWCa7hFiz3E/wF7dgF7SuC8GyZtIN
cHhtLxhOhmfAl1OOjFoQNFDGr/OdO0PrfJuRt2So9MFTvLTtK5utE+YHMfxA4kTxexK6N+IKW3fv
PVS4IEljRW3FK+ObuB0/O6fP65zt6c4eXkEoQr9XE29HLy/6gV7FC6niBWHWq/lnMp8ucbg7psg9
I0BDW3e324m8qsH6Ak7k/Rz8fm0LwV8lSGCVbDI2whAqBG+34kmooKvvkKh3PIDmQlWyzpQqQLIW
3t1AWCumCsPphEqJGVb+sp0AySIimQS0UUUb9cd7mazuy5O4vK6dqPnBJ1+O4tCM/CEXJ0BYIwnk
Q1hKS+cwxXIkbdB29Zcx3YaeBMvYwoSVcU7Q07mBPK7TW/3gszrOJYXhewRCTtOD3iQgKOm2uJM7
9RiHknHXxtt4wLn4nBZY3I4Yyl6+WhzgYyJTNIcm1gq5Pr6zm/vhOU1Zf2TCUqWZ4R1PCn5HQdAt
JSWk57JLbRU8CYtLH02TTphMq06CZ4jKP9jYcHuU6q9rLtBQv4CcDZKwlttt4O7JJBhAuJcQCy1H
f0ZdLr+eNPpOJkKDrBTBrWmn9Ey4+oLujUqfiTDUTFuHREE66uEwMRKwG6Ne73xNAOzMiDp9MfK4
DkmvALvCaVOCha0uwjKcKCO5voFq4TyG1pp6aaRCHfGlrXeBr1R0OABUlTW+IYfhRjvPx8qa5SgY
FfAtj1O6A2unBw2SQi4l+T3h2P1SjFKJtciHPJESM1GQ8i7br8Eoo245jvPvvA/lSjdeP12Zulcy
fiXxR+8ws/bX2FnCbjTalz2ZO9PQq+hpm3+gP0qwrMHrpqr3rFZC0DpWHzGdn2FcUaLv4sK3OYts
3wYqvoaOb9pah26ZCo0bcfQLopMMpYngO5qV7eSjcIvSY7Kl/fJEeRvxSzLmRLCbB9HJrx0o2Yhl
o7uAVJg8au91+IuJgUQ8GldTHdY+3jZJt5EMcW1nss9bDPN2V7CIa4rPMkHzfmmsMbGWevFUlRtm
lm+km5mXzn7g7yTYeSW4qIiLXxP2YUqu+fAJyHrJ1zoIOJR7PfmIQ7lGzIZOwWqPWBhI+zSkYZ0I
jEx/he8wfGN6heomUCGQIpTNH8nxyBEysAxz2+gZ5MUOFF3+FjyQnam2sIMvP2aCuu8qz+mOyZOJ
S3IOFkAslIswuHsQnj5AEqnrJ3CSyFX48z6KfoVJlgQ4ufKxeMn57OtHg/Qa2e+J5E3u2Z8WnztJ
5062EI5OQSLq2+0QDmzQo5Wx9NaICNB0OtuYWQmB3ffqThxt+83vzsORP+VMMtla7wJVm383Ovqt
kLWKLT4a9Pz9ZBs2B4ll6ErudEhRJBz2S4wGkS12DF6S2QFfsV68N9fy4/Eym/+Nj4bPE3JiTc19
ypQ11csmqvYFXD6JaQXVqHCkEqB+BXXTdthOoGtwMZYUyTSYm1+sd+jer4ctDs05Ixf7hokvkxVU
DeTsCAM+jzibpIu04yMs9ySKkr7Ou3SSsdiJ14p/gE+/j5aXwu4qFrU2aK1EoUBe+qSQ60E5eLOb
31QN9Z7jLM2Alian2M7ZVXkRandXJ77lEH4M7ejDu/iTI7L5iqx4iSz1i1dq0aaGNLqTWcGflHVJ
ZniMpotBLUjcPOnd4hq873lZG4I5/fQiTAmeD+ZztXUkxbBvoFks0HqwqNm75hxd4g4mfJxk3wIe
bP4NnVL28hfRlf0PWpHwB8gf48U0+pt2VOw5jCgT/HlICJjLDA97GMOJ5oOpVfrGzqPtFQFChfxp
m7ja2CdH3ZF0DGV9K+bSRKDeaSXY7JNPRNzMpMi90E2YourthXrHJeYXAJXLhhriGGFHImzvxWC1
l2Ds0jP1s4UxzK4/0j2LddccTOZuZlCs+8XolCQXO4SPPwgQHToO263GPeHLU8NqmVsBgo3N4XRQ
1gJED8DlEBqrHIBxgEQ/u1VDwokID8t0vQRWDXCAm8zsGP9XcSPaSgvjTMUG3gFea1a3plOmSwD1
s/gVlYV91zyEqBrX+qyaY7z/lldvMh7vhgJR3tOSJXo4SByAwShbRw1BKaiP6Rqio4odN+FETGb1
YasAwv5KZL44WRoVORtzdR15PfahIMNg55SmSWIiXcmE/Aqqp/8x0x6R1leaBeWV3WBfMw+6xFmE
zAlTAF/SHnjof6ELR+eFBSEKen4FQv9LXDSj8Ult/CA0xqR0c5KgyJ1DTv4pkOUrJsHjDGJfwOcW
MKrn3XSw62sQvTFOmwUnaQWd1va8xZElPo5hIJ66nhy+bFLG4tqa3qrm+uuZIeGNhocfPQWeueOZ
0l/67V+N2QXq9WybqhlLE1Otk7LEzsxl5gazGClc9VnEi/KrCf4dOj1HZ6S7mQ9ByJi4goBmlwu0
MZaj4m2NWI/JGv/TmF8XB+ceMSv2wlLaZJoCymqVZHCnuPCAjs1d+zedbWQ3V5Aj65YL/0OGQCj7
SMcoj7aKfTaI9N6u1a/9el5nlo4d+KsvZ+hiiGFd43IVW3YRiDUyK0zN6qcgiHVkvdrWQNvTokoM
oLLeNMX3TG0wqQMFJfngrCfGUiRnFVFhxXjF9MkhfY94MQPs9K6IDo3kTeLUKjySwc8JmMHoFxgS
6aCLlxZstJc28dAoUqli2vb8tt7k60aaAj6634mZ+t8+t2Tiuo/GR2lQ3CMtEeug8zrP7I/0Ch4W
TGm7aejx/VmHZbXtsnyBfjp2kTUDfGwYgG1V0knw7EjgMpFS4jHPODZs8V4HJInXzIzPD/3CZ9gM
jGiJVSEpCA6g+rqKlG3CfuVPxvj6/3tNVNw9A2J7EAYp1JLkvLumIziLGliCB4c+JhSbvzQ08del
bgnSxaOmedct3c4cGJn8YFufkgLtjP8PYPJURwgg0ndvyOuIzK/JRx8NowZxQlvLUe20K/6N942w
cIkk8vDWBrdxcrSly4mrAQPgO+VPzlGg4SbqAbPb7M10HbImPcWVfVpBVAk1L4bF5yhUMJ/OzceN
H42iboMUJPWdSa2O5FPNIZt4VODKFZy+1C0+JTAuH6gUCkiDY0/R/3Lq6gJml6hEKppovAcJYAjm
5ITAvCOd5PD7mMZp66m8Twl3ueZlHyQF7xB4UtwRnEd2nf5MTGq1EchlwpiZDY8aawGbDiHHW7q+
wRw6relK5QxtapwzNxP4I19P4crzTaXu0rmSBTJR2E3d0AzxD52qCw0Clces+WmzWa9DaB75a2BW
qlv3xoj0JxutYza1EQepCi1/Bu35jVw0523NBHlNtVzo/sfB0ZxKyBBDVPmgmDWgeqX1MHvxCl+R
ePHIWUGylf7yhizaLXwn9WWiL4G61Pq8pflpG0xB5Vp79JhlK36dzUVKEPEY7SeSk3xed33vvXUD
Iz3u4+pW63/QwdWebBJBMCHNwJ6PZoF6fJIhMMxb/4lnZygy6t2BMd8It75Q1bEVLExKKYvFC3ls
ua7Ird/ZdDq3nL4JdL5+GsmAh4Fj+9Z3/K/OyiHQpPetQesJTFcUOpNf47DPDvQytkoUXACAKB4p
xYKQtgDargXyWk5xMRKq3479K1QswZWQEm5Bcwm8IjpOlG3eOSNiA8sWJpNHXE6oFag/Q7kLLGYz
1qLmd7NnAjOCrx2N6KSC7e7Bfkp+FrXDx4kbzBmYTJuxbPR84jlyceCEnEMXyUgYNSHUkRi22Dnb
YPih0Wa09/WibzdrxmeYQJrwgg8v3xaBa26mi1GdP3Y3El+qTYr9F5/JvgrbcHq4fkQNck6z63mN
pO4sTJmcxAQjLx41LlCcJjKozC8QPnj8QVWRaaHDye4ckEkw+39io/sPd1pdYVDXgfCBKeGasD3b
uDrwqXt4uYCloGLEbPD9Xl3vcsGzaZh4l9kPu08kCGBNEHn+k1PVwTPnONbvGq6dndAU2FcPI9Il
9BsmRGdUqWV2Lt+JvwBJe27qkbxOh6AKXsXKLMKygRZ8u7WrE8T+4ydFeWaPsjARg3cP6p12Trxe
3pDPbNXhndVqDb1zKlL25pzd5dRDvvKByevP08ewaeD06LkUPQzq0qdNT3c9lvENpzCZDCt5htGL
FgjXprthG9EVNdVAbL6zudyy6JTOGs6MuUTIsJTdtcthMMo0Fcwc+f0e28rdGmHoqSsf67nhhiNs
grKg9tr9/5EinHrT5itMVq1q+xsxXEZgd8m+/le7U/Ro195ezBcApMH3aETmvhs9Kwjn4BQ207aD
UcShhe/SdiWPBF0ltxrKSa5fzIKN9EzUtXr3b+dtxLs7XR3i3lccvLGkx5gF++1563opbZRT04PJ
35ykMNk6NaEcnFTZTAq+3xfZmIMwYqvyLlAVvXEljySmPA+JrMiYedpEe704tsFgsaqzPRrLvTR4
VfjlqILByfvk0k8WIa23dosZ6uGHjq9smIYsGrjTVhf21gX6CxdCAdocy/IT5bIjVz6DGnYnNF0a
OjQboOZAlNdhTdWMyLWmPLw3Z+TNV3jvqsF4nWtXshxSLmtTxSVWggmRtMXCU4IuI9rcNhIS1xVs
1K7s2eExkbSy7sDR7xXPyK5c8guayJxFDzXAAneoJHV+ygYx615s8mBNR+9kAcoMn+h8bE9NmeS/
OLIjbTWRkgP1uSXkh61XwSJdFW+tjW2hUTlYvs8UVtWt59zui5ku4Al6lsSuq6esp4fTJrSreEgf
6T9GZb/F/jqy3c8+2mQIWY1KFLUPuZfevWUwCboWjmMBLb/43ps/pbO+JM3qzEPiodKckhCd+55i
oaH/wy58/nYGwwpuZXMEXbw0ld5YSmr7PoRd3wwx+SQpo0ZNNnwB80nXrUrgVFYUk9uUUIVawXrC
TDZ49V4B7ZAdSms8fvsxRKCxOxRh/NCPZvMDlGmFBgddV65c27OnSyLa+V8LE9esSSrRmb/oPikW
uerdq4jhKecW/DcSWV/sfFScOZTxSMOHzbnGR9mgfPLRgErHP/LiHXuJxI/hNv5xNJZIhZm7wt9s
VsWdz7uXkbK9nJd3Xz/sVpK1B82+ifEYrdvWgxUgrGXvwTfQt15NCEpe57wET/dWhlxvknKSlEfL
RmLvmkvfVHBkFV6I9MjEqHLP1HW9r7Ffnt7SS0iN3F/USa/2PZBcm/G6p56YSCxO2nrmU9K9nozf
DiDdoAmyWqwkiBlKz08+m6AybIACXKO9dPihdRIRYJmOeCu2L2CSr/WnID/vTYYh350aayusauGC
ELjfqRPe8DqCvAiRFIlzXuA0d/7vxHZ3apFaNyPQ6VhWVx9r5xIWFqrdifoTTF3KnWnezks5hm/X
oon5NM5WD/Qn4LhLY+BLvATYmFuumC8hmznIYw10dnnhqJ8e1dsbiFyxYREq+7jvhbulncDF3xM/
Gkfk07F1fqZHtlhbVMhstRpCQ8uLogkhVW0Ll4M944GpxSMVJlTiJA0Ldj0/SFEC4bz5f465iW7n
ljfW2acxpy9NK3cB7c39iVhyPJBvP60lpO2JaazIeddn0iAl8+Iiecg+uoIk90xMxoCREaJGqzOL
sFxQkNvzdKVn/ScTKmRNfEy+vbIYsCzoQHs4ODMtACQJsreOUWsREJb5OWtuyGQt5986jsEMWkbt
Izuicj8BWTp/p2Mv6o8dp1JJgl2Ly99ZWFQfqc8b4T9X9or4RVInv4LcStg8ZOjpDu+w+TpaYIv/
3YXzcYt4G2taGYp4fgiB+qlva1W8yXjqgtEJ5Ug9tU0HtPC1C8ccW8nKQkSGa7hvaYIzxBldfYrG
ZZ6KYVfHzeUChIUtXrN/zsUFygQTL32kovWSzruTMJkLa1AR1uzFF2sPRx/wJJ9dCoccZLwVlgkG
U2S/I1iavqH1W9b8CvJID6REdQdN3ghcjvI2nuGoYDfS9wwWFAzznOIjwQqhiWSFdrs1+WR6wHvQ
lYz4dKK28y6+e1e6HCzfZYUjguQIZDzBFaiQjeREUx7l7cKetafCz48GlvoXw/SUsOBXYq9AMe7h
04UVf2nGY1VUdSvcJW5xyIuuXQXXxaE9SULIyBV1CGt8NM8q9m8kxqWmbPc7I3fIMGyJa9vzOnIY
M2dJ2KVqicuFvZUPqZqowWr/5V2Yrsk+llzNZuXGbmI9SXDkilsjvUIhbIIiVWI6Jk/OoNHGgQ+w
ttE3HbNXwrkRwdKs9hbWhDMgOQSyfz/6WduVtJB8IPmudpKkqkzokhVTE+t9fEuNgL4KYy90rPR5
WdE4hNjVmDPzoMLaKLVozAQ3lNNuFTbV720v8jIplkeC2y8m3DNQzExOZfY3xOQBrwQYZqrnKwpU
I2LqyHLHFUl7mOPOz37+dZZq/RaIdmZy9qb0Do+LdBLbHSkFsOcBkUiPA5lx153JxopbIg5JsrSF
DK+MqZUTTutPbQ2smnwkKnxVKYn1mtdmW2aj73Z6RCa1s8qFRJCa+yuqtn5An++7v0Jq+6GvlV38
/LoxcSRhlOtqkpGBu/svedU9+UkiR/ktfg19NstcDZvxWfkkOGvthQQRf2iRL/jo0xVYbBuP/wrR
G0tEPHGttFvia+TXwGsReOkFzZcQatbix1/6RbyZQZbkE6ccXq+yv3SatpePHzhH/ePEczakCxI1
tVFH8E1xR+WLxfbpkJEDWq68Jel3MzKCHPDUYXA33FhDIY7wlljBtsLJtHABM3M4wNnAz2P3eW2F
/yV/oVmvURna8PfheCllIdAqR7hvo2g8sLR5muOXydjuv9LQdMM1wxaGRyFZ2Z2fCle9fr0fHSjd
YnGXeXbVww1DmrVaMg7vh9Cjs7iC9YYth2YWoM7m92FP9tMWYoRz1A3x+/4tFY+f4PeSL5BzjBbF
V6PSzVq/Yy4oKIsbvOAL04nIwri/9HzsKXZHPa5wkMRDiRqpA5VY/pjq/PbiE0RK8NMKt5vclMjr
5lrBmKZ2DEoOiU/hM/7exusoIKvkIHHvXVsViJMh5hADkJZRUpsY/xsC2frSMGLEZEAkWcLd2Qlb
B5G3oujcR4OWcbkhX1pzhf1C1oZNX5s+ywfyG2t9rPjLjbIV7x3vEd4tKux2ZIhWq0gacQvvrTIS
V8wcKakju3FbXvDq/brjHHKeXNFtsZhfvcfaehFsQHP5FFFYsiw0p/8mW/e03XfmcJ4MHpJIxKWo
/1sl9M+tJmjDIuQdNavPim8MjflN8dmnSj/exECWvJYbN/qiWo1PRHYY76eFqfLu+O/vcgZNsx/e
Rice/JbZX9tQz+Iu9xIUi6CvZTdmHXFuvdnEQXenc560X+FnMez1ZfpAHaXtPCF4C14Bgr0CaLNv
ADoEWkL3i6d8xXC5jmBrFoV/SqHgnaOKQLJ/qkgKemlkCAQKEAl2HnJbrBQ/C2z3s/UqR+sJAVj7
1UVqTmFKvziGsTMfFSodyOXPOlF5oJ5lNcSX8DF1rtX1Tx5ynF4S/jtLDisYXAqV1jHoQy1C4BAq
8SFJu0lCnXZQGdK0lrbuSen2eq9CuiGstO15WvojoJeYau3r0Txe5XNRjBfN5DuD9l7rKB5tfmWP
P4jACaOtMbz3vcb+gi0X8Y+PLmbbOmsIerJJVEQex3Hf4tEfSa3wBiTQcwNWrprfsR5jPRreKeWm
J47jJdgZ6CKNodcF1Rp9Pjglmz8yiJBVUhwcAgEwkjlQAotGRpzyduPobMt2oxoJAuZLi7qGn0id
u1fpBAiqKGoOmhMexhlQhoA78Rqc00Fz8k/XGsdC+k4TZfWuSwSD8q4cbsfXtXluWFoJekMaztsN
9vQn4ZYmLRRmuyo3OcDoNxqR9gWLXBcITTdfNz3y1ikGYlRanOvwYS8jcXMLVk4RoY0IPDo+kmrj
WCSqNoZTnD8acZ/LqYjaz67OZg0OX3ERNQqr6iILNiG1J0MyPxZKXZfdbWt8bFRQsBTz6ryUxKhY
g/ZCcZgLsy+Tk6QSyeVUnvM4/aBPytiicvAvtOt7KOzqrBF35iJ9cnSwYlBvWvrLl9/vwKfBaI80
7zO0SbmAfRI7iicvDh+6Pgydbh3/V3QnMN2sf0h9RKnnvo245NiEhvpA5kAXoWF/eguv56abUH/+
QSXp2JwaXizKy08E6JoFwQwrCU46FWfrOFJx0sfFRNYqT+7pl+9ILoSrzb1OqNDWojsn7DRKZZN8
AVgDBZigowI8WS5YhHOyYabhVPCCRsRlcw6TWwMEesghxy8Wui3OwlLRW4TCPfZOlTZepx64+MTd
ag3hTezIQyWsgQHnCpEcnPVyeWfJeoLAmo0ocsXDuN6+JbWiTmCnQwHVIac2IQUHrZzyCOxUdpu7
XtSFRDsCq5LWPzgntK7kkjnTueX2lm1MdqpF+DODBHEV7tcxUs73u4RxXvScXcTT3hhnK4LVfu8E
FwApMqFeN+geV7mfAgPcG/eRk1tSoTCcqAZ8FJhAkKQoisEMj/qubXalB+Twratox7JmC1vS7GbG
qyAfgTMrXqnVKHQM69pRnnPDC2e0SxM1WTv4kie1EJdB4mGoAPYhbPQ0/WEyUU2MtIkkW+r6ZG1t
ruDNc5gSrZnYM4jKVD4RQS9nFawffhPCZI1E2YRvQQIriHOpzs448ndOUb9Be3+AXCM5mahWJx56
Ai9jFXMPMxJvB5eZleTx5/b8ZKmUvXnppSZbGVRTH51QqjDSjor8S9Ze9yE9v1yoXJ7vcejDcVSL
fb4f9r4iEAhEywKjeYQn/iUriUtdEEXn0DzYStHqh28H2EmvLnQnr7p3Q/5veFmdaBkZy/UnbShX
YKOZRDcv2HkA9a3F689MDfUuZWChXiWpxfSqnW0o6GCFitXVTH63J4SGHA6bBqVymce+ZiMVUjOG
TROgdTQLOW0+aOzItLuRIyIyK/f+7ZQ5zJeI+KDL9lYOYQrixePnmPJ+htTQeHN+1t+oiS3ahbKz
00A5HBk1b9nvAvX3WcDNH6ERDopjMnLIFbyZcn8f6lKx5g9OTxqF3ICZL45f9s9KoQVVaqBTyfoU
/axp5b6+sJKF4KHGxQcc8QnCITI+u9d7KUTW3StoQTgOyeEqFLP+o1Lz2LugoikzirsrVSddRML/
2rV5V1h3A7v2BKR8v4WZ7rZxQwSOKqwj223VejT5z852bTHQdrkcFCQuqnSkfYgmLnfsPCkkP7yd
NBBthofGtkh5TYLcq6zuwHL5VK6ERFsAx4vE9Aj8FYwXGMHlxjo/5LkT53MXmjbjPprQVgpEhqMj
S8LThPTMvPh1R6qYezhM0lxVOB+6ur6BUbYKn6a4ct0JR0VarTqhOWSHyruuOtpay90ihRSHW0Ww
uRBGddyjn5NEUiou3JFMrpZxJElAh4APKaIEnePIgrxbwIdXvKNGKqpDEDibL8kohpMMJNChZSdW
8eKwkrHl/mNzsEMHx0ESHvDhikCP3gst/NDKF+22K4Z4rRgkSQZDpSWJ0RwBrHh7v+iOZ0zYx3e0
1UdBBzYx/4uXQ073EBwREeBa5uRr7cTb27SGsGHKTo+AuSxwi/EFw+fuKelp1SkG4FiP4DbpP712
+XUMuHf9tmqjpjVcHfnQLeQ/tSYfPIPXU1i7yxqDZYmhoUoO/ALlGo9ul2CMa2PFiQYewOTz1bQ7
u86+m/BVxJbUzbWw8HLP52yax08PRcx2vwH2IoG/hAZ+aR3ue/eOlPvN7a7oU87QJW/xr/E1VOmd
iJbs/7inHCghSFf4BzbGCe2/ZNgXvofbjB+wHdqNr1YlPA3PBD6D+YcaKwHCt0xBluXs116RbpY/
1N9TSivyWydc8/IkdiHtI5QpZxHxhrSGP93wYhbHxxFyKGWX0tv1tbHgguWuyNb/1SDe3MzF1htu
GqwaxpC++6D+n5ic3+P3DxiKK30mw4GSpVUUZYde+wyYdloCBJwHrm57seHPPQTvews1jLlmjkqv
xNGNhQeTwsLPOjc1vnPotfb1W6dgRVrWjr1+xEx3S1heLMXI+OQXwdBOu5KCnQ0kJKTvnJUnfq0y
bB6dIVfBHXaOomq3/DIX45N6MeX3dxqPmkFVdeEB0Ib+4FcW6EID0tKT5VTjTkOgjzqDM87y+kKt
jj8qZgM3fuZYXBUfG6ZBOWqhNq4thMEv5+2Jw5MVoR6PDOwaaoHGgBVTxNFrEYCqpJKGcytI7l4F
5m7axE5mMQK78VO9n42pNRQ3hzH8Qz6ijGkw4sNVvzYheacEnFd74C2aYELbN+2mK2hjFdloB3pH
Jg9j9zeV9dxosAs+DLHOhaZ6iNFchiQneW+L7cwCyCtA1e1ynTyovLdFov0lzHns+xhCzITYo9LL
Zk10s0fjhhZTETzhNhxd0hcl1O7TbebY2CGKA5CB5rk5ycd97GmzQutFMlLgiZh1NkCzbY0pCGYB
5n86K+S4prls57soL8DtucmXODm+UyMkjyDWJomJyqbi4By1gmB/eme/p5asvnbeNiq7rl/hV9Iu
9HjwlCypv2vMQk2aVoJi/L52nk/qtdvHz8sraxqJtPpMhMZBGuh2v+1Du4ZZfIUrYggPc5yBpk0J
UhK5Gfx1H1fA1rDRBsyVlfXcY9aZj8V3H/AoKv/8zpIEzmSIQStaJOfND8U0OYjjY4C5Bu417LAw
ZQWTe8Klz2sSnHrzNIZ6kb4RfbGJtTt3qwWNQo2M5/nDEO7cSkj1d7MzlznDaR0qNPZtvqpsE2Ng
VhD5LCUo1mBSsgy/HrKVa7hnxyi0x0jLjorHmU3gvhMFIQyHpjXfNBmNQ5dgCmhB69G41105xw07
V9CQpOE+fbkwG2vSVxBkbiwgPM+bqW9HrcbLWwGyZTvE0w1WVfmGiroAuprerstJW/GOUcmaZ5SF
8mc0b/CUSKwy3ict7Nkb+Wggfti9SDIhVof1no4924IjGni9gWPbG6isTJxnpxam5glpOBmfa/XW
8Vv7BUpEiDdx3X1gMNMCmNt8VowCOydZeoY893ugTHcYTMo3nr+6AIHo13YZ6f4TzgE/Nuq5dXxe
zTeBwsjZtEmI6DDAaQmE7VIvy25E02QpC6VDcgriKeCN230Y3iq5Nfdx8SHIgSuUEG8MytnQ61YC
6/oTpZM4OgOmphvqBoWwg6kYs54glrqX1pubx0aSiIfnWo1Mx1JCQbdVr2ggeGq6nex47m2pE1un
jGff3Oj5QN6T9GQgvub/Alm2Fb9KsjD1Ktwyu0QLBQmTnMGPtbE6nutfI9+Gr6hqOkRdw+aLtOhV
28aHHZf8Em6GWdjfsBU3+i9XZ7H9VBHysGaN1JpAeZJzBGTixwC7r8x4R2nI+J7/gK4hQUaKfDox
/rC3BpDjZ40mcsRuXf5/XmD9bFswi11/XGxf//BZReLq29jY1UAQ4g1ETATfS5eSXf4j2CmdlHyJ
zfihXUylrkULbSvkF0/jQ7glZ8gpbEKOl2qhpfOYkZ44/76Cd5dgMQKlbQcIEIFxTdwFkN9WMWyJ
fI228RnVCoSx5BnKqB6tfxYKmym6YyvKgi2R+oH8nViPRPLPE+g9+X2h8OWVjci+vTeLXt1kvp/H
vVogmxowbtm8yrjTbYx2TsyJt4G7ZQG7qF7vhngIalx9HJmHLsSI96AVPnX6tWCP3Ap5xKLJjMol
Y+8sgYVyfLWtoJxAvOlnhiQqO2xZ6KC9stuXeYMhUnLwuAo6XsgCevFzMp9zTsy2tqV290hnOKma
LiA29c8Z51c6smWzNQJMclWpjyhSixNXo3tzN8zcuHgZNvpjiFbjcNaa0lXCRm9gNVbgiZT9HKd6
LDh5IFjE9cxANvIjvpVItkREjVYQhMqU0xCvs09SkokfRuTSU48f0B8qHvIsiuaYwaJ3JlA6jaJq
vpOI80UI8ZfQdu3MrQbKBXlLR1GBkvM23mZWB3/JzqGDM2IGhcZyeDJ+bhjIOqTx4p5Q8RyQcZH4
dr6tSSSDDIMAKqkR5OKalk8iU8D5cK/OePm0yGOmwS6e3Oyo2uFuOkz59BHDlYWFXrf/w8c5IFhT
DKpLIa2i6IkTkyMqKOoNV8ry4Dpi/z5uYQkiRYsCwlv/edM8oDtfq9AtU5x45NzxehJ88BYti13Q
E9EcomMJEKs6JSJzjXKyzGCiPqFBUtH9wlBVJ37LTsEj+sg8puu6mvwEspoMckfTV5KiKiYGncnA
0YhvIQrPks/cTbA5JS/VSkPd5ap/FXp9VVFctDebTaHT5f+Sr9FZgr5Eypi99z74kejrnWw6m8pJ
XXjfifIWaheQz7+/fMse/oGALS5rWi9CB+yhPZ0kpNiQbp0THWNciQ07nvqSJE0cYDfhryn07xaD
/hIIjCn55JMU8iqjaVSDFZzFBOM8wxu2PqUum/tZ/w9F6dIDH1pV7gACXb/XcFs/s54sRgkCJcyX
klYDSjYiAFW6ZMkzwXfwQRfPPzdK5F9gjI+RXbAmgdj0gIultcBOEfFIw3dSsMlrzcYI81isM5rz
OZhyC4AxlMHg2ChecBD1yJooi2FNc5tTBwi1BWeJ2VY7O8Ve328kBVPIvBDZ1KbhW5G2kuhlOtIQ
Fmf+nbLNUGRQpr1UPIjkK0qGkzp/T4jotkwijiGY7VU1VdxIf9nT96haB7oKdATZ/DcFz9eC0Vku
K9/exnopir1K6jem4mqziOj/7dFPlrTP9cAEc/MPb9EuY+yMyvOt0o23yhMEp1LhPoDxGTCjsr2T
HE7SQzWoDMZJ7ZJP5jQhpocN69OwT8atzEJkq6pBM49Wc+VFN/+LIr3/K7LVGb2l1+mOdeoXMnXs
vA0uPnImfRuyksU04GIIpr+ITmNeRZL9b40fqJuoD6K65HvhtuiRLuu8YODEmXAMykNBVV34acRR
OFw5/yMzxh7UvEu9Ii8wJVEcIN4FHbCGSHYJt+pIqlDW0/QO2NfDsGQ8cxw+KfRDjgzPiKi49o0A
0t3tHTe5V1Z7x7GVbmkFPkUn2N8JagIV6drAccaUzeUxcgr1uzmzdLliN7vhHBZqrxsAE723Eduz
zGushEuV5i2vmcyCLZN0xFD57tERrtbS4fuQ1b7GlfdoeusUL0utU9SglsOWf+vklUi2ugSVaD8J
T9n3151wHnXPDHk8H4YULGr68sPi/0asJiKGKxElZIPm8sgt6aPNR+sjXhzljqqMtN6USrW2KRUK
j/BKATh7AX/z1UbAT9voVnjVauPDyMuQL7tPLBtL/DBPbbw/np9/6b3fbJdgA4dKSWBLhh6ziq0K
xo/8eq3RqXgCXfBjGLMYKIDF7hhv6YV+0b/aTZ8/9ro9PFGj3T7Tm/qgxkg4NVoJt1R97Wywfx9O
2tEiGpogQWKajL8o10mC9G0YNgSUyx2ElqGHffQ3QXNSrE/62Ma47QbYCnnJVo+5VbNy1dmLBnHm
botFL7BFfznwqkQ5iWsmPHn1PSvv3KMnDKFoukSbQLoKgwJSkUEGza/M1xCARjQPnYOUwae8EFRH
AKdAxp6GGrqE8+LuzfeodyN2yexGFlmAtRrqQcudVQ3cKfvyxk72xd7Zt9Wgecz91aIUUBHWLfle
OGslSGJ3KFLQjyIHltqlwnCiKgWbfVFXq2zov215ZieTUVeRzKHRmYA+4ZShclJxsgMVHTjxfug+
dzu23d23i6qudacW2WoY/rsc+OA5ca/imP4RuPhHBSF0mJUeszxeDBxuLG+Dkq+A3P0lIBFYqBNM
9kE9ZcmHPRtt6XOJtaMsVevUi757TnMUbNK+kRB+yyTAwcI5+w0SZNYtS2OMBdnypye47xSZeZwa
GcD+PXV5JE9CV41xNPV0dqRZPzTImVp5HfdRmFeYNgLMjOx+uRolKw4T8JRTxFD6ygzvLJ//+Nd7
q0g/Igj+u0Excs5/SxZVq9tNn4cCZcEvpa0slQYI7u2YSmrczMX9/5PtHHqBMxN5Gn4CSqt2hBxA
JcNEYzIsKivOKhzVYNHbxkhN0jgJkucRYdFy2RenzpRAcqGyNUCx50hsUQDjvitmzFKgsf1yRiNa
DgKD9WX6bOLb+yiw+UNZYSKFsCT71GpxT0/QWGDE2f873Afh0pYcsIaJsFMy7CFafNJdMKIpTcnc
+ifRGXIPa5rQHogB0AuKkh0IKmnIJbJVS9126CK7auNjjo6S06HlinM04TTBwnWi6vubOiKOCinq
B8iUzuQAVSZHhCFaWIeOe61SxALJhskAEIhOatwd4PDL7rWolrDPmMYT5v4YDd9UJTnhGkMy+HN1
4Kt/Br0bPgC/0qg632ixSze/+JSY40WrK+bMx74LD/jOkU5pmtwZ4nCAj54okPkgxO6bmxX/4svF
xbNc6U2hcSgCCFz9fGpOi0JAebPYm0FlP3nxVQJXIct65kqEkGfzjfqjdX33n504ZeJ49K3vfABr
EYegBBySdbxT3tOA6brRtdsAbgDJnmLIzof8ZuUjG4sYXMOgHZWNsiCrEEjDbXg+5eqYiMNmCLeL
IQ458St+xbDo1u+8CUtpdtITG8zRrISv1slFIWEWEbrQ+uMsvTLFeMxl29b0flbiMWOhhIyTuMtF
o+O1zzGShtLKOR1/YHB6/BlgFvfcsc1xzWbn0O/wC2BYDZ9wRpO/i9nzViHn8wfQEDTpRvXh7P1J
f5jn8ykTsP1NTTLvyy+ATWBMwVJS+0sHixTgvsqM2JhdFi6+bkkjjUCPH1EwQg8KDRfVGo54ACPH
AlYvcXlPBf+W8swoi9Op4wUzdxCZKj6w8PFpxUBntaCweMOTKWNFpedv3sE1bRk0gUR3hTeSkKai
Op1CPNaj9hjO0zZMRJha1t7oF0As20wpb46S+lsnL88XvKNvLYi9AdEiPecXkv4y8pIhOGSU4DWZ
v/T2/tSDGIIx+puVoagQjHhV82LP3HUHv7pW699jJjFHEbaeBZ9FL8y1ju2vHgrYNTnswON7rQnZ
Zwsvo0pBHiG1Pdp5B3fvSEQmlc6hym7Umu3e514hbsPZZDpxEJPQ1hT1YTbBic+//VS/0bEQEK7J
ijO06HsXApsSCXDudJQ3Svwvdfi9ILpkaL0B22C/lPzTlF1A7/nl8s+fs3jJfps4xJfXOhsr/rAh
oBmFr4Esneuf4PBLFQYo9mXzh4Uvy0PjFXQgawuVm/L7eoacxIN1vkdPoXJJ7LswV4qsPlYU6x7i
StKFHLGzaDsWeJHTSbCC7lD/CcfWdcvu/sJ1uZ0YtkvyF/JKKFHy+Bsy9+iR4CBvftsDr/xdthV5
yAK6y5pIuVJsiOPsVjDI2VstHKLnxu+/zGByk+EfHh0kMT6Gh535OVi2VZzykrhG/XsdcoXN98AP
sBaz0rmIM24TYVrTZuqum1BK2WsrWFoA2out/oyRg484ypSLBRceQkB8yoasVjca0kN5yoBwiSTX
z3L5TCKaOyil/sZxemw1Dfr0nLN4m1Qer/u2LvAVV3a44gKqS6/5P8TxLm9z62JDyqkesiOrCjsS
0E4ojzKJAhO+fzAlN0/S76Fb3u7oxteb8jMhkS/Dscs1iYvvvNmeklRikhHkkuK/HWLz1IQg3Nq+
t1sdkwLHihA4aQNFAvNQjVUOd/QRyE19fSdmt+x+pk0Ovy9526X116Gtg1jRelp8zCmJX170Jod5
0UVXFuMromy9eZJYNZPiM2PysiMRZ01gCvf/kxrtkKhROxk1++u2Vc7e+0k3fKmoPwEVbm6kpF//
8Nla2rSKL4EBW4u0hevZ6MexXxqeuy35ByimBUUw1RSStZs6eoo7TbaAVQxDUEQ3hgktlv4Tnj4A
RQqI8E5bWb9tGpFQzuoLY/TR5q3tV2FJcqAAH80bJ9wAhD80RPDf+UHPVMimFuetabztopicFDK9
N+b8Ir0PDfn14kdO1icZ142q8reu6BO7C/7zr7UFCi9abRGjJGSBQDIIE2rKdJikwr8ICVJ5cKPI
4wHOL/pBRWJrBM/eYRRHz2ClzfUY913tk6nJ8ToSf6Ct0DwajE26Z90qmBMSzQrEgojmFz7oVdOa
gE00uAr3PTKaUVYxcqWe+wxhZzRgz6o23jQa4U3IcpoaKN9osJmLWgP3rVWjAaOQim370J8Hqm1v
58FVvRF6/V2rw1Wj/RXu89n5thmVfEq1jZHK7SgUKJ1IXXyzcXQexptE06LIckN2ar7wdctBDjY5
9PCz45l4Ec3MoBC6gc9jQF/2beoL/C1xucOAWGzLqEmtma+wrjKtqE4SpfcrSGYtsxuK3MTozB+M
yFVkKt6TpAHORXZrrughHJ2A7vxI4avkikNoVSoZHKjgjjH12Q5ULCkytr9D0IZKz1R6HrTSv6Bq
z4eT1XvQ827mErkDAT/ck4FuGUzit5YurCbANtKRCMit5ODQvqaN2Bu/nXbIwZaslni/x6HhZECd
eqss6zOi6B81ZLcMUe5FvlVggDaRg3YuI0QgA6XErHz5+ZKxvs/QzKwKmlmCTohTuRjbgyguHnPK
XEeOlFuDo1r4LoftdkxslIgRTWGbDFHR4kRONGTprpl/Iv/ii+EGCiM5DvLn76QASPtANLm7A3ND
G5z5W+tSLvhGa1OD3O33ngl4Bf+dac+ChaMX9RjO1pmaFUsCKHytYeG+MkNq/vvL3RbbfGyzUqGz
dqkHLlwMESrSxulV6oE1Nu24+4BbKDWVV4YrAD84qHjeHkOxCrgjQ6Dtm06xJlDZlOO4n2AKaRS3
v1krdG716XMhAuIcgseqhltln0/RtncN9NKl/UXTTYw6hQwHdGyL/XvILy/CYy9nnUvUfp/b3i7h
Fx4kCjDASeBH8+zknXmeqA85L3hagRzrw6i+7jFEnQZTnppDDH29yzRql9OUmkO/LP9WjEe3FZ2p
AVsWAvPwvjmkZev3BUzXd1umLWMYbqOwfk5hZIZqDLVdKY3se5kHWOq7NASt7hkrATDtlvV/CdZb
mWS6NPqkHTkxK4SlPhiTEZtfnXr5nXt2ULscnobyuYgYJeG9+L1u0/iCFlatHvCOs19Lv6ByWrhi
E42nrOybdzF7CA5eNtzhMM3hkfH19gyClTaZQPwVK8wWtUOnGqb7OKQgk/v1b071d+JDnVGezJKP
NPSFiNJRkVwinirkkzHhL37wuNcjK1IHSDbQIQfknpJE/Eia3UTGcNgc0qP3dhfabuU5gF3SZJxM
4tIwriXabcHPxuK8k50E/LBOs0okpK4BHx8ha5OnE6A/wfSwmmPNKQS8gzEJ72ZXE1agoo1M7ZLx
srzo7XJ1CkBFCrzid1V5IZ5QHBE1MzXd1RbX0mYiEexxQCK6HHW/GhYWjVsrYltEPlFGvUNhTF0r
nJrFnA7BO8+cPhuSvkims0vvTRc8S+vY0Wg64LU6gb9iJ9BxegbmwR8bFjYLpikqzPQ9z36BY1/y
hNgPQC4tsZQVulGauURh4ZP9dPKhZnmc7R9qgL6Hj+cE9fA3Slw1Aw5xL/72ytUeUwqyV6L+VXH1
m7Aln+Tw7t+UT8SY25eef/rNMdZT2FfTIxC4LUn8/suGoXUxyFB/UT8jnY2JEI45JT1ZA8jiBBA0
b2C2MWbYMKQGMUdKv4LBtxDpsHmwtQFbN7D3ZXlezh5JT8F3LLCsYsHlZuGtkHBmwyoQChYdIdEp
ZLSULHSVe+XEJOM53XuF7oLM6MxhTHJClCkfVF18gRYCJXMsyHJKE3C5nVCkCkfTCA3FewoDgqm7
uCTLerWCs0O6Pola6EtSf9oB/tB/YqCWICR8wANGT7Fy98agmVHHssZqJ5cDMACmV+1EIdvs25F2
GHprgZn+rlp+HYSiPtVqKTYCi1NCCyYcinZPSx3owdDaOm+KgaRC45wc0UigtUIOm7OGZWvNWvdJ
B8/aI7tOEFALTMu6npLvAamUlIOrceOiqXzVxs05aMmVSvZdnitTqutv81cuCilbqOndrToVA//3
9S17tFeQ7puz7Tsi7uVHjzFxh3C524Jezun8K4r8v8jiEciExk98Es+F8jIXiHLx4TnL8Ga1i+L9
/BGk+P8rQ2rJri0Jgme3RxTcQ6ByVnEa7IhoiF0KEqdOkxqsUZjLrENlb1qKB4PrZ47ZIZtHIs/o
GUcGRHwKzJE7PqUMaqkKvOp3/iPYee1P61Yd3MFx4oGxgnUAEQurjOs4h2WUsrpsqU9dQLXtjPZY
IWntjkNRQpIIxoUMrAQiDmFlp5rcthRps6/EaOnrmH8cWhoJSJGpSq1r87mpBWVsWqikcvDj3OS5
6ro+IXAe7PacGYvlr8vEfWrlcyszsCUpxI4SIAr9HVWKn2RJzl0kW3iPxJ4Ij4QFvc5g+pFIu9SH
17yI/hl5hI2RR+tj51iMygKrUKbaPEWrOQQlqrUt/wIZoR+XSdLRhav9mW09hNITt/y/tqEDsAYm
Zur2nGkYADR/aWPSV2xjtOymGwqCns+NImI3bzcjjFqaEoMuRbopqw1XJXvrnQmKCHyD2utpJot9
pFNFHHNtzAKk4QVlxFz6nEh7cAC0oWXjD7yiqCJCVlePUQTiq+g68+SxGqPqUmlFfqhfSyIL4pgE
+0yzzLH05ScnpEN2a9Zl4//mExrEHwJsdEYUStxYAnmJHQRcnDjgx3dVKlje6F/7/hT6UV/xtasQ
LtsAEFwOkzXjGpKCm6s5Pl03hV0v/WhtQjBr55m6LhqU0hi/ohAR6XyRCopYYP2vo1xCj0ldl/hO
y3MV/NpNNgu4mkzrFBF6unPc4Jnevyw97QjDkfZFBiWfJeoNhhthuC3zzfb4DvT48H8qsANJLWB1
Mc3f5h5oEF+W/PHb7usIsjqwu8ldEYGlGb0naDW3hyzwZqhQ6nskEMNj8BIgGw25558vcNkHTuFb
0utrK+c9zb6tWuRBuyuGuNWS1gg36KgGDL/VHHk5qU6zvkT8/sR0VdL27MwHcBa9BGtDIAR48dX6
6nczDpRdZMpdLUa/WY7trNnRGhbHTVlPDg7rtf8mXSv7NObw360fd3rQJyzAiTl2WGCSE4MAsxt4
7UVVgLnnbhnqZiSO1lz6evoHSHdVR/8e0I4ENqqAPwVIQW8JTcf0uz02UNDcn6MeIJwuHTh/GXKQ
C+GZ8pdvXunduXKntaDBOGI1emLFgcKOOq+pQdO3Yslu66shhOZ22RL5XytysAnGuE3ZGnDMpiYX
JuGIdLIqzoON/GhvRtOFMftI9xRE3pCGfO3qHBHZbLB4PT3b4SBmEjAPnDzp5Jfa8v7xVCTFRzQz
B2TIvuwoS8clJ1QKzzlUgLEq2HdDNASZlYs94uK7igS69LMkctFgtW0tce8ARZgF3X35R0QmJk/u
ivQdIkEeWBRpFJqkza0Oh7mr8cRwBE+c+gJaOyBtR5dXQ/+QE5sjQeGvZAPyAXbM+Cvs9HxkKO7C
sXyWHRKCdVmDnp0ETpODyLGlwsqEW1zNTbWJm0OvZ/E96Cnagvgr/4b8UQaT5LZf2df+TbMz051r
5pLmW6VVfWBm9SNDmWeGfTlqAVRtFijxl7s1Pme9zDJUx92JplBYvwFIhQWBcjbCPeL4pPhnNxwY
KonQ2b8xL4oz5ChUE8UqP/fD0sDb5TJoJVCiJ3Ync5NPQrRUr2Ss8WVTzQyxTDjkB46T9PQEOZj4
szewoQhncOCpzSzWnGPNe1fgB3qmjuSdxgLv5vBVFUTrB0U9DeTvqJR45WmUeCuSroCr6vgKAq9I
d3KYTQAdFgaSFv9Pf00zeT1fvUUutdW0Z853puyd9U1YCfK8a2QhC3NimWyKsuzzVUnWbf/1CuqU
5rYAUaLvq9fxBtzMeBpNnW2skcM9W2zlLJ/ecJQq0/0teJMff7SIRvXV/Uz3bBknQdwDckeFd4Yy
esRywivCG8j9fvpZKsXgfbpXk52s/WL9AqS9TIucjUun7tAxKleh3T63BCjLcxgLQrZ4exM28r7Q
8Gf3jBvS3HuWrOeW9ltdUBjSf2CMuPfvEJYEzG6IdSwCpr77pkzlRiTIPrV/U3zcfplTVhtDJUYg
AEZqgjeuUbMPLkf6SUHrQ4jotFzlOf7X0MDu5nrfVuDevNbJAxfL7bftjgjTQ4gSYJFBLT/AMhl9
k5IkKI35eRMpmMie9uKXRuASjtSXBIO86FqbJ3E9HExjg2JUDWFUa/XgFaTGnfAB/OcocMbfB91J
NotRPruBCkeR416VKD+MxHVgpJATlyABpOEsx5ATFAUYRa7STBsXS5zYQ8PpfzvWmEcsvb3RMYYP
fWiVb8xIB76VxXLmIqwsvQQeBQF7TcgFatrix5bABlr7j8qBbqNhk5HxFxKWMZab9nNzHTYuAD8w
jvtzJxNsPD8XBBabLZ1otVj/3oqT62uXsU6v9vGMf3yX6mPq2Dia+BxQ/nng17URQr0SvjlQcQ+o
6kbhxUClurlGxWSE8C0CzFBiQtjj7jpTjj8j0GlTgB0JHxn9MVyh3th1JglGOh1PFvy+7gFYKKiR
c62cUGV3iM4nJ7r+bxwNDbnG4kZcKuu+l9P4nmeDeIYLejb0nF3mQ5lOzPtK5e7+6PHveVuonC9B
5UYj+0kUJvEU5OFdPEpygPnd9zleof3qbDG1l+jwWC37KL9FKocN8jm100gKEnFL2sYtAWHjWXkU
G01+HrOES5F4yH/Xue/6u0ubrMJfURxV3jBCAEwtzfHA1ZqRkppE1MbqYcDq6NayNP6JwRFniKhU
PV7+Fe5DOFssrPbjIXonXVQhbx8kucF/1BV7WhEaJ7Jx/dbzsjOtK/PJpo7UsTp6gpjVH83f7cc2
J/bfp1AFpVQoL4ZkkVjGL7iiDZnm+dBBWOxZysAVvHjAA9vlyRH5xYjEjF4djaovYmEwX/xOkljr
E16ob3fTLwP/U9pJUMSLQm+dyOCxCfQkgO7P9TrGJrrpZ9CHK23Doyf5zKvQ24rm//xL9H9HFL4v
aCmZ3dGdqpUydTsQ/dPEMNp1Mn71BDGfvnpopDAi5S8NhWM9tWUtBUNaND8rEk9oh7JGa7L11wxP
BimwHsoqOQS8TfZ2np0iERr0UPk9tYJ9PdASo6Bj6CZLH/uofp4XWb5DlDtUbGom8p3uMF4VGBKU
wT42QCU0KugU28UJJilmhPhLqpQVYfVIEnbSIvLScJ/miOPI1bisbaghfeyrIkQCQUsxEal4bvBl
jLyEUvhhs4q0PXj1PwMb9Xa+Xsw4tdBw6LUW0ze0KScJYRD0SyWMskPhgyezqefKfKoRRYLzOEsp
X71mueDHLsKQhJV+WAl1840saS6wm1GdO/O+pw4qJdptKeVIWzcn/NImzhwKm6BSVK36ADaIcTEq
IrdIuGguoCvtt1aN8f0bqfcXnFwXS5PU65rllfamjPXhUFjSO6jtfBJhoPCXESc9X4kLqhZ+zBFD
dWef6t+6nzTmkh1zIJNUe9ADPIpMEKSy5+S+g7RiUEx0XiP4owl6nQ8OvI9Q34JrH7myLXE6zxqp
SK8A+HAzd1Nuo+a67tMxz+meoVFP2TMGjotMl3OTmnm/Hqaeys+9Mo+xm566f/V5a6eP6ycXExbP
MdtDHb0jITR3jEZBUtjWg1Sr/RAokdEtr8rzxII9DgMzPirxGnoFmrCWTZbPVA0CLBvhqkxt4q7S
X62cFKFW1HiwvgvW/4p2pcltrnAXe5Xio8WJ2fGpBz5mbYU1OKaSEMC7PcHD76nTZfENENy90TRm
xKzhFSB3H+/Sp4DmPePucEQseGr3I91IowBmS6ehX1zLSu5yJHiZ4EVYjPXw/kpb7NBONUtKj6PE
7xUIqQ+ZB0JtueLUlUY7vtSzo4leyUJE8W1Z2qA5mkxwy5p5RiJKNN9KJyS9NIJwlFrZB2fKAOVo
IaWc4mz7KbM9kQrb8YPmj+5pP8Xs5Sl+tdSX17oH5Z/XTnouwY47L6ko2MTH14kuFaiqOiQNecmG
swQD5/bH7ZCSDOz2YTmQur6aQVuN6bP96A+T9ugxy+c1ALHYm29r6fJ7XWDE74U+hV5kE9d/qVEr
3rXuHYuD4bQLtcoOMjpggFhYaw9tNZsY/XOgjMG8r6OTxKF3t0urGnXERhD3Xj/Pm5y+jJ7zyY/t
Ik+7n0xp4iZBLZym3LQOOK0Z1HXJhSVhS6WoUFXAf+tR29mZE2AveuZN1odRKfduqT0AiIodGLHd
Ppy+Arn/eeCBaxqVGoEe6X2DeHvh1W24WW1ZRG4qOfo97wpjxxpNWrW6jQWQGszJ877xiw5odA7H
6obuNfX7p3Feff8Zrse8Bjm+XAub+Q05OSiNJ4EkUvmWSF2as2d3UIigRy92X76r376iDDLOpPip
oLHRlGCxqGd96Xkiy33BKAQFG5H0GmSgJRa+7FHxql7RbqtbMofpkG2nb4H5FyAlifNq7xqiJWvw
52DmH6CE4n1AyGTIolD1zZ5hQmJ8PW4XQ1eOLuxNuSD/YXMklxjYrjiqUXyNl2xc5ULfC7RR5pZp
rbjBhvSp4D1aoHeOtOjDOtaHQzXNvrfRyXO60EoLEdJgiOQIB9DdlUekulz4Hh2rkrNm3WbR0ym7
mhX2cnvZQWOK1FQKV7m5UtxQJP2gMdR1u1CIZ4cMKW59/HC1Jn2T0/ZQKC55gIKZWYYh1k2q/c4v
3DKh5LmxOda5GntVETQcUYyi3aawJ6slf5OvJQDEn8C+PsF002kXXiiVcTrDtWkTAkPu1UNDYzrb
WPpLwE1YGYsSC4yIXLryv7kD+Ui2bKLhdoZUI/QYxfSuoI3GbXnNEuv80m4Cclg5bHXx1DntVhF5
rswETCksqvXvUlMB1crxvZijP/Q/5ytiPxyUWEyu0iOd4ZWNC+Vd7xaVh7XgnmXN7h3f3uH2bvb3
cPyZa5O1rGFrnEax9kwinUcGLV18XWyklzYLIS1V/+MKbsRULRyzSh7OO9s1U1B3pYM9wuT+3ey0
B0ledltTEOs7YJquTDY2HiymhURj/9DyIui/PafVWZMoksBypOegggEls6SPoAYZTWolGnrR9Xcf
da6Utd47ej8A0UAArocsSPrStj/BZEMaBs0sM0UfqWSSYcSgAobIg9bqHLOtNHaqn2hzIK6kZI9F
ek0rgt+2Z19AUTs2XO/KHVzbyKe9xT///HqH3EHNHvshRJd6Uz+TX7w25pO6e2j4j+ao1HxlMDsU
5kIH+iXB9IkyCOVuqFxonC7419JFzu9hpzfE1QzPkavkvETLfuCPJzKzDfaXHBa6VjSawi3DxmaH
4FsM0NjrGSzuOkC26vDwaOHNLNTA0FfXWkA/5T2vzFfa3COTom2Oz5uLoZ2DSQD374X4I+v7kao8
0rPJ6FWwW3dDZms1XNeUFjbRvk27wX/BwYidfmmsY0yLTGs6G/Cq64JKiNOviHtkzYBEkhfdkr5U
iSiK4NMQsp30+2SgjeaKGsP7Eakl/Ac0VheZq3DcTEWcvngkYlF4EckTTJygX6utm4ibAzLKyB8O
kiKtk/p7EPws0krDVrkinyyXO+RlMRNRGf+qaTseKxAn335ujoOktkNgC7StcWEd0b3XLRP0nMKu
O/a1GGQv7vtrWRAFKzeBftjJrCI3F58mSLLgdfYk0EGX0ieZfRZjizFpUGrbREFvcSlagOac35jV
7h80vlylUdV6LXS4lLWCe84R2Y9b3h7eMuTDCC6qC4PWx4jwnPSsS4D0tPA+e3rw7wg4kM2H2bH+
NyYJG6fIJuPwkdNyGQkGhTCMLnUMezQf4mBsKvMzoPUmxdAuH48Ic/108/QsAflvPLoIc41yhf4g
284z6lUmwKtFPsyMDN94v9uQwx2Uf1DgxB1ifYEbF88y/DVbCg0rih98Jh+tZCa9+gvlhoWAXWcC
hkjNeO8JZjpE0nBIgBRMoud3Bu0iRI9/nJgDnoY3vGn0HxT7FHyzjBsqgFn5Qf3tKIE6caGebbZx
GWuDA2zQdpMh7Y+gT1JQCqp3oR3Zim8kD8xuzk48oy16AF2i7uckXzl20c99/oD/mJNoqpWWpcZU
OA/RdAhaIEGmdZ7HXwsAAWoDOA8cd+Uq83qWjovBQ+A1htVin5OP3nsrUMVTQo/fAYwHF66muGiE
cOCfh4n0EwuZB4Be4K96nWNej8miwqqs1X4M3g3uF8UtVQayJWfs1Eul38HMFIgdsULipsnOJV8X
U4WCTc+XIj6x+6D8PFmYzn2fRPzx4QbPUSV3UqouUdX1bjLTINX7S2iBID3jPysnDZbpEqN2RHNP
ui1ckW7iKBAUVRQUi47HquMi4zCHRlztsXc/LXLc7bOH1oZ4lKBBtDN+1j42aSPAa/pgBkqMqXmF
/fT1DINJv8l2Ud9LJHW3E861CSx65Y4XR2Dvfkf8KHjA5lFD6/mbNARqt3QnwRO2ApOMbKHr7GQa
0hF2DDxq29n70Qm9hGCYJHRTjuFTO7/WOL/g0viGH7WpEqKbfSWvAmSNjlBCHKNN+nozELdtHLRV
e/TxGLbWXgWCm0SRo6JYmlZFXFXAkk9Zvm6er9BStDY5fbXRHOYhPvrdiU4cSw8U2hPCJK3MXrCg
EEkP8MzrTqvL/UqJWKQpS0maowqkKDbDJo+8KjON6EOPhdfaz9QlX0A7UKoX2o4831ZDFYuZ7R0h
efiTRIb2+4CnctcyQTPHnxEtvNyKgDq4YXRKr2hVQkVCWwCppSqdpi+0XEtzq5r7XTEzyuBlappp
u+GVjcT864nUwbwbp5dS/zaAiARanb5vtgvZJyDzWR6MonN9gDQ3j8rfIVcyzEKUIvrTqgw1oqng
SREctaNMAa6P/lpq1NTIibTfbO1PrTlRf6WyiMyvtNfmXSUUt5tWBSVQrJ6n3KRtHQeDQRd9La/z
5PCTh7s7OEajt9GXCFzv94EKfYoS56ul8hP07kzC/CQetPXOpmC/Kvm/vyklitC7yhN6Dh54RtaF
92X7mxnooEHi121Rs6L7xYVBEc4SQjmyiNCaG5mwWB2m94RJhU6x3LQ1Wiyfu1COK8tF6PnjX/zv
WWIa3x6c4IVuGT3+wwtmbH9IcHQln1VInppvrcV67q8Kj3dTV0y61IIDGfu1v+T+Qcegv6KZfUGE
glzhvckDZ/Q/fIzGqBCjiN63P0wM/rPJ7e+eGlIaLKEg4t46ZYiV0b05P1lJUi7DI+gocP31ab2p
/DNk8LkDBIpIw+CBlfwuZ2rxv5bOPc3fC/gU/c7gTGdr8grA+TleR1TvVI28Gp9Ciolt+MZQDGkN
rOg5y0q3OTSaR3WCTRhzVw26rRwp9ZTC4ZXJfDVuqAWtMMTelo/nPKjipSO1YN/7iyxIAlOCADrs
JQ8AqMRCmIjqlwOcrYALfKoL5cfc1zfoDYeWVJaz+Au314W9G3SFxhNjG3Alhj6uTrqzUFNcgn4E
8iNWp3OjNCF+W41pgTyPQMcm/ClxX3QG5X0IdJKTEcwlzASq4DSq5UDSUYcynKwa4N3d3OnLQwQ/
WlpkFELlWr2fqAg7302m6UzCoaUqmi+6gErj2w3bjebX6mfsIMBEkW00qdGeqMGr8Ssx3l0xgQfM
Mij5fpErrmLag+jYxy5k4jEim1WHpMv817nx3cvFkMHFZnQqIHAcFVeO2R/QdmruovAacHt1XniZ
N+QhzHKfDkfEQHX/ag0/6Ys4j1EYlXK6pYLsoS2/v60+PEoj89Bx/P7BaFMVnbfWfsxgCcp2SlZL
oMyywttFmc6ksghvWU8yCUxDIZIoDpK4R2valrY7uU7xyH+MG4SKtbPcYsPX1ySTn1LSWY7QqbNZ
QXOCZMhxGEZsOVVO7S5lW8TEYNqwuDVYs0EcwXOJnNs+97DJZz54Akihz911VatPZ6LjQ6yRNpUe
ycwd2kkLcOMLwtjdg4tmIZSCjH6EauGUpd0/CcyG1rjj3XE0SossdqnYvvu5vpt3VrWCzG99E0HM
aVtW/YK+QmqHWMzlnEEAlkOhhi1RVhyqizdIL2RhbO5njY4VRI9U1UdS5W6snwZRe+Ev3G5H6xan
DTjtTYw92V1L5gvY0cGCsCjdGLrwTojFaIpe4wBSpRj3f0X9I256i5mliCTCYPPB6dZXRHHOs+jD
mgSKqOl7pZBMd6HloQAglzd1sG/WbjOeVX2/ZhK4fLwJrZQesHC5NJyQStuZhsO8oOw9VIftNIzq
k9l1FYG35Ct0LEzTARsVa9CLI44svOKsko/khOdtobKhFV51KYFiogSY86HLY/FXW2gQ12KDaUPd
se6dQAJOGyDT8oOyuABpaSxlbN80I99VgEjA2irMHTK/xXa3+opcqLxvDj/4z9Fu3xEWITU0uxpP
cV5e2aeAvSdR/WMtOQ1T66C6+2QwfJcwkJS0ju6ok+6TrepeNvddsW6hFmGlQoCfDWMVWfF3jzdv
tRhOqEaQXUVT9xkSkGzsaJNr0kl9TZnifbiwX8lkRivGm0F6ZwiikNkeox3Ffmbf36t7KmXs5gJk
kAfy6qxnrcu+mFqtgwP+9q0iGANO/Ly1c1zPCCWjXs1bOkBI7ZCwh6oT36+qmz7fxRG2UkVz8lk9
8fB3QbpkY8Wawpz08hya84sTNqhtafL3vFxTqYkkhrEfPDzq9UQGCy6+1VAmTvpgGHOT++j+CvJ3
SOT0YxYGPAfmvTFaKtrSreZJP+RMb0EQxNpLSga+Xv7xq3+fTFeBLjDMiWVr0+8Jw9uu4S+lomkE
Ao4T20IIJXNQEinUF5is0UdgFp1Gca3kzInkZyceem3Hb0W1qOvDL/+RPcMy+b0AghF3VmfFkZpj
x7f68ngIgLCdpSFiJPaxBjHlZ55zQK5gyguv12ZzfTUGO1g+wJrEwJlM2JJhTz9zGMfBGtjk20+m
Eu2A0ojWEaoSP5346yTx1C6HtxYzBlWZFyQAdrKDxqt+k8scctX7KTw4qomntMMK5Cn7MzN+t66h
38wRy9WNWL3vPXWyN0g2P60rErAf23//Txe9KN8gW9HHKH/QSky1GoOLSP0ulnRKFfbtvE5tLZ4Y
7mqxvRWN/1I7yChUy3qlSfv5Q/rKTMVsRs8zUfdCVgkmMikdovEa2CiGVBJHdHabYQH0SK1YCHzA
P28iXL3aHpSOjpjKa852TmmFx4Anrkwu/0YeV+24dE/VpQ8pHpsexF7u5030gzZVevCdvu0QXvK8
mtzj6NiqhxasfkoljHGFfAzMxmIgVF3JgZK7GZNpfUJzPLUessVfFHXuMBtk8cAf4X9r+Or7XM43
6ysPVaV3Qu0R/9rnNk6V8JC4fD+2zXcKbF9MS86T6yj6+DHuEAGfnVeR3E1Hbn5ZEwiXJhGr1uNv
sDc+nPLk8yAyYb3BJ0Zlr6XSXVdvlJ0+n63ys4F6BGFAZ6BFw9R/5KPwlTuwJCH5lRQovcSgc3NK
9FDynRpQYvnVuE8AypXQEADSXAUeJq+om9+/bMMU30IU2llOaTVAVK6wAKvLVAiV2cXwqUgRsXhC
dU04GoTr0aW1j61zlih9of/OdOGZSV3B0CC+yuDmnyysX4wN/HzOwcsm45Af8blIM1TEhTBHDS55
/Dd92xxKiO5jMGtvXMITWOMZzpTfvWSpMlqWLq8Foiu+X0Jm+36tBcs5fhifzGzQWFyq6aqd1vf8
/TBWWcMET5qIItpwHtgy51IykmpRZ3DBYhKWlQCGUEdyS6RdshdzPekx36ZqoV+dmjzRNMJ9YhKv
KJZ50PKKMKbk8RtnHgnRNvKbMjvdviqJReu89yklb7gAotufuFVN58AgcHh6rvvBGiOehRPuCMCT
8pP8umKaUhpUdQsil/7kCLNMM+UiFjeGHtks39lCB1QLvX3aAhHA6Nj5gaIt78Dr5NZHWVlS4nRh
Sg+cZhDG/Fw2/cliRjuM144UkIjXvNf2kJB+P84QO9Y6NJM0LHje7Tg5N4e0mOf1jnD6kW4/Ep8v
aIIvYViS8ZyOw3aG9/NbA5i7GuayOXELd1E2YaCcY+AhwOsBGcdNL7UZ1tJogVc/F5nHNHTTc1d0
S4GdakYKaQBbZi2jsUrCed63IobOTVTDAwVp4nfSx8TuKBuqFkFjzuWGmJQvTREtzMGQRBnD47CS
WnISbwSh/qfOb/OXNx+pUnUn6TjVmkD8+qIlE4pPmjFi3bYlN8iHAqVijhSYYqnaxAVRnC/SpOrY
FV9sGjbXzWrjXTHNHm3JolE225vLkW2eRazWATksLZs9JUe/s3DSsbANwikYzuwAor4dnOCpfDyS
GqVLTPyEO55TwJTRTplPfOWKbZ++0Htdfuz7nK9Ubk6+VQ1KAV/UqD30551rpu9WGHPdKhQFjB2n
mrcie1RKTrbb0wTr3LiNL0IWY+taqJmHOfl5hjm3p/jdWyhvCpUfZZuXIGrs2vwhtPAKZwOgp/xA
kkuk7YOEJaUQ62a7oCTeghfL4wvgF+CE0lxmoBEXsc562q8wHY9eaDklRDEV0f2WN9MWwmLu/d5q
rkGiQGGqkqXI6iCMIHJPENg4x5QjyL8WbSrpBxE5kiZSm3ibi71wWSDC3zwiClQHbMqp6DJU/0lt
e9sjRwoEQNvqzPX28hKtnaA/mfKnKspUSVX2rNbromL0gXulgJikbrOUIOdifWSns5du0XHiE+6a
KJyAru8wm+JQyTLSt5RKPFEPl80ML5+F5OM3LS/MrGu+oW30FOPFrW46aji66HeK5X4yBVPK5gso
PLY1QXgEiwF/WO+9pdv4f78mmx7yVuQRwoYs+fhhnK5pcoFfB+B0uyiFMqK7XYYYjK/aTkZBeH8Q
N19oh/QeCXITCf88v4WcZUGDlnCVqu1dWXY9oBc5Q5j1+NN9keamOkb7GwnclH6jFfPgY/ezzXxs
R9OADhWePi/Rcv8v6S7OJuj6hvqU4Tem+kqW3IaiyFrsirTQMtDoKV6wq6b1LOnD5zavCy0AuINy
W0H2IXbVDkWEAWUHZkRvjQOpzGHZ1JftEskgNBXftIt9TnFYPfiuqn9x7jPsv5Yoj+NZQx52s05V
DdDT5oAtSz6duFP0esAT6g0lefWi1vL/kV9vDPtE8HA6wYdtOGrE52VcBM52S7+KW/g70iRpJER7
EvdaXxKCjje7C+y9sjUbVMl+Jk7jrWY3KNQGMEh9OZElt5poKcLv2G5OZxOj2H+p6jlqBXFogH9V
HJaoz3smAapbLiZUUKp2Sf/9ljTFfRK9wLTlSYaKcN/l5iKQ3EZ99tisxkaOhZnA3Y4SUvhLTMCZ
dYu8VdQdEMUt8GwxlFnY0xp/4r/yNRf9TXbXjCOtG1PsaXZIOoWbtygL72vowN0Z36DYwwTjtk0/
xsxuEv4hdzVyw6vBESuKcUWi2hSzFKVkLsAMj+T0OD93zFfTL4YyQJ46PmPwVCLorjBodHbExX1M
c1hevhMSsSiRhDn7xYGfOGozZxhcTyuyt8jFc9T++R9TUIyOVrZ8287yMSXCDvg1+1oB/e5W1vYz
2QYps14lf9qCOrnr3YPltODPv+TTHf7mH8PhUPIZZ1nVvtvolNzkPXOl9CwiBAKDRl+8RoQzeZEH
K4ELRsl+fuQVO5c/nVy3WIVnAuIdkPjoTMtPKIEtkZAGb/PDdo51UQyneQlwTvrJ/ie972jqzuow
drngqxRsKIRJ31oFMLjQuYacFv1KNLkAXVmWvAKwp6f64rlj78Id6+b9rZYgkBrKi1eaoJNFwYjX
mVxgJCTJFp+OVgC2SFE/l5ThhknLbKFWBQL91cvpjBTAQQLQvzDR4q0fsbtFXBk4O2zUzrkKhfSN
jz60/6bLOvWvVHNl7n8k+foTb01ns8JQB5KZkilGJR0x9KFAVFGvNmutH+ewSyfDcRRY0+IW88xf
lzhaWZr3Mm6zdN9gOwb5Q0+bylMUcGesp8zHL8AU3wsCtgmqUCgCC0vSdttGZhpOMyzrT7CQ8BOE
hGcvtdn0ZqCgZEMyDlm73SOrbUGlu4yM/3/O6wEouyAnn4HyCiu0vQOVoYX2s7FABCmZPN0a0ebU
HKB9R23Qi8ceR8OlndS1zXvaSyLmIuu8360ehVX9zz1EFFO5lZ/RpBJt6yB5HJSdI9iHWdY1QpOb
MG4cuN9+C/0gCi5twPG+Kl5FC/tYpIiCRjP/4iNcT5pgvKdbUaWoUNTpsjgBUlujWg3/YCaWNSyJ
bkVRGEsi4QHtzpbOPIxp8aPSA+SmgddKEHBkoufzkhrrXSVHn8iIVWEa8x2f4BuVd3SxpAGe22yi
qCvwJQgWnBH7VvehWDfqfD8vx4E5Xwjlq6g6yg2bwk7FJNOEokKU38SjuccRQehwcutJmCHw2XuA
KFuPgUBSbm4mRd3aHLVFJvKptSz994TI4MRRa8nGFMN1T8KHJ3N2bSmbEb2WikS/4lx0Ptnh9E7e
P1JzWeX62y4RzLQGGWYXdp9Ip9jeO/nlpISpRsoAW4QmHTdZUQ0dGpPL7x8nBLPjJQyoDPmB0emu
BDl6i7t9svWF4njvGzXrBDesy0Ix9mCS9ftZ8JjVeFB4X+gK5NHZpU+yQcY7kL/ClAbChj5mVkkv
D6Il9+xL9Sx4YI+EXeQcny1m9NAoIRdPE2T8xKn1X2Q95DAC+WB5GC5LwT9eC8TU+ggrpaH/H0vv
6GlkNijBp5Gi+SwW74WBbuIrDmosJbymzx2WKCV7JLsvuh0/6Cl8Nzj9xasqcTSoTyWyQ3ZQdIlI
l8hlQetx+MKg9SRbftDGMdwBc9qjnZUbn4miUOKrYBYzeelrP83xFe+G5C0FHM2OwvYLw74key7+
DP93qu5KT0B/0TX7qkKhqMn/qLO0wYgiA5AusBE73pbE9fnLqeB8pYRXsZdyAthZXB6dhsB/gnDE
dEFoMjX5bHLkb0HHehbTIoCDpc5RXIPzW3Lj2jkcyU9qiKocFLXDs+bLzEBJUJt6qpNhtf9z1mnH
KzzUSNibaGQWiKtFhM/Nobv4ioDRKmwIKUAZulwOURu3iIigxYM5+gqQgXbEmyRBtE2k0gIOe4XA
O75AL+ohAKljE9LABK2uxAWP/C/Ku+WiVOCtwQH7LGLbr8r/ySoU3Km/Seqfj9H8fR8EuLfe3QjB
jZ5Kpz+ONjVIDcbiR3D6e6bgb8s4XLU84DPYgQ8dvtUN23M7RrI3AmN3uum6l5rwIVqEERn4vvUA
Wha1lkZV3LRhZu8XfGdhObjdfNpLgOsjkRQvt6GwGZZq7I/QlpLWMNH866bmCOpNokl5ZXe5b/JH
tQK5RQBkv86s3NqiC32EULK4/E0BB0YmhN5Y8nUzPMahyiH6aJ1k5Pp+Onq6dQyCgikgbSKqREwW
b93aS4elvrUcgrAyEfl8l0kHBseMa1ik1rFEdGrQR9AWXdqHFEmKaOiMAusaQ0ye7uiTdNLwnn9T
XrHOsIJpAyjA8XvbX2GFjRULx50b/w+SHDo/rhQb9lj4KlVe8OBOvyAwsPkATuQCRZkPZ1fn3LeL
EJQeLTqVr2NoSYZca+IWk6ZG1xwEAwfgF28L3bJ+iaRW7/mLW79xX9a78BZLbxXqrvca35KK9haN
peSOAfxx7SXD4Fyh0IFL8vsvNVxPYjQ8fYxAmVT8KvOypASJtQRiNbPqTcKZ0RyZM5dPM3OV6JfY
0INu6NJ0Y8p+CE1Ra13XaF7uS96UEB3isEP7IKTz0kp5IDKY8Twf5z5Nil+9cPpfJ7yZW/juOs4g
JscK+Xp5keKCPRg2amrk4h/1jERhPj0yC30Ir/if20gaGfZDyiBnNnOXlQthzw03tA5FddqbR8B+
+Bd6vbUSkrYsm+XhmWFzECzdA7/wX4Lg5t3gaA876KhOKE7RqwlzvcPAOqy79FmndnZL4kPPaQom
QmYHAkLHZmFc2j7QF2f+BubVVwaCrNcvuoLmwD0v0Q1XHmJW4ufdt7rry52IhPTUT57D7umpPnEB
WKK29jCxDuM6lQDmMTNCOCU38E0U70innRgix2oFjJQ+UUZHmxlyH2BWsC/OHkFNT8hLTC14YsGG
5bsksGHCLUHmC8/5aXxTaox4F4EW/yek90dzBKek3C+0YtaROneNcD1/e2+YZYHu+b4MAv5xZh2s
Jd+9RqH/dJdCIcwW4yncRZxkzIRR666WmQD1xusO0MnN1L4jcr+b8p0UGEgL4VoRo54Ioto/5Qx/
Uq+H7NpCiwBlk6w0pj+mLIVuz9QM4kXAE1C97hHaAQHJAH7T8VhAwlgwEJZcUe4UFANt31XuruJL
thP47RV1/9gHpI5P5yXnwqVv3kvxAqL3H0FjcEVvACNY59qSqDtajok1LErn0mwAEb4CR7NbGjUF
6I0L3GjjfXz81EfkrX7hqOkapG8LbPvCHKOEKQOVouEZuuzlQQMqjy/w1Fb7S/HeA+EIybuDnq15
z+oz5hcTdMNCHS+xb/4rzOjlqFHR35nu6TKHQI7+4Ge/w6gtRqhspxzz/gbN8uz00y+ZbF3JwnTQ
7LldgYowm18cLNDEvi31iInWVrMSMsDeg+p/1NBAoU74rfShR9nVDWL7vzXavhOLf1XhaJFi7y+8
ZJfL2VyY5AwstjFzGWhODeqrgd7ptxV0dWfMjNYyZqfnq73FwT4rZCyih5K3poK/x5Pp53yFBZBS
BqU9WW9kGUkCXZXu1LNPr+1qczeinLdFkrn3mCKW7szI23pf2BvrB011P8xTaHJBKzuNerfbuJMe
Lb1x+npE6AjHywWCw6LO39ywlFIro2teqgJ4saHmSFSXGuYIzAz6kf4Qlq/GKUxw6lZB1l23zsmD
rcmE2AuwKlrqtDtBLdkmmQDovJYXTWH524a+6BOXZLOWcmI8Q1WR/92aNwH1oopcHpH27jIMri71
y0ASC17/IezVgYuuO+kGGLwbM/3UInfNYM12bX98cVQUYIigzR6I2c40J4uVbkcWRjPIErNT/zBn
FLdFK7DTZoYnQU4ZR7yXWYpiMjjlR09SaqRQHfvnLYWjTF4WOe406QWVjy1hvXvmmXCqqVD7YD9V
FCeAn7+VepSWjs6RVDtNfz86pKjYiP8+oymWO16HLRhh/09M7lMPNWycmQSWF7BEZi3LV1se1+bo
aZBPmYd8mbq8u+XQKmclWa6d/xPrzoMs4oq0LsU2E6NhYlzPMVLm1fPq+mqPvZpXLWwBJbO/jEIN
8LFj7rB62ZP82rd55oeCeUj3mpWNHyeYSssxWs/D1M5anrywSSWVQvvgZyk7I2kJuDd2rIci6SAZ
EqvPafH91LL/sU4RXuWI8p1Otyo7tFJhTWtPCkULpNK9EOTAiDQlfdg3QDZMJjcGLY6Pn1ttGwbC
Bkd5OH5fP8wsajeX0HHJ+tsryNF+YBqJTrh+wqYdhp0YphSzS5Wmn8rd1vK+b4HLxD5VN8sXZaeQ
xBN9FS2uNW3/l5CP+IWzyZI6MyQD712Enush05P8t22Q8DI2F4hQ7O7gLF9su/x25oTr1Z4dTZqB
YcqilXYoL1fHajppBeRd+6PwGCYiFazESaHwsaB8pS6fCnlC24ewzqVw8cq7avqb2/el6YnLZQRr
nazraGi2YywyN/V1jmSFtQhLr1xdKNJ2iZXjIMiL8LHfXhxMG4ZiGMbZkSvAefE9AeA6bhsTPpfk
wNeOg3ZFGAxyvYKx0arKk0dUi5n6EQweoFeezb6N1agDTUkJZfzmzxoUG/cmI7UD2OWDn/m2cvYJ
ozUNTlZwikmZ0WBo9FxW16USdbhQEvVehI2av7IcmejBjADlZ9jmAUFloy5kH/KoGtKFlFTsm/DT
uwvZdph4xpPp5LsmnEHRGzq4/Duq2S6NuEs/QTURs5BTrksQYCkwkQ/LbAlaUlshvZUycE99b6Pt
pVWyvRfIQ5GKjzsbCbftiL2vUHz3QbHM08BORjOebFUjGM11wtbFSXkDw48SBvbu9RlvX5ODb8pu
i55TwJ2tBziRW27sMU6rjn0S6M6qJTGpTPLBt1MMWqW6fLWOTzelQGzn9dUZx2w1CqiDP4S8XjVW
eXSAEz+7+YKifJa5Xn2QNWZQK7Y4oHcQ88/S8JI6d/T+MfvijzA/lQYIJ4MVRQV8t2sp4MSzM30m
rX3Z/nDjuHIAivbdV6F9BEWthogbrirEw2L5Z5au16y2qzabNw50VeBnnfsh5aoFYO4wXFHpX7st
bVWAgN4SU5dc88u98K7hpMllbLEbbp0InY48576F/UUWPXOGINOLSFReWiP6FEkSGhJZv+nvqIV1
G9zurlQmxviP70jSTcW8ubE/kn6PF5AQmwKg0TPVu6lx7F+f7+fu6AQ031u9lBiE5msKNcY+imjX
Jo70+aYr+eADvLCxm0tXQXs5jaqsvJBTmwZRcHQb7sty2CZKac7vLlsXE5ddFk2rXVu+Pjddc0lP
bCvPxlpuwXbi4AQ2DF3nwgAnaZd4XoQjMfvK3f7suqLAo5WrzrqzEVCBZaC45NLihvB+4L+6k/h6
3OGkayuTDi3wTsT5PXJ3DG6oSDzlhV+sLqOdJeQbm0UzDIO3mj2z/AZTXhCPe2xxG/rrUocKtnRH
sq3hujGS19FfrV30Bv7I6ufiw+CfWYGc0wuOVvtldfmDJS5/SuLd8XMjJRpLL7m9cSCB0vLUSUWz
N4VY1tIId2aXrqb8XKj7iL++h3zabavCRn8YbEE7sFvZKTDxPc5tc1cusIAvEw9uUdSD0VGdv1Mz
wWmEjjlLDPWHu2M5Kj/BYKJvQPCvIgZJUl8Xb4GN8rMIQGvR3ThgqInuJQtYkuGpWSIJHqsgzh0P
0sWd/ZojyHizJm8R3wy+oSQCcg8QkV+YnFkA4ZjyfWwX3CI/6+nlEUa61YhrZ6OcMHMiAWHtMT3J
Gq9ueaz8yUvyO6cXPfDBc/90zP5ZjvHeiHCx1UBzxDYr6we0f19JmPY67Hhzm9QBnFwFQlDUgq+T
xQVWqDh+G/4cJO4XCnv84urZNGnMko3PAwyr+BIaZgSmwntexM0UoV9eke5tRA0V7zWQSOLa1+sY
kbGO6q84I3i2cO9rabXk+uJ45WhvRr4ptedIY9yE/zNlkHhaedoYfwPkBmcb63ULU3rnj8at1Uy3
VB/2+akJye0qHlkpliYJjdudfvMlyObT2TQmUGrJQC0uQfQkfblqu7JtbLNAjMQq515tJDaTHOQG
7ofXbkgR5ZEVnkzq6i9DQtZ/c9clKr+pmSlsSmSvFv6H8mU5CMwslPSnnEeXTtlHGxfOVipbMlqn
IV4A8OsqTLrW6hevezlgbAi2eh4QZ8UzdAGBTo0UgBpSQFW+qoie01Gc+6796Aojpady78NBTFcX
ovfErVcnz0Vaa4lyWAJpAjhDsmacOqxeNu2E8bMTjkg19yWDiYxsfe4mtDsBOqRefk4gxRPW56aL
aFK/C/DKZVhzU7sXAjSNh47F8IT6YfkKUlJhb2LrEMTn+X33rIm9QsIMPAdAwSaZTqk8JGzme2OS
VnhXnf+oKfvOC/n+RKVvn5CrDDA7CRUd87gwMbz2ughysbcjJkMqD2g6lpWbzwwFjOlDeOwC7wyy
WXLohgYLpzfOURno+czH853dCwz9NZRwI58/aZc4mkmnk6WWwQBkxpWcTl9RYj1nGqXFSu+HiKnK
SCsP/1KZAbGyP/CZdYVTq/fK7Fk4ExkO2byIebHuQDXJM08I0mrPYWpgiqqL+Wr5mFNCUZZwtoYu
/ndm98syXFHciVxBWUK7XwLwbgkNlv4kCWr3J3VxLM702QTV0pgwgJChbaaAUklvcJ9WRjuxcghk
RbIhgVmTJiSGglcAMHiSPqsGoR+ez0eUE+tSJHQ9uF9UGH7u0MfJvVVuLSryKbMHRv7wqbZMbxy+
WIpiACGqJ5EHPxyFWN7FY5QzsH9mjPnYd7f/CFSZxgHN2aqBNp2BlYceCmiJKlI9787/J0UiUtQR
kc+PQB3Hsa6Pzd1kFigPnmgH0MRGRp2joxNucCjYR8peQx18AJbiXZXcRI0rvGaiMGCEBx95yTB1
ggUa9i7R1kryG5wW69sxG7qIkInRGWvOBxFmj95DcOZA193hBlZkruDj1Og3e/OIo5oWeIu7N3Ni
jPuiKzv/n0NDIaTAZR7uoNJcaeBWEBzy91tyMoi7xT9bpzElSgqSydZscqWVgVBwQ1Lm9HKHUwqr
R3JSjgpYaJh3I4Sl8HdcP/Hpb8o84g2jh1LRHA4tpYAb8BtsGr5coMXVB51MGUXt614oocagaxhY
sMfBQmgRmHCkE6a4ktKjLf+sstcLk0tQ90J5uHFHSkZYFoYWehpubvQdtGXJz21eauAl6vWWLLF2
qXt1Omod3j08sKkZ8HWEMo5chtKVfOFasSB0d/21eHK6xHgN4bhy6Vsah+++/B3HUj/OyN4Ejok2
D28T9ZeOmK5FCl0hF2VAmVWTweB6eOUrNVkM3D3KaAPWmfA9S52xQMQni9tkHgSbjI6re4s3vttl
yxsMV1qO9tGm5s/TfMwsI2Yc6Jh4CokR7b0/i0iamypsD33Kj9AIY0soRh1zte8tYeCpEou9UNBh
Dj5IbvhzNnwrtWs4x9BRLIEJDHjO+fpOLd1H2XmwqzNOTRI9ePgTTutBbytbmyFoiFJctFSKG9wJ
9TTj3cQAwnUgk3+/5Heu4aWVsdt7Lia36orQ7CyYv7YsSpcIOkLECEXoOE/GeAiWmzqISfieB9AN
Qw10ikJQT5q4t6curJiagkQtvOQrRBnZTWsIm63LUAhsJGtUV9K6oRfX+ZotCgsHASts3s7kpFoJ
kabzbLNGBYVyKT/Y/0cppLaDWBU5MwW8xVTDiOPhhYi/UpIBEwXKE/Rcw+8Bj3TLrR0OD9wQYHyL
XPz7wLPUZC14nMLqbSME+6auv2GavW45cbbueZdZQcma6/3kp1A3UqqUx7+RiQO7rVPXeWuFihb2
2JDQNAO1FXIelqcyp+iU3hp6yavKC5smGenKNfgxac+igZGDTfQ8WDQLhxWTKlL1FicjVdGDY07S
Qt2gaoBaavakZTajmiGYeB0RpD2Pr3uJA7bdabUV3BZw8BUG0LZWRY7kev2oVlKLkekJdn8DzxH/
c53Lf/FpRBhAA3gASLdn9gTofk1Nqjtqzmtzib6DTmQbSi8XIKhbOZw4zZsdcLoirW2Hgn5EXtlZ
3uHcS6318I/JAAFi99csWAYCE+Q3ViF/XPz9nvNiQuTlB6DI6FzSgXWp5r6ttSGDbS2dMFcNw+Ul
nY6GTg/ZvOquM2wWz5DeTZktklSv9bNhc93F8/jYDcfcGrHS15J7fuLVRgmkqKKLfurvMQ7GMRNw
j9XGHOnNhW4Rh3w38KjzxS+gQhNAXjOWS6Fv2Zb6Kw/uAuu84a/T3eEbTXD7PsF/5xvTmesDFcXY
l9agNjxFyvyGyDDloe++JGaDT7qzPSyiESgc2mDMGQWh3T6Nxb67jq1J1l+RoWFVWwZa9yLNr8b2
9n7WnJ0x3bWh0Rt9FEHRKpF03osrRTZDuDxcc8BRm7EYaUK/eJa4IFxW83LWElQBDQ3J5lJ7yqXT
raNSSI25O2KoMHtWK4SvmPlRWDUKT0yxi2oM9wugewEMQ04kDN/+ewsHwQw7h65PpMJf3OymbQ1F
8Z3lNqn2Q+qVVlDZpZ8kp5v6l64ymYAtYOGDR9SgBuOM5aLSJVCzpMGrZVDEphiWfj5IAZqqVvT5
pTCnxMvVhlgFQyaq0LkMcQMdwHqCzrVEb/txXcBFautTFmUYuovXLLKtrECrrqfdSYXVB101bBVQ
c/va7Bb6MuM6UIKHoIiqEJeMfvv/2m6lZyhxeu6AYui/1vLHFlI9MjRAFE+fwoBa4oQU3Er/qLEH
iuhny00Y406RHKJXfYs1CgaaA0gY7IctTaF5CNGUBimlIgstwVilhC9gmiR+sH9fwQ+liUukWV4M
fEiPf1srW+0lf6zsg7JO0MU7j/SX2UXlrAkCK06S1f7jt1duQD65FuoNKno2a97RIK+jWZ5NgoEZ
Aqfgza/wLMXXHWXENzf7whvipmKHH1Zfc8vDkvNuRhDIbwA9JhTwHRGP8Iktd6g8DpYC3P+k8XWX
rucscFOj2e8+UvYSFmw2H+TA1bHP5XoyylkaMPiVbzvHvd0pvaO8cGI1oLsf46YcjtZ2nu9rfxyR
nMaJFYU9fOXEJ07nzxt88F05CnpQKCLHQc0qMivHbYIBPTHBrJv9ojCjhKJnMduraXQjMhFveB02
D9RatkpgN4SeAQgsg19RblPWpa7ZkJ8z4m9sOYrhXSNzlAwOFiPKAeWwddYEInICpeu+OyhApuQl
g0Ue5pjuBhJThrH8Z0jRB7rrjyW2nvs5WUFbr6Ks5rJrZ/nZlBRU/Jxo95x2d2ffrEXuBQ9EiSkn
3bKwPzlxBzp87Kr9qok4E1DeZ8GNRCWxI2dHN916J1hFWtb0c3QAanOPaFDG2X3s/JX1SaRXt/bx
P3Kyu4FXv8te5KAdPIVlC2NNHpdTX97tbEjnDCIJ3AlT1RWY9eoMxfu848bsgv3VU87gDx4EtvIB
pEOtbGnHukRMoIIyAFFXxq8uGTALP5SRXgalZihA7Kxst36B8bs7JGYnHmhXuioB4SYTtpCl15TG
FYwzXgw8Rek/cRiGaqNLgT48w0gc8txuCE/RGgL+QhMXhf12nAYgwR5qXCqXjMKcy/2tldlOK30f
eFmMmUrgcmTgGPiZwafhyr0LKBKSUhcHi2XVcg3t9+gUece6twA+8tbcKq9SI+mEAe5/tfB3CX8j
T31iT0CNa7gWx27jfk4d0QS0ZnodL2LcdNCyg3bWOxFBNvystk3ayzwWKFtKhHw+eXhzdRAsKh9i
2FNU8CsEzmh5Ug3QiCoplFNnSBnER6Gl7/UDH2OliXLxl5o3+S008yvyk8/iBcPF99z9JEFJtn8Y
KyV6gNO5npei1krAVMupSQ/JMFmA2RUtQzRUq7juZ5cfWzKUuNmWAkvSXvZCJ46Cf2WPNAyKQUVP
V2G07/26oHGW2lc9MUnG62wnWnk1759v+U4idDC4ePTCrAUxLWrutWNrfRmGSUEG+DpvSfFoaviT
P8cs2U6cT3qk+ptaypStbtA0NZpdYeTDFoEzmt6zOekAbp914zm83YF4Kto7tnE5ShccpR6btoUC
oT0gIWxwvyQKdnpa4xiBLS1o8Sha+53FIHWZF0j2vIGE6F2ptSXocrA+PAVN/8QhwA+holzNg+wb
m0toTSli9G3ZSU8hGYqHIuaS0DvHOSI75TbKa0rzcuBJ/HLli2tCi5HTeZ5d0Ev1aWeIJGJrFnS/
tw8JxukftKI/FVS+u7jWbj7nTZpjDDL1beQJcSDEa6xP86SBLZyJLovxOAV2SapbNi2S3c0E63mp
bMyIn0q00A2D/huuqH4GOmWu5hZ31CudduZ4BAu+8xksY2N+hqSH1jEXQIscJbdCCh4vHYup5wHx
SVzGBN427zLZGca3UQ2vS7R5N/w6FSqgHBi8/bV1j+cFxYZnP0A1oXav1eYBChEkanE1dkgLecxL
XmUXqBvzA622djpUNgL2Rmx2FYoalN0bk7ppcm+nGu3i/AnelPPkaTUNQxn99KzmKKzA0KFzF9Nl
RoMO570rpq7h7BcSkhsSBffvv63+MS5F10uu5GhDZ7eFwEdqVZZ4ohXGFVPIunogpIFgkdtQqtWM
Ras2zEY5b+93cYFFFc/Fo60NqLN8cy6O11Ag3zPiMF7dLq9b1voryitRTMVdEyURrasmzE7ICypo
zGovue9gKokRD/mCCDvdUv3XVAwzThNLW58JZNP33lpxix9cDZvY4kBw2yA6lBj3ddmv5OyIM2kR
R4gVI8FIitcIZkAwizqLnFFLVf6x2xx5m2B+938PwU23ptFiKUosXElCvqjPI/0aWDnDHWkY4QGc
FsNQwD03iH420ju4BnLzZrInZbJRig0jV9iMWI+9JZxqqpVdOhcEK75XrWCo+PSNBU/RUK3JFWKl
rYWCFXK3r9ZYLBjI033mj6pp/6Nh98D57QbBeWX1srXftzes7bZ7H5XBVNbDwITn4I3wkxe2+Ekk
vU/zKz6AvV4Rco8JT4D291AIokxOqOgDg6qtyvINidebKEMA+XvH/AdBLAvyRpXZAG/4JcHaPlpR
TEKUI2iFJt/w6Jg7jzwAL2oszbZTU8XzSEu3Lg+cSTk6iW0HQTOGhJyaJoE9QMJE8UPKBW2gW+R5
v456WI2LIMptF6GNyzq4Dh7+DRHTGKI5q0rH6iwcoZCoU2xLoAh10rr7i/1uk47wNUqUoeXPEMuB
75VDgBcKCVhHdrsW3ORar9QL5ySIq/1UT3j4U4nleVHV4I0sXJprmjP3OElIB38q3KIY/ZNoYIfs
KGARFTWvJ7/BXDI1vrLBBu74XGUcNxv41VI9rFSfOW4SZTsoeTbBPS7m2bpw1fKBzZ+EOpXmDs2r
Su9UZ6RxlY7Fw0IWm/5lnhmW/SNwQo/5Lxhrj0uciPsZcxYkMpFhGTPOz5Cw12sPNl8Mzan8nJOO
EWjd1QIy5EyBCscqwRB1SxdOAGJoQn1wm6UG00RTDkSKr949n6+Rb3m+Sz/KvRPyRp9Vz/2fQGfR
dKbgxA5kjg2KaREv17JfXd0cz+pKtSq2wamGgMvbJLsQ56S2IJ22lEReJhdZ6sDQkkE621SxFspK
xUuyyOc9689FckDK5dwAvxebcl9bR7MPPM6pcytLSdX1Wz4K6aOBNoAxxxxnzpRVAkWe2dmw51Vz
fz3jIWzH4BizxlFAgDFca/LrDbQ7WL9DuMRt3EXwiogM43ItfAxCcxp5OyCQhKTHe+j55lANPnqP
rBpmCqB+tubZGL++WPHE1+KhQdjg8w6P/l13d05ebejtyD0E2fDxu1VhBFchEhNT1MU426ui3cK1
nFkz8dm0LEMD9g7UIykaJ71YhvooHr/kHyPfmQB1GtUgZpS3pT5qwVWTOy1RhhaJ9/ZEeORrQW5a
a88LQW06ic0F1c8V+8ruTV2QfyJbocZeN058zdnXs04+PpThtUgvOe4MGu1hlUAvOxNb97k7jxH4
rj5N7OE75xTkYab10RhzcQCQEs0z1CNws2d2mQgBQtQ88ldz9bvjW0ZU8q+jI+5l+exWKltLqHNq
u54ngi47gTG8FD9P5BkQpTYRNKlYeusFVymQh3cJuDUBZEk4jzsGG3zF7ln+YlWWXYzJLzix8BFS
LEzkfC5bYnlrf3oqV3HvSJewlVxTsNFxsarYU94C1s2BR/QajoWIr9uAJPptnPFWMOoOwJYM/eRu
YGf8GFEwlBWznqA8FTgGaZYhGME2hmmYUsSEMnYwh4sheEoAO7IGq4oBgQH7755pfbEsG8tKcgmw
oucRWArURM+dRTANZwd5M2JSLnvdjSo7xH317wsilHeCSMPM13p/8Ex2WzyWngy4eOMnvjyZ1PZp
1kF6lC5K5K1N2PQebU0pFhtsBKOdx6XT4FQ8p9cHEDKVSKsaU1o9qzKdHptKIKjYc2W1xM6PAKOE
tSp0FRUCQMB6jqL0ZuvgvyE3tW8pMLam4uyX1r4CmYNO1j7NrusLFVFPsHlVVOAj7tMwV/BBCLdz
DHGJiBwSbLxhT+qMrV3ffklZ7sbmKitfViuClBrzdW5IWvWBRLk1SJJxBJcCty639ED2JjhXVeUf
IIztkYVayY9LWlJYkzLyPmKLamN1vO/yK6h0xbP/Ddc+Cq5sy0OgA+DNim/73zUyZ98CrFsZnXkD
6IjlhrOdz5V/qgKQYr4vhbS6jjTuCY5qxMC4xboJx62vcSbXaaaferEBSFM+dyhA+MO0aiWVtXm8
5EhsVV5skHZVSBumK6/epgCsAltL4zesb/TnQBRIPDbLb3L0nTNZYHxXJ4aDTBAKVCj/A38r+sSO
Tsv+6i7dEHG7L7LxT4Q4LIghnOv8KVr5obPdw0BJTFcq+UIJUvMUzmAOAEKRIJeuS8+p4JKkiTOe
dIcgkjjal7DBfPg1FIooBQ/YagytyqbKIEKWzbszLuh2LyEi77QhLF/KBVVpzWaI4XGb7jX3iP0Y
pykRRmXxgSjdmhA8A6VpZMZCOQjk29/qPEYfvJdzcKOFEaTSnyDHRuzJhYP6bvBkbj2mZfW7yJVo
J4LKUJzS9EnAjwZkRu0ZPm94V+xhrytiaBq83fHsI4IXazrKhraisnCKVUc2BlhlH5EgEtEX/pTh
gY00LUPjFxgWsMI5eNc59+hYIF/4gPAkw8d2rZV7YJzLXVPzGBNlOU2/xlUIpwtobWBU/6JLLOoG
BxJUG2iWWuFiObQkgmwAt9cPcZanFzwbFB/eZ9T4euwZxYLs/M+Yveam2GJ7M7PYZMVr4XoMxQQ3
WU4IKSjJl84PEMZqa4GlwjiGpuizUGNyUbe6kcdG3TimXuldKpyKu8r8aRPjO41FYtQ+Tqt0VFpD
aggZjnD8LsuriONs8jUNgaRGMWDl3I5RGUEOhr6NB2ntlkYPhaO2O6WhaqkwkatDbUjTzpBZ9vlO
QzWn9TbRujC2AMR7TcfMvH2YmpYZzYWzPD5iPtJMMIxQcGGDB106D6Aj8tXIawqdCMmz3o3DNl0G
48vjlkFNjWzZZqR6zE7aIidrA8XNPQUFwt8BDz6B3Kg50r87V/7kXiak34u4KBUaNaP4O9KtlcIo
qSS2zC8EkqU3UefHhKGNEsxiFEhOHnK2cV3BqFV/zSxaYIgPlwKYs99WC8i+5ze1xeg5h0KnOk7A
Gs5B9eIDH2G2A9wWYOqpC0AgMTc9VIv+QKnQ1Xpsr8LU6neiOScxXeEW08lMyebt1wrEyEDit6mN
7GjPHAaHS2gQXELozt0Y44V0IVs6JXvLD/AmwbvB0HRvsA2298bDcm3TGHZ0So1hhiEvo5i9cf4d
IfFnh+7N1wrQuzYGD254MqUpgfTQwtcv2FuOfC28E9VL8lDOe1aSDY+JryrRFqtGeWnBoccjrOif
MyTYSCq95eEwxGAAE7sjN/SGz4UrWI+pTWXJy4lHuK3rECJX7M/NGVsra/REH5+1YggJr/fBjqto
aujXM6qjk3kX8JtDXvIrHQgyrm9yxK0u8SHlHvJvvjdT+wOQhetVrFLmyeATqWrSLKfwrs6WB1jR
CR9REXsTG6MNv6B3f6edbF+AHEUFCFsbfR2PITJAUyRHX3eJBVirMnqQfOTOntnyCaAXCGth0WjO
L27R4B4DXBLZ9uzdv9YFqogSLXne1JGFdXXQVPT71Rz+oLH4VvDpUDTvURmrIaW51IQ0VLtS7eFB
Rxn9ZxRRyPeX1kH1q69NPFhJLLknk/8kZ35QXXU7DGDS5Ea5RC2nKDZ2NcEU8Q3L53jI1R5XLSB+
vtvh3eZ7e1Cbj4nFpf8QZvIr0e0QHZPTWvHsqnB4eJbkdF9KZyuhkmOlOwPpapFtLZhH4UT3aggp
G4KEUoD3If2DnKfc7JiNQNBdA3jEKZrrW6dWiwpaiI1FeBEqe0/ya/qOn0RGlDKZfV2PE+Jd1Cx3
fUy/iIneAdcOi7gvME4DTiBj2XQlkVOu47+QAi01jWUzrtKlwpNCv19aLmpTKXtYlK8FHABeaRvy
QeQYdntN0MD7O7fO8lml7wL+3vi4CsrG1QnbV9ffOtxRuVb1jUIamwiXXHn7hNvOaIXvz9jybL7B
LR7U6iR502W5ztYX8YLTwTmsv2FyV2Ax9Yk8IIt9nAxE1CHmDH90fvAs7BkKbUdpranxGR+47i8m
LOmzvRKnL1SkYkOSsH7AvdBf97jzrZL+FLNS8wDvprAowOiaGrfU4RjFR4anuM5BLqqy84anwlNw
HtyDF7g4LFVyB/XeY1Nb3ioDQzocs7dd1xkereawUQ/4iEO8Sys6ZhXCT61+LyuxLrT9353at6k3
MgqFPOGUjQRoBI5IRGquz2+MEwH2jj4epTo6qFYsu0foXD/fRMHb8hN9TicQ2zffnvU7//tDWREF
dSM2z9soKNQHSq2B/YirECCOuiiTdIPBOYimPmWhibIlkmSd2CschmzM/gpnw49KQqH/XKkpbRLE
rKlk+t9IuvH5s+HyYREd6GkxGtAbEitEYzvRTgshkUAUJTMfSgTbRUOz4BBy9jqHEA8PCg8pFEkD
9TOZRFtr35d/B9q8buzsB+eABiUrbsi9A7DZh7NayTjkRLOhxG5iYYRiThyYS+Ma4Chj+5JF7IWC
7IBjxv5RahYvhMRCLthoCD1i+bodZP7WSLvOr478oWfOdpMjvLJ+GOs59HDAseVJ6rmJk/FOSDZ4
WFVR1QVxhujsekGOIPmVmIvgoU+2ig+Ns8YG1GnqtbNQX2DYv8aPYQlZJRrM1X06/IoESxf276Uq
TberR7jZZb4sucAVJ0eEbFVQq/lwximSstG8VuiXUZxpZ5o6dpC+iZTqnl8ABwj24CJgx7g+O4FZ
N89DEPM3bP6FmZyVtL0ASawB4rU43E+22zVH0bu7j29V2FP22EhahDtPDh5bNflcxY77MLu2g+4x
kZXTx0sYc8lCXuvHx7VlGRLzKLJDMSggqqmLAda1EoVqUpM8/2a84eHe6cZGGOVLkj0/MeJxs/mH
AarpMy7aQFfb/xYXhWinmYoghFed6papkrP/c00oZWKBL9QPtiTa0Evc/KDY+wJPufnm0OKQSXVa
ZeiIYlhSSCXABXpSTLwp2f0nRFq/UO179YP4RUK8FSvjo0y6LF40Husu7bBoQqfh4rFlXufkOEOr
b1PCMQvikL5lGX+i7jKXfmf3I83TxN/OBQFFEz5DYk5bI1Zo8nh8wflRUHfakBRBcxXTOg7uMk9c
nwX+amdUCLiPBzTgeLzU72FiJMT8cmmtJd0Ak8mQMF83JM1S+ST/OfPF+Hcidby9tiFWPaA21x0s
IX/twAf1+MhBJW2fvwn8I9EQtbP9XL6kq2rX8xXQi8FPINrjw1Hak/SRjXgFLkVZ9FMrCPQWbZeA
p2a1J8cpmEmPugRoFRQnNE+h+4s5sE/usbsfbfS9llcN4PYB7IwyD7KN9WuZruK3CFeQVugdDqBK
jpidUzfitiYtTkjswOSTS8hEg7kfYteDkqWEzvdJ/X7d4b3JtzrtMWAtig3V3AQOSvBsFAxMLJgc
0/2gak8SM8WYktwIaSBeleocnu7t9DwS8Af+j+IPeyrR4VSPB9QlpKdyJVVmzuqmQ+iruhX7wNfO
AewTYCD7XnTLIYY1fFTBD+LNl/d3dYV4b/+oMGrTm7yG1A82vpMdyc9arEqwrpXWa3GClxUIT4lQ
gM4dwso3D52S/H0yWRjE0LAGFmi46gQEzlzQEUHBnxd0uj+i9z1rFybD0s6H18LQpcHYs7bXneZF
MIgoln1wFdZLFfztXsi+0BtLUxvcRpYfnnEXGIAGnw4h0wo93tFIKiUlaedH7+rXWTiyoIvVD08G
CH6jF3dJ3Cl7Hb7rsDVbkRGe+S5hEev3to5+09vn8ZSAs9iCQCHPiAiYC6mIAP2U7auPvNTXzypw
3sy6FJdHXSZGc+N9rxKHkqFp5hHEV4krjJD265LY9QGCQotWgaGV4yBznFgmDprprVMtoK07BD0s
BBGfZon4RA5lrkv0y6gi7hOe9Pg3bbYmpVIgtZHZJyfKT+Hx4qB4jaiWDazJm5duICDwr/JV3+qy
FPEbcQJUfc1fzEynDfhOVWwOrfPxT2Dtkit9Qht7sziF249SLmF1fonoMz1nS4kzPIZBtYCl1Dlj
tb0s4XSzuPmigSZ57/3G7TrM5gwxdTFnU5xgQ8IwAALMXdiKsOPKWHg3EcsmoJpvHprSRiU2zvD9
MV8Iylr0+Ca+DF90pWxWQtA1sqSDdHBmL4crW/yf/dkuOnvwFvWitk3V34dvc+tFiQDjXh0fbflV
6cEhTUWINBI0sKS1MGXDnO31Wc8kOEtR+yZoOjrCORHHX0DIGjLDnBFphrJRZNcMCDB0iV7K3Sn5
Ewt1jR+uzTnn5B+0Djnrg/eaecWDqQggCjS+7W9hectkyXZFif7shEu/tWDIol8fsdZME/GYEumz
3GkdpG7m+h5UF4dboLPuWHPLjGUQarG0hU1BgYuazKxIbTtmPB+mOYVQPgaLsd74lZHpeswqK8LU
dXKLOeEd/Y9eyLB3rxQHLsGnvnb6KzWmh+aJUCQZn2kF20yghMDeXRD2JbAkfBEPrJOcmP4o5UQx
jZoLBZhNdUhYAq3Jak1oIJ36BNkZngXqeq0Rl6ASrgk1AVjqrIcLszLu958Ebmr/1+p4Q0/fMTVh
wj9xExKb7xt0JY72wT5pL/mzNTERuEkieLf/xRYNcx0g4bzQ3Ipdgf8jPANwkCvzo3lyyM3VPfjU
bPU6DmPrDj4EB/6Bdgtv+lGGg51K+Q+M5TAlhlJB7hW/q0JBBrMUqDS6F/qzgx/rUHO48zxvcjst
33VVhspLOlSj5CaVlV6PRXXps7FFlr+1SD4vX0lLXOzf0622URYA6zGPuBWzudu3p3zpNzpU4UmK
1iMMnr2KroxL8WegYkWOuqcRGdAFwRXoZ6pGggdjirBkvmlMRkC1gCyzL1TV8nCeekzEMCXGhwpk
17YEkGzclpaIDg6G0lSPU26bUjauDcwZilq+wDzVmp1Pfqx78FvDOLGI9zkfUMSXyWzLY91SM4jm
+SQIyNAaQBeUWfU/aTIljIPMvzkAPBw9AmvJ3wZLmkyWBf7sqMvKSzPjAaPDurRMZNtMZP3H9NFp
FSjZXvghrOY4l9R4FLktUDclOpSXlBaH8lZACcznvZVUDNWcwVGZu+8FRCB9f90gb29zfSaYnTqc
k2/FUzsYpQPeRfWHGxN77jOtUuBWZ14UTTvHtxSCzl+J24NqapDcnZzAl0k7P3+ajZETkYx8b+RG
bnV+WbI47IltOcMBtjo6uwmgCOAs6dNePZAo0+F9yMzycOdt18oJby2SmlW4hQstL8foIKWUKVBk
faa052r7OSU1KU8coYX+FgIh0gqlI1pMjSbqTlA79CMBTdn1L9+/PO5Cg3HF8C3c8ECoht8kmwAb
20xTc778LfoDfpJw8XDBp0sv2TUjKQXH8KTnWWWX5zHjBbgUenB+CLSeODc50JTXthS8tT5RSTHe
N8aEyG80E2vNV7P9fYbTWqIXGUFSjvFfmlJdeSrdly1Pj51FEtPNz7ZyBdXhpMOuNBcnU/PezmFG
SO5rNkaRToQq5/ABuDs/xS7Po2ehCQarH3Tjkpi1387SXM1fzXjy15mjzbqKURLb59UQCMtoNL6V
2dG7J/CeJ8vkSzqXl44aogP6KOCeixDCr3EpOWVBcyTUilwFq1SqkxD5/csz+OxpOuWswwAbdl2y
WmVkme24ky2SQov5zdgT2F5NSQ1UETEA0WaHl7RXzCsMxFhJWAisucLvhDO+btOjFiXTpQzSNym0
TunPafu/gsFTdwbwa1xigT1WJKGd0mCtwLK0oeh2u/uvmLlRjQwrlND9Qcqf4pRyCB8pzrMomWhA
OkLq+cIyp0Rh4NQtk8zlI+O314H6WHVoiNgl38N9Yb3G/t/sR0CWg8kEiywI94IPSuwttxsqI4m7
CoFOIh4uvd9ol/KQnNuKhPQN6vwHWhnSGI5fa2pm1Mvq+l5yTlRr6Xt+aEGcQGW7rRhXIgNGFjCV
DA8jzrt9Gx22fFpSAzgsKo1Zu1sGlLQ7UPmL7WYnJW98rgRVAmXtmN2Fu4akx6/+/vM1+xcDs6V/
1irkQcsguKlpWTaGKGFX6EkWbm3FUZxtcnfBVoUVk5dms+A2DjCGlxdq1Koj1QrPTFADDgyCAWXx
slztG3o2aFgxRm1d2JlqTYoa/fRV39KKdctjYlRCYdvBccEFDYO7UG4VFkx8A2As0O5ZKTgHLmK5
mUaZHWzAtEVaV3rqYpOB2BFqkWEGWnkgeOez89E+NtLjI4ZYkJHU94OiCuf7YsBkp43/eutj0Sfq
h4/pfyQlPfPVztOx4e/Qeri2vPKUTYVUZAHLRWnEEnACScxxBHaxkjcBtsalScAwekbIbqOEB23t
h+4EpLJsOnButxC4YXeATpWXb4NeHYGpkgbHAaTCYvh8kzdLqm32NKK18lp5gTTdAuqFx57ZOsD1
UesxmXbm3dh5QR/2JPV/pkI1OOXywuLDWRrS9KjqpF6GfnXSbMeQukkKJS3gqwU1f5rxuYl0buyV
thqLn9DVUL/Z0lqrqMBeltiGTem8tg0OJTKP2EC+M6ABdxQESwdB0EzMHK+L5/FaQzCwokKltv/v
5lzOJMBCRUM/o6E+cL4KhEfgH5UJrpKytGnrF25fk+4CG8xXIZ5dYIR7Pkrr1Vo9TdxislYINpZl
Hrb+Rt51nWUtU4PoPHrVSP0wzf9TuY7D1as2wFOjJsDNOHKtXmQCr+3L7bdBtRkexusYgy1iO994
CGzkglJ3oOO+DPE7h9jwEUsZP2+Yr5L0niXDQsXlPdKDsaZ4T0lZauegxeKgBSoOzvpTvCakgrHP
nVoSBW5UMReRShn5FjY1QI0MgJF+y15doNB9JsM8g0cWJYMCwIBrBKAMWJCaUpZIkbwiSMQWj6bi
7WCxCb3vb4lB8ye45i2K/SShujSDbXweCL7BGF7KvDpzvVH3k8B1zE8b62i9Fk+mCleYFvLLp9s/
lJ3wQ2x6UlVDAgskX2vK+s6ZTuJbjs7CJldwd/Lbm56msV5AMHF/ekZ3oKnRFBvZKN4hBBYyEGMl
y2XF4PHIOCc4p1dfCVgqGbldV0jNNOcvNikQCG7j4MEZI/EBMcCtu4aMfuvTD78VcDneKo+0cBTf
5KlnBwj0x9nzJq0Pze/Ltct9x+hAKLLhkpIN7toMfTD9Nh4S9SRaiQlCNJKf0kUBpjh8nRcM3CY9
WMkECy32Doxc7jTnbokaJ8xtQzHtPEEsTE868kZJBqXKzzB9v9F7J8tPPdwlgcmf3UNo7rdOCQR6
ekEKBzr1KzFyK8FI96RF1jgBmsxGmjopISeDXeuaxXbAOfwcRZCfbEb5I6Wk1jVdEhgxYxcvvLpE
ICf2bcz6WubWbNYF6ainAGy7UjII+EQWNaWZX8C/KDSkqSV+e9HNPxOM27xgvmtWJbKZBNfvYDK8
h0Ub7ZE/j/7inNqlL2oIERswUuGyexIrVP9SlN2aB9dqi996TzIUKUmXSQ6u9nYtY2sIi93YGam/
ANOsasVeAveICpzec6Ykk5g9ZpwpbwL6c9LAUFzEggDx8Rqjn2F8nNEMEyIP8gGMRLtILLy3IlFj
tvQxynXqbO7W2dMpfC9W5XHj7FllJwDv4Wc6nZziF1TPh9XBvFI28T0yDNFD+tS30pRLak32WpFR
pfNzUQ39bnEJ5Bc+L/Co/dQrkrcgmBYOUokFpc+1pnXd47KL+sOiQOpjBBRbLqp8qm57n2wGqLHo
Qo2eAfyvQ0JCibxSMLPesIX0Qw7bhU+CbRV+D1bZDWCEXn+eFO1vGH5suNxPBFclvORm8DEtUhsh
v4NeIT6tDCUseF8heqTDkAbFBA17pZ9ubqn/LeOEE5SZmwuDaSbe/BD64KT6Yh9ltLA4ERa+tUOB
COsXDOm6RBP5WLrvjiodZz7P798ZLmEvk6hGaFIBizwUcHdtYL04ANiLh2Fx84j5/sPGL0BmsTAt
PLbnsD8MpbnPmF6CY30fHRKyOY0vjnhnvRgRgvtHu6uKyTt3xNKXK0gqV/B8ephULLimxPSsw/HH
mUsEpZeGBi30vMb4ACssIDk1h15zfle9CsQxsqVFz8qTJE8gxtS81x+Oo/wVtWJmFgiDcQ+PPgKz
Q44oocVu9H2UQddliOqICnlHhN51A6Ut0hutu3ElBXsSxZ9t9V2bhmDWI+cw1wOgHP2JRHBzYJ/U
PFpYbpCrFUyZpuOm51QJ3qRWHpz6Ow3hSlgZzE7nQq3rHXVx7WCtyt5Ly05Zou2mHvdERpopGfIj
rXJgDSItS5Pq0syXOlkPZ3Xp2poPpPzshT95TRwKh5sf7DptHFmZWtWI4ZndrInnjkiHtYZuYoBZ
2ZbxSl+zphi2T+3QkPb5nC+gSManiDsyfrnHDMLEK/7ehpVqQY1ambF/OM1iQZJn9hsnWcmhiXEL
rawLKfn9cvKJ9fuxKpBZbyktpdeZD1+Ue4kg6XJdZBg2WuHhZi6exbAs3GcWcgl4jTpcUyxy/JOz
jxhN08VVPioOdbP6GSJ7Azgso4Wmv0H5GKX91XPK9vPsIg36I6n8Tnrhw8/OKsd4WMcsRxNNNYvp
iENHIzaKDoAzPG75u/SvSzYirvrN0u+1vN71x2C1kC7OaC4BTZpFHgNtVYFlaJjbwmoAI7dsxwGu
A+NLBq4EYuRduea4ywbvZauCtGc30w/0IJTwJaGBUH6og3twSfAg3tV8/roNiot1li635z2PuqeP
oM0pdsBMTof4WRwxBjwNnJQ4WV6kaMMrOgyCtZyc4dCj63C9Lrm1LavuPvTERSFpB4YvpCpHchKi
C36WR3LeRmWScdiGPSeW9QwUcszSQpF1+qYzwPVRs0aUANxPmAnQr5qkjSv/nkZJGeXu3CifoFoT
T7i+c1RnH/xGua2oISXrF5Sul80M5GUVLMP/kYdhqc8MGyu6rhaSx0/mzgfRtcpNuiiKmzJOBlX9
j/y54+BB4NygLF1D1vTNoxwyfxnl5RDpibIN+mnVXf4LSUcijKjNSgTqEtwedTjVs8zy3i6reo8T
xaUi1dRFJx6No22HFpp00zFOysZu7NeHfJWZxtlzOeHVdFrgIidmYHCBiqXuA+HB144HvjEF78yh
bplTX1eVTU6QwQPOdko/3EfET0bDDCmSE+XIjiWXPyJp26TW3GjU9p8QzFamsAFsguNyOYLoMw9b
Vhzf2/tQVzmQMugdM+Yay3lOg/v3hcK01XRv2I/HiKQLNrqmTOmpacmDJqxdLRr8goylnD1OTBix
0k8v8mqvJL0d8Re5DMPlau0GbgbnLl7pdDFkBPi58ygVxkEBnYP0NXaaZYnFBghF5k062MiZxbjq
YgZQ/huI1zZf142fq52c4ASbY9d/v6eUSXbcSJMlI+iCdNnhmuLVWxH8yQYaMUVMsIuNHgiATH41
NR1G6QxRfVNcIJd0ttmcOfwUBNFKCql9T6wYUCFntVInZXh9jhujW1hC9Apydm5IKslTH0y8Ssiq
H/KuGIsxaPeIOZaqqgyTDvH0aedyfR978BbH0cljrUq+N5R5Mzbf6qi8Jl1x6vXbTaJBXB5mq/xU
TrsAQGygAKCG7wpEbtO/YIlme3CX69ntBuDiIKun+XKi9d65f4LLQsL2+cN84L2kcin32zOutsDF
+0s6kTzIhd/8gn6TJD8q6+fSHusxGmuNBpdvzWVkYY4NA/g0MwzHW7JWj73JqwTCGKTKTyNEM4c5
wdioMBxAoC2KVfz5GIRlaDjPrT56tS4lkZGqrzIqfh5ds2NWYitI4qRuUw9VGU4ZSYLsmepCcGjQ
RC6BiXY6LlojyusQzzkFdXWAJP/rrKbKh8nqsw1Fvj5/zPAexoQ59zoOkoqc6Y0+WZQmm3EpomEW
vWeovE0wX1IVOjjfIge1o3g3srBvKuFbS/NncmE1luyG3LWXAs2dy5C3fivX0kIbTmRUdLIhmmY/
RgFiSPLuVAbr7S05vmxZEd6XTk4k0cfqsFvw2oIKcs4uNzDOni3f2WTr7dGRAw8RX7DZVWxGfBw5
EHLCXUwuCtWAdD1cIQQO4HLUpFs5Co6HvgrDJTo6wLj/8dPJFPFwimAnSrnBVAqILd0vdaLSkIee
qbAUBK2j6nkB8K1NB77R4Ylj14XaE2DoJvhJt2gpVugjWv2euoyb0sSZm9eN/ADPlmA0OqVAVTpi
vJgygThtZUXXWjgdxgXVnYlWU9yPJ2nV/zCzpMyje4CE8nElda6ePOd8zDHlKcOHUTbOtbZc9itE
so5YX++OVcKp/Yk9qp33ND2/+jyTAaj4h+y6oJz0riEni67qAyIpMi0it2X/vA3Ai3uyvxxLAbNc
fp19g/xH4f7mnxRFYvnjr0xVyUMMRlrao0UgYLUHg8E6wxjyr7VHkem/1Ui85qdpsr3l5zLQZ7//
ioxbshFHa0h1NWKP0EC/4aLU/AmqM7skwVNzd3CXVxXGHomIEnvc3EehHAb+WqL0WYiR8xzwViRI
HoPdfBLmVwh170BWWe9+rr1TJc0fl4hlA4Xp3vvK2mBaPUjdP+iH/KaIbKHLDW2tSOYoNoKGiEs8
3wYH8g0IUelJKUymPcM+CVb0gRyZ8P+bCLiAgP7pau3DXVDO5NmQmj3k5mKib1nLaJpx0x/jzf3w
xwqngsfPmKQdSLdl2R8l2k3FJaj9CfhBu6c94ITN4QGix3OLdX13wNfMoiEoYHZkxtQl0gH/GHN+
7SU2Pz7FZDFIcjkTQ8WrP173vzdztnuG0dAQnZbozLELzQ+qHLY+nI8H5Cv/vTyv5DBBZuclHdU4
D30qTBUd+N/HthxmbEQxTe5dG/MaTrBFf8Zu8eOE2W85aKBFXrB1BBnDhGARNtX9B6pdI2zXGwhX
Hy+oqLgvJUzSYp9kM+sSTZDSQt4+KCdjr8XgOMlWz6NDWwX0NHMt5TB1uuRFZ3xtPSDpW0Bg//NP
/iLoJaioSPBJ2kJtiDw68nXcBOsaIbSFK8LySt1fN2z3jn3hnj8PXmW0nEzoc+vhKSDquBNvyjfC
jBgncNW7WenloeMuCjf3h9ofUCBxEENRTTm4eYv0X/uhX5s8qypGBZxZIng4hfpbQoGR70j3cvbL
YpzaNfufCKiPs1OY+15NbBb6zc8BRNAwGIeuAkB+NYmCrqEfDUrA87dRybRkv+5EDQr33JF+lu9T
XFCgCLgSQlVitKDm4J0KO0v0pbstBd7Zi9+r3UHHe45Mi99YqhT/WOW4zRFreMtZmttxzdhMGhVp
qUe4dN/tU8rpxkSNd4jeE66aEjLtJDuxltwADk6Z6QQnLyskX9LWN2OG/RDOyCpLMmUldbivmeOj
RMqK11G7t+dmc+WT7fL7LG+4TEF8HcfBTvAF2iPFh8bC+pjacMr1WA1rhC9mw3I+7aA4Bk1KkfGf
D1jaVGhOyDFVuEJLN6f/jtSoJMJvLaxzTo7k7h6qY4KYFO3YbZ25qqKwvYWL9VGTTSsqVEpRRAkJ
szkZwAEZcy9LzFVFLTyiYEgWu6W25G2UfkCw1YI9Ioc3cGtT52Jq43rEr6XZPUSRZwG8Hxs4l8/z
R40xh0OQhOT3YXHYlSIN004ryvVDy21pkOpVVccYyDoBBC0/aD2VBJBROMIoadzvb5QFNKtUsuDd
lNE/zd8WvQNaJdiho2KAPHn2yHinWGSELW7QGHv5ZovAIBCRzsFVD2a17CyxtvcMyUgfNwvXUWp6
wP8VxOJJf/oIjnmzvAvxGO0NkKON0NmyJvfzZGiF3uNa7Os7WP3mA4KHQZMsuj5qG7Nv/MNuhzXB
pOrLlcGRJewRWJxIXAVnERBaPecqSooQpkdYBS7SrecxKsNowyENzG0ZIH000h+rwvq7GeFkjX+T
y6jOccOiZEyjwEG3xAjtEWzB783/RGhkxvHBSXZfPsgUusLwf9NZ6M0uIL3L3QtvdhrVf1NYWfi4
1fmtviYI4iKGKKCSHSBHWJrNf35vvo7JJ/SsVinB8L0O36zSeGXEa6MqHwv7RynPEls1JyUm5RFc
2VPeppMe4DnAsWoQHKBlyE3WIlME4um0+GrctEt0PJP7x1go+QF3MO5J2qum5U3vbR/cJHgwP1WA
SvROKO/qXehOCFGZglDd6YxNI9WRTRs+krYJbKD1n4mjEAbAosCbRUVzr+3mpfLlrOhIM5MBWoeC
pnkan7PbvyvFPsXh6Gbod1idD2YoEkTtTdrQM1qc50fr85ykTc5R+O/nrZaiB1GnyZu1ccR3BJld
dF9HpGmf5Tt4HnEDg9w30st7FSA6+GEpe7N6IFAO0hWb57HayXJ0ZpZwQoJC2WPsIizcgZl2k71n
rUjjck5lugV085f+zhNNAyG3XVlYxU80SrYUc50qVfoniqLz1/guwNOTge9rfAlgGB50ihQx/sVH
/m/mgUgg5E2wAyy86v0MvPz2uHVHLSmoTJN8XOpALu2yILj4FCqe7XXj6Mm3WF/+M/+ULy5IPO/u
BExR+yQyPA4UYDBwHwcrl5hoTzy03JAz+rO0b4PApQFxyWh6Il4A10Ef+Id7yIx6CiZcUzUwKVdu
VaCIIilCcCd1HTzEjERuIN9cqmri3dNfnLHDZ53DM97iqYb5wpwdMxYUC/Zl8bqw2CHJxGDLG5by
0Rg+TWtX051Y7nAJ7ZOS7d/Oo3Hvj3BVkHsCbGoswWkjETTCs/uwBLm2q1l7f4LmrT0N8Qc0hxUt
zZocJubsQSsxNOOPyozc5W4p2lun+bgWzrGlcZyKSNWpAp79bFiSCEuPuLNuJ8seD7xvb8WzCDQY
I8BzYqzVClf/LYRzg1KWYDyRAb2Sl35UGIOGgfnM03a7shSojCTzqz18cXDPjBY4uYr5bbzeOzLF
aq/RXvdhWf+R9YU1ZldTB0rE2hhBYdKiBsW3W5Obf7mtPChhVHweqn3aSW3qj9ZXDy1Ubyf25o04
YKBBk/jxqe9fUQ/d1bgjrsS5otzXhJ1p/C9TjEVR/WYgncL1+8eqDANfOVXB42su6KOfenK03tlQ
3fb0si5K5LFJpmH8I/HNZ99/K/cz3fXH469pXcDRST6G0INyMDZXkekBuNIvGty4lDIRpqjsglHq
gy3IK1EZ8snCwQC7sQABPliA++SL1k2oO1WKthtYArVTvp3C6+jpu4+QdL5WHf9jT5fAgzcy4UdZ
Jxnnn+tNC2egu+cqyfjdgVpJbeQMdzUA2Vu24/15yCu+DW+fDOCoiM3LnIg0Wz8BnHl1uIF+4Sx8
XfSR999ZTGJEr2oPsyCmd+wHKJy5vUbPUMZOWQzKMft7o3LEfkyZJl+Uafn+a9wplDfUvPrJETkR
UNr9viOITvqGdrBK5u2ZM3BFdw+gXcw1rm9Rjw/5Y2YTNCC/48PT1nU9uKQOsm1IkYaEbgRXmRgc
IhC+UHNsU3kyu0pfZiHBB9nz7iZ7VqWjNW2MKhBbGwNgkE1H6uV8j68oy4SbZ4l1TRfeuHIXROtx
budU8ErPD2TGV2Lm+4VQFJXuapfkDjonm7dbXn5/Y4dDC9KZf5HovelJvu/whUbn2py6c2DoBXEb
G8fEkgCKWgqCBePQGyzsneV6FeZdVFltHPYBnMNIiRVJW3RTNiQshU0e+Cgv1P4fNjuh0DCRiWqA
gybD+ekc9Lf3Roo7lHyKgBo3ZNnsuPKOOGAfpvmreZPPXwfNI2l0jG+ocsVxEkR3aV9oT9soGzxD
oZ1GACeckJh0dOxSY1V5jY9BBYkwHtL2vUS9b6LtVR+sCC6/p2SsEPtT+N++GAh+rOJYkbfvKy9I
C5fU60GS6D7TIbSjLD26N1Y6WoNfD1NAjDtYPuEEuGoAI/dkrWlEgZ4rGhHOqWI+j9NVRviTabFu
aINj4dy+eHfCN5WUnVj46duti/+sStEZ6HbQ09+5dSAM+7BMmygnmedy5SDWEhn7lGOBFZy1qYxZ
op6QFK5kPo0ZCKZ1RzaMML1o2JNLWFn3Ze80AKjfIW1mU+b31nHK/TCfskGEfdZE3Tv4fsirHIAG
ye9lYXhgEsALsvcRd/G71IlbTms6WWvyzQ2+9yHtLbEqe0bmIZqWnryDwkdpYNkJTlx1mWDY7UV/
c2V8Zgz+7hM47kThA1sfFdoZ/4TUU01S8m2KncaFMH4XieSxnwOS0cULh/qK+uSHCuT9UXUHC5PI
UY+CZ3AaUxuIkcSyQbiEwdQ6p5i/oZkNCDMkRJUliuE2q7c5FR7bMO439PtgZYKtiqnomHSbXSA4
KvQJ49cQLWkqXx262dXDKXrJDNoxrJdAT3qsGzMaNo3S61ZX45o6BA5b2x6jpUAGegr9kao1DdQi
ABg0or8U67my60yWVUSVhUqGcis/FtVB9W66fR4qHM4hKXxgSxjSbReDBcreXqdYE9Tb+XMnPngP
ieSarHUaSf0FWwh1r5ozG/JUQbBgoqpEmbLU6SBk74HDrjCr4P+K+wfFNfABZNANzjmOV6ZCnDS1
qrpdb8dr3B37OADDZoIEIED99CAL2y8pg83nL45JJjcixO+qez/fQZyCrHVfhYvVRCDZi9BwsM7X
y139gzCvXsoJenyoLoh62UVVXjUsfi0MAkb+iqPzoO38OUdsP0jaEXwG1Gjn1URJjwgPtzEoh97Q
MzltbZDpu5hI1VMBIai28c3/ZsjbHw7MnmgVQp88srZgN2B7sx8J41nUxs8PREIO3hTOooxW3s6S
EHIWVjHAiaKwF/z/aT5rQ/PFzfuK0CevO4U4x0WFy2oWGWDdEkrpgksXBWeHlpV7irt+5veKeC0u
QyiCzLAIGwb1FTzR0IV3XkZRgQdGEzFSTnA6JsWa1aa8dgxZg+pEkQyWH0JRM93ZmpDfzxZ98ta0
/xVoTwgvFtF5DWh6An2ZbuFSZw6/1pOBJt3J3TALLI0pK2TrNdnGQBZr7ldez10tJtiBLfLIE3pP
fimBaa7bqvbwG8W4I0abUvvke8A6dnAX7QD0gZwrundvlx4zdbax7If2tJi8LYjWd7/gXCHhNapk
V7bOVrHZUA+0AE2z6Wh+S5TTexYpwOsA6j4ZBHMjnoyf17qbo1RFY+77w1cnHBFJ4fYEyeQ6Bhah
ZxWxF20Y2pvOjiUl/V6v+nnMjfZLxIHIs5EOcyTM1DMj4FasLuzR+YM5TFmRnIOZSJ21+pztD7m8
1MeVcFzCi4iIup/saIC7p9vr8o8Yv2U5+C+ddO4Fk6HGy0tWwpwtOw/CZFIIsUUaFrNttpiLffyd
QuM9YVD0AKtSktltgLljSiDesJRKVmrfTdwg9J3gvIapwqQblsirhLm3INPf5G7jcSQ1T/eoLf5l
Uyt74Bz/jqmYQ0qWrfKGwvq5I7XEt3CZJfWIw3pnCNrCrmlx4bp0cm643UU+cv7q8BA9k7fjiX8P
H81Hd8sQcBELeQ9n4H/ZKXnqpJcYFI2uOGjtMykXwBxmau+gTtRLIz/92B6fnHkNotTfSyA7nCVB
zvCDCNsHjtFiGm4CxXXDzTwJ1MVVKpu3/UeTZDibzctaEQ8RZYUWU0HjbBX8oH1GAJsRkKKF9l44
jypJDY2L6ALwXp454zgBbXMjkjx7EWy+cE6Y4ViqbDywbZ3WOAqwm/lDUPfTRKKinTj0ZYGAN/py
cRk9wQwmKu860lfjJKE0qsucqzXQ6Nt45Sq4PkW7Xa0N7GBnGBMACUFI6GmUpqKAXzeuK1CTcP8N
aqkxhyj1ZknpeNeR4ygNiLpcZUyYR9bw4TF/t5mul8W8jg0AM4s3FW65BeUFwbxnyAmg4GqB36QR
gI/ElH1bD+Q3nZG6649wRPVxFtOwN6v2N8GZQF2qCIGtc8+SWn3F9Q3lvO9GwyqjEo+KaGCAOQT8
5HYKn05d8XXyWYj6b1PhVFhmcPkPLpVQwDs87KLEDmDj7t0gBLRwEndWD0GI4mpRnHw+vxX0UfWv
sFcHMqdGOmrDnGcxIa7Js3X2gR0X21/WFfIDU9OWs8hJoQrY2MzoxABs9Fzt9RpOH/Sewi7I26ux
bHd3Z9WpdNOZv7pXJb9swCG3FLdgIenv/vhciamsZWv5HbcNUf+3W4IMDr72XGBig64gX3arcx9F
QG8JynGXWo7Tk6g4CVbk5OHxqCqI15w45KHkudxZ1ieE22u/xmjUeoZueRFC0YSGsBYv5FDDux+Q
69AaOVBkluWIWPaH2hOyO592yTU1uEqJ8d9EyxL7NMPY1wGewi6NhqFbvo43Utskoh0mWZ19iUs0
ONaCcaJbMv2AHVnZKLmak/uZv0syvSFOpPx74ysGGzKuwYV+9J4BCk2eq/rP5ZkiRJ/QdX+IDADX
QaVQ5aEq1UGXHbn/BNHODta29R3xsumN2ae+G+6hHTc7uBfl1l4nyp8rz77I1uQRNG0bSHFw97kN
PoGH+2nsPeOyYA8MnUMcdI1mV+txd/UFC/bnmJAAfffhy/3O7QNpjCEW8wP4pWJ8EJ3ZGZogDu/D
L13HgTl5ULTNO7w2DDafmAFXlx4IMaRI/XPe3N+fBRkYyBqbsHJtcJwOGa86X+fZc4PYxsAKf4rp
rObwMXKbIc65yCeUc55+db5V+FoM2hXixdDhJr3onoA7CI6ZWefAzicurK7O+nNtKsm3ku9Tzmh5
RsiCYyToZ/zYRWlVtmWhbur63sHA8rZiXY2kXbX6RHHdngXoKtAshRRXhFs8tajoDwOLTuvquT8P
Mwdta7YPflNnUEQ3d0Uo8E1AbLFFfgahaTMz2S152jnD71qSmxteLf9r3TOfJLHgAGc0x40cwo+i
a+SKjla7R1tJze4tpRYDcC0uH2A6mybAv7NSRA9qzFVzT7g2LAeBeK1+xSdEIZ7dLbbcFsEajCZo
X1L61vtG6n8LA6DVJVBP7vWKvYETL9SRVo+rO0aOJFAzli43Lk2ll/h05ZPYELmZpjdDmAzIcZZ6
p9qSN3leia9spF8MZ/FKwkB6uWSOHOtFdYqvqCCsygV1Nk05XG5i4bpYyGhiR0BEks4M3bqXk/25
LzyyE4WvbrZmeN6MqjswlIqacixtxy2K2sM32m7u72v6EPiHyDsRc1I4lwAs63q4CfRjR3+cbVEz
iNSZvy2lV1xCCTKLAaWDMfmp4pFpaCESccCUe6F1EchEzazMAOWubdGLfhMXkf1nZlngyfmMRIWd
LD7sWEmyqPtSzeSxPsONcU1Yh41ZDKuXfFlMNvHax4r5Xh2RZxw//LdfCJJ48JEJ21If98fJ44RJ
apVBWAuiqYJrXpJa70ABUR7DWQwd+z5CZwAtt5FVgTD1G4084avncw3mBtseC7NQTZY67V2LiORY
D9q/W+5s0YP78keErKiPgvSqD4RSuXd5XIAbr+99u8T6gmSAYiBV+BabzKDb0RuhEDKte/TyCsip
5LctXWtsr6NvkwaRVfswFKdNdPhsDIK2gTM4o8c5SwSs9wa6aG99GqyG1Xdtz2ogFlEmItg5VZbK
ANS+kKP7FRh4TLG1ZtS81jr7mDrVMYQHVgpEjinS+j1NetAf1dLqMh92lsXv6AbwcOpF/gNxsiOT
0GGiW/vQKvwH7ueh3NBjrV8hM9MFYeXVc6aVltfcOIEYj/FZH/l0mCvQeaTST5wAZkTwXmCPxvNL
ZPxhKTOiak7tZmiSU/9X3/mH1S57HAdCAS3oFfuDmZokUaP23/tY1aB8ugXWOA5QOBSbS97GtFSi
DZzg1zJjGeB2rahhDfSar8w/tHgCn0Hgqfc7cVnWg8gpqBz2hDM6gOKJNqNmQKNlWyLbe69RNytN
PILEJRPuwPj1ZDlN/kwj9WM4caYsZu9RHZdAot8khRaJFh9871+re6exZ2tnOTyo8x0JDqGWfCl7
OTa1vecIm0vaY4125xAbFvc8seRvsZT9vIFYF+dlhyxrGSmkH4JXE8TMxUYlky1BzxSJb+0hBOms
HTkJ1FsLzdQAH75BNg1c5qPjKG/umMiJIfpSvzFfqtw/J+AkCZkZ+SVPcX4VARLo6eC6PLcx5+a6
0/pYE8XoZGTDXotheprgWRVvv7orYxQun8CIOA+OC+r3hIZCWwRIPpPR++JR8nhTWiccddSnCTO8
SBZWgX8gvWnbT+qf86jBYdaR8u9W+nKL+2VX0NTEa2p8V/94/a5DaPoZ87c/MLbqigh1KgY1+myd
yS8kBScl19PmuycTWd/24ICCKPQPJ9mcZXqDcPZuDgY0ws6lL74+bcQ5X/8L5mV0JjCftyRVbo5B
9Xc38Qkwdyy4sN2rtH9mja7fnWLVRG3MNJMbYD3/ILXmaQidg53fRFB8jZ7/IXCvEXssbZxqm+ht
vupo8+uasSgvdZuZuayzMUS+3waSVL7TXQCVL3er5iq5QXiFocnb+V5euaQWVnXAqBNDiY9xo39A
FXrr8WUB6Ln+LWiW/GvbqX7SD3URm5eBEJ1VZLebeV511CPKCxvtmZ0FWmdt/Zu5lQXbcLk8pnNi
9w70UGRBPHqVxoQt3U3PQCnYARHRmi5+f0Zd/8+0Q/uW7xljV5D7q33hVghZU0qPmZYWsb47zI1O
aIpljOGGEHb1XA7MNWeSaiz/nJyqp7Nst5crvacKqrgaGwOfqEE4rq+d5d2xBGWGBViTS68yOtWt
HR7gZi2FSDO/j4e+4T9zvHX5A5ILnYgLLdi9l32JC5o1i4F+4YeFiz8IvRI1D49HXi2OtMobYqDX
LCiHY8aDhk2fl7EGCMcQA8KyxPmfhwWciVWMaZjIHov+wCPHsekrgR+WvMAyjg1ugD87JfQP5X0k
1zqTaFlyZ/ZQP5NAmFUvSDkZ6LXoNqdyrJi7DMCIlfHYGgTF4YXIZTJN8n3m1hHCM4bSzyUAaUr0
KRqU+d7M+RwLK9hdODWd8Tb+CmIrf/bYiU9egOdVci71uygdCqiq2WGq8EgY9hiA1Ia05aLgigEc
G8nk1Qsc7x/4kH2t04TFR5sYAcmQjtY0xXA7wN9TDcF3e5h6a8w+seFoEeHSePtjUGpkAve14Tze
6V9xHzdItciXmnNchjWIN7GZWrjb458+O1PGECOJJXXISQKNtdtbANtNqPEQIdKoWf8NREgjVQko
Lxqsfg6Ebh9P/6fzk6LK4PNnZNdQ+gLi5QZLjOEZxV/DBu1jvu4kRjaXKCAIdvdwe8dGxHJekOZr
WjCJCU+yUrGGL3K/mQ6C7njMea5ilc00RjyhpbTxTzvr7qR19l5YXsRbEDP49wS09QOO/BGPuSSk
8aGHLW+ZEkcgd0KpzMkicpU+Ns/pSnTt0aHx3PkhHsEtw4/HAZrzdciTIuY90sm9aljxT2vTxARw
YqvQme2obU94VZaiIir+iU2MwU7aSeoJj0GChedunnwanQtijjys+f9qrgTgEb8nSJ40InA7jbzw
wsNLFwe6b5qBg3RrBx643ETB0jfdbQIlNmEWmPfYqlF0dG5fhugNfUyQbOC2e+BNw7C0LwXtgd46
PWtI5fPZQA+6vMQNA+QCliCYSEp1Iswg85PFUehBXBIZAXPR/hdmNy5C5TDukrdCAVp0Rl5TFGSp
/OczyD0tDNbib22NlwRpSkdh/TJyYS86rmb215aEV4xEZeXDxP8UPwZC5VIs6i6ne9apq1cRLIhy
i2qGTGWxMIUewoRe2xG6FI8kc1ItFwJzKZOHCyoC7IsT3kZk6oXZlzbhJt87mv1LKHoOtSIvQfNu
ga7qCB1gk+oubYlJKtEgSD8rw+8PaBUtRFL5o7Kj8rX4UeriO5EXlsxHkZCpYllqctit4h9wN4M9
jthN/WdXuzTCvPj0I1/NDAgtzKAT8V+Qws2yYKpf7XdG4D+Z8a7Q8Gj9EVaH8V8RlvLhhIvZV//b
LsTxh1rrKpYI5Uwb4a7aCHvhiBOVg8tN/sUUO1COUOB7u7Vky4bKM+VLKIXxh/2FF5/rz8FvJ+LS
VNJQY7R+lyaJbGajAjl3JlTyZdG6Cawada3A9ZdHdtH9MfAjbM4ONBqprdR1iYGWcnLzA/Wm0bWy
0l0YFqiSUIF9nkft60s87uf5kV7y9pvjfOeQ/WSbULD5oj5vAdSXhkaJCgN9fvNeu+ZPm8H8XCpu
Tb94GbbggmEXlgmTtNga/mWb7u82Au7/wnqGqjAtFfa2pNT6l8G5XVWfVGQ8IRRuYpfhn++pfh8t
hJdNtYxusYKfvtqj/JaUgv0PXmoltC9vNw5sp3dms7x/fQKOysN35N3+iombzlwJpLIB02kYwVnz
0WVaGi/oNqTBC+8uA0sX2jDWTDuDJe7qqDC7KiHbPQiPnQl74BX1xxzytQRpb97wO9y8+OlzyTEZ
LvzG5weXWl9qPacFZxqLDwfYSk1D1rASCsSHjmuuOU7xhQE4KNrMDWAuqrTAOPqcATvclG+y2Vb3
l4Jxj0pSd+DfqrxrBY1dhcCizM28KcqfRlyzmuWQbIBIRnKrb0yb3Zvl72U587J0WKSVUWVIrDEx
9AkMWzGhDzPn0XZnpEaq3yYlwqkwLsjeeW9B1q26vg251EnUtuy5lIjOp98G296JSN/z7UD1XPCW
lNzFY9MljYYAC0BD4cuxdzBTsyNsG4JptAuqhJuHBCXPWj6IyTuNerI7mW3SUYYl2ZZat4a2fXaW
6/7OkwW3NXP3PIBNTOP0tvEP+3LuOFT/sDQu3DsVkiFmq9uloMuWhAFgZ2Q+Q2XrrMEIi+9Z2Lo7
mVmUOL6RtlvBk1om4CL02VTM0Yrf0JI/6+pgHmJXR8FE6XMS8lVmgJUA9CzV9bkc2jaqvlTB7d+/
4IYAHpvQdC4XAvyK7n9xhp3R2IfpllbivoDYbsgZfTCuRIYUCTkqWthLbOJ9HwcI3gA6okXAcEcA
aVPZU2KOhi/ke1dzfawfq9WpVn1glEZmUfc6ctdAu5bxPlXop3idRldxSlzC+MLylLRY46NRsjoP
eYL9DC3p5xky4ifMpfrJq3QROHbw6MdUypKLrIQI/OsKiR4O4c4EQb4ZkeWLu38Aqm7mInV1XABr
Gk6h+9bx1mL3V0orjzUMQf5PaUPn2ol7Jog/QEEjLZ0HrrS+qK6CsVodLr+BrIKNb8ZKYVtNRp1X
UVYULnjRlj8+qeLfcdAsgfUXh5auDLG0Iwg6PFEo0yLE/PzqIdc7QTMjMjwlQrFg0OCqXzXBZnMr
iE5geJFHpsQB41JqqIWMzsaIQh0A2c8gjwUh5vh2aNBtIDLe0oNqEbHvDVQ8c0iDLl4cW4DgQ1gw
ebdSMYpGjz4bppTOeYSqq/oDqXPwP2mE/gEX1XCcal0eWC1UkG9md/DKbB2l9kRiDbNTKY3jiMFX
mU1oLZTmJ0PHjCpHWP23oMJIzNBNXQFWBNrAKYz62iH2evAYl0zk4T/K0JCIEnxC5lxJrXuo0uOM
3Rr0YVQK2O9VTiftEnS1L8we4nOhltTalr4EaP7i12GY2kqcWs4X+spzYLMXj0DbkYbhiXLLuRKJ
l4Pl3aN/nM49Xfam1g/aY61o9g+fn+h2oBnOhgflU7YIcuYsytYUiVJLa1+8cCN/4/JHQH6+QRlH
f5YcicunrR40i21Br5KG1VRYuC8jBPXcAMQVLMjYhpJJ1yeyNBx1QB/uLyiv96TrdohojNmg7ebS
oa+sGiOxiELevD3iNkdDzc39ixH/WtEQn5KZN5hArjYiPfJTrl0ccWAklz2Pz91NHzlzvw1+Aqnf
RpEuONqJXWbI7BSOFLqB2BqJdZiyeUTvG0Qcx/2LR+SE/vBcIILeasdzy3xIXTWDqk3ZXwySji8W
bM0kttUoEpnHynKimm+JRstvdS11oBSXELoc+/ou4cLUAWambm06SSOr8oGuSv9DxIbXFWYQj674
0uRSozeB+ZqijWdb5nICu+gwkV99MWnHBCeYrbyDC63M3cMjQOZotL48VElNBxIRhIDtwJj01SpJ
UbEx7gkKhyVvqycEFasjcLg/F+gRC8/kkbD1Eb+G7TVuMXZ/VdmXReXtsSAqoBLiGoI4d2xreQX2
ZBd5p5r4GIJKnOJ6OHCtVKDqHTDS+1Ge4gclAvbtSUVBinGoONAmqF3DSDV5QxHWUiAHQLKBX6T6
4inyUvEDJTNKIOneiE/r2cHaEW7+8SyqJvf6DDVUeVM0y24bC/KzRVuedF2nl/DhUO6CsCaxM6ZP
VCc6oNp4Z509XPZcplKTnYhvI3hjCSmcc90ZfgdPM+fxYQWvJvZbsc5HRjp8XX2ZSA1tZMOrCzkk
BOyTVncUSUT5UwhD+aVcsIafpmMTmjzqapgIOGYOwuI3PSU+g3dYx79KQUu21Ah46NSTmsRNETa1
UKwhVBGnC56KjjxTqSAEp68eyIMVHiimihXBjAUEiQJZHTHMPGUHjLQ4iC0jtY6V0bgLbHtKXkrf
AnG9ONjOacy9mWN6Be1gFmRP3Rfn083UZT01gVurL8H3dM5+nTHnNk/DAESm1Z2XewxdiW1jHi3b
qBwmbxrEcbQAYLBlZ4urNGg+0pq8ajt3HBnhhBciZST2ftMIzJYrwx7CsA2x9bVjPOVf6WrKP9Kd
w//u2ffonD8e1/jHBpjI2I2frYi9b6WWeXndRBT3xHGmSgLm3vukMRUl+fSl7fNKrflZH5+ToFD2
GOaxfG81phIlqaAz9Xvpe978qFhwq/rle5loAoU8J/82W9eMx29Li+jsS8xKViAPUSIi3BJWWZ6R
dK3Hmmv0xQuIFtzqudcZqx41IwwFG7akccQjhb5arfjBAfPtOjZus9I/J0bpE6qLS4QZ+fpRw7+v
n72qZJ6GKZ+Dmwo556hUa/XXmrRApSxMbTFbKpLXnysrno88Z6bXFoZpacAh0CACXxZwCDr3pG3Q
L0tIaGWM/jk5Oa1wqkiiABBATapRY6abm6p2ekuipC1YcWKQz3MCuftojUCkTPgChdmNtyXgPDf9
jy8Yjqun7PzPKP+IjDqcgchGps91Prr2Ue6SVosOMxf6qgWfbayiZ9w0416qa+HadZzFnsYtoGJ2
BrzE5VZ8CPzscuSxVtSMBpQ5b7NuW1aMD5QARQkp/8TFHSs0amTsxtOH5jZXimgb38m9KswTqoJp
rSsnvcxEBK++OZJC/6JFoYfqjhtRgOWYTNCjxUrEhCK7oCW4EaZcFD2PxCn7oCw3tM6KH8PMlCKf
YrlAQ10EGDoN3eOUxIHoD1guD50kYHYgikBfKR/2Q7WO77KhECIPiS1vZrFtjmGsSt0yLnOEDfvg
iCJ2bJoGI5OeaSaUBUvhuPa8gJ6gNaDyTUsIIpfdFKsWo2TxzdQFajQoPhPoliumlXnH6ISJ/Otd
l0whq7cAoWz2mEP6BEjQ1SNZA4qB5Yr99BDOTBHCHjNIdwtqEHlrMFlqKPnIfsq5xJroe4b9J3YC
JWDNlTPSaEtyI/IPx5Y/w/xGBWma9N2u9SLjzKWiSwXgFWlxAMb/8k4CTogMhkCzJn5zrkGomEnr
f60VB7KbFeoKiuOj6vJZpZwgOYcZh6flXVrDijeX13bPoBfMke192rIYg9gI0k/JigH7Gk+czEiO
Ps3osV5ffJDCmzvYzY/i5QMcsyMmYlSixr8yES484d3uC+ME4bFL15Refv5XnDb2JST6LO95YytM
OjAqA+CInAJpX1RJZkEgkjeBlZEQxSMW4YPKNVcSEE43g62uYb4286ElKu380X36UlkstmB5aafT
U7gLSUe4aNgzq78JjPs0E9yiq78yOnGfzIocKYeeoZoRgBvwwi/iepHgq6bRh6NoGyDIvp1OgnBA
NxY8fcoDwP0gaRjrTOIPly5R8aEjkCUVvkBGx55wYXFrr0CgJ+y5Onjo5zFeoOwWAzIoE536nR/d
pVVwaLNHapPVtKYyO0kfmlddk1cIJWDhFC4nIVFoMkcT7zukmmHFt4j7H0ZiPwt82BPijGOtv1Vb
7/mqBeRsnT/GcBCdUL+/lyIDziAO4JPoc2mwO9zMhRHkwSe6iQG2ooIuIxH0fQGDRumCrFnB5tAQ
jRE2YJjoSO0AF4OcgCLX8JjLUrG6EvgOesf0Xc9NUOPHq5JnHj2RZbRA1K+y6FqZUXpMUaUTysUz
sZBN5mqYXylYOvhcsbrgcUMZAdyZxnwLNOBJrUvoahQ2LklY/vLo3jlvU1ln0zppkaNkN51QTZBj
sjG0LmmXJgNpnLriQnswIMmXvUlpQbLTusRFL/Z5490brQxilEC2sOaBvEf5Wr4N9Uh0/rQfsRGp
X9jxaW60fmXDNUJPnvM4DvWDL/ls1Sc0oNNRPFm5j3DvoM580rhrx95Zt3Rq/PhW71nj+LXYxq9W
vhNaLI5OZbBKpxQeOM269Uv0cz8a8KWF0vXugppe+2DwApTvuTXrNkaMmqEAL+bS6oOuhF9dhNlb
XkhuDKGblzV6aWn5360bvE6w3biVlFJ1ORV3CL+JbyYFSrgX40TqpbE2LfLODGmqrL8ue+AR7AuF
nUS1wEUu0B9Qjo4cbmGiq+2tl9bWbvzm2O/asqefDfTvmQs61gcF3pzI0yOi0ReDJg0rHMiPll7m
Ex2DL5HjKAUxV3LPh76xfNtKY8e9Tz2OXXd5ckOMM+YjhZCE1Fng4REwR5W3vLOsdrxwMtuy1sYi
wVvW8lye7dg8Lo7Jcxot+0bam6SJapzaLYozRyfBnU8sbpGKqogipn6wtaZ/1KJ6i6eh8j+A60qt
gzpcu+XdvsGULJi3O1AP+nDnZXgp4iTgYBUItPimdzE4uIeVzfhSUkuopuDFJWykWWJGfhpz9zFt
nYabxxLQuaDu0/2K28OKJ0GyrBoc9lezKuSkF7QBQNf/GlPax3k66umRh4jNVoVsRkwbPx0gCX1/
YOZAlzlAZg6fEXnONQ0uLaENYiNXKZxERa4BGX6ebZHpZ4vjkgQcnS5VEhSjRd7FjfI4PrbYL76X
sWQ5+j60dP5E4cgyJoLkR789/T9C7+abMZVPqbxBTzghHv2cMGpIwunJc0hCOhvl2lcQ0FJMbRE6
Lwsl7bgnzMStRpmZuaQbBt9gNRAwCaBFMdzsWggqA7ltLhZRI1IipEWcNnxNgqIpCUrT1J3gdcvH
p308Dtj8P2+RhpaDTxiDb+HK9HaOGdmxjdrolvUaOy9B6IHeuvhK1km1vGflhZrF3le8VvRY5l0F
/lIR2ofZZWOO81uoSJt97EAG1RrqBwiQLJ+umaEZ2ox20Nu801ETYKPw+jqJtjpwh876ARaSQKCf
AwgBBW7CWdxlOFTk98ycYyvi6uzeWxMVaMbihFg+o+APf9zZ9U7N84xHTDUBEv4s/bQ99Pj5j/tt
EJOu1xwwr2pQmLep6vx5vu0FNZXzZP0QT1O+x0EAjiIJehBAcA291rjFH0qICEcA51CS8JxDikrV
X1rLJMKQZun94d7ZI7SouFzW95b1qRc2IpliolpH16bbnmNFKljjqcanvPAl4sjze7wSD1at/J5H
fzFGUAqswwrP7JXfcediG00mjePKh19xhzcHZMH5JM3GAz/achQPVqKcpj7DTZMzLEtg8RA4aBds
K58HD3kuZt5uS4A7i9h5CSrfzdCK1GZclzcF3m921RTXBLbJrWS4+JqHd6Vz3tDnIcE9/fct8Hgj
7wAqzIuaiFgQ5jIgZ1SjcXIsIVXjUQPe0HD5vm3B776q1jO6zcIaxN6onznp6SlrowCqky0+Hh9i
fj3YBOnWdpdQi8bnawNWiBL7ADhBBCxdr0g99PszyNKW38V3VO+DOScrMszVN8bMwPaDdCZp32JW
1IBJbCK6D8ufgUGZRSa0rtfEjKdu7FdOwds7BNvppntEDhPn3PqiHKuNyuj6WK5lC7t0VugLrTMm
VHqwumn05pAU8vGwf0aH4gTL0Y8KjpGIFKAGcEFShjW0vr6ZCs4MTA0o4md0PbgikH2XPyQJF3BR
CwXaF+s7mcr7Ldrj+VVls5pF4ITC9tXTeficxI2+TWgZ9s82ajEE2ar05Wx0MkSOJEEgmGf/u5e4
M+k41vgjB12TNyW2p1yAqvgb5t5ZZvniEbtw6y76p/d5zBpT/pex9/EZ/rFjfAZix5KERvTLebDo
FpTCAM8E4VHKmILugkGc95ZD7A4BKcguInhvoYaXVQz4iV+EpbCpc4KarOPLc4xDphXqfulMD2is
TZTOEnPU6o7mn0lwztttWry0jQpcG5rKwXvgBWHePL6+r/eeZkL73pfGiQwezot1UyCL8EywrCp9
bYks3Ao8+iXvGu49l6k4IUHHMiUf9SlJ1NIjzvMXarJjb30qPdrF0ZpolYdPYdHx+A0JEvPbAmof
XhXujdHA6Mq+pbD3eQ6c94sfvX59+OgykK55UBfh/DSa+IX5N3MyaAFOCg6e78crIMLwrie7j+Og
coSe/ufqJonBRjZQHLiDJJHZThRp9zJ1F11KWTjHS/c3SXc/OV6MbKS5m3V/2zaC7HR1rFlScwbO
7tz0rw4NFHvw9jh/6+IHXMabbUDZcVdPqZi1ZfEfv2il/oYbMbYriiXFLyN+C9tzmRPZZHxg4YtF
/OHW3BSz+ikkybdE3iNtKfiu0FAroYrXdm/FZ4Qzq/0jLqoQFJd6nrPrMwuelobBC1Yq9UbeLJAW
sghVIFdFNLnzL4XZGElKCOnD8JZSkgHi02NgvMs+CP9FrHgiT8vkgokaHZYNwowZ1cm1acdbjgVw
wUUBrFSHaCoM4nl/UyL/bAf/EEO7jxxgI4xgG+PT8V+y6FvEEguGq3+ZPHIvMew+WmYvI6tLoHCl
dkQWEi0aBAo9apRmSQOTTRZfhcZInpKhVhsf3yCLnq1FFh0lVY5/OaOTTr1hDO2L3nUt3AoNZN74
e+tIfKu9yS97qOPFeupGxb3lXcq0027Mk++4SUv04U/xb5YK6fOQsiq6VWTHnH9hFSpBdApoGy32
afGk7h8Digv0vN0SgzRAHiFAWyZwQUeiyCwd5PgzzJcdU/RE6e7WyU0RUWsx07V9pDeagMgAETIy
HhqUfVtX12hhn6HFwHD4Cq95u7/52bV3hwEW4otT1Lx5jUpXMY5rqs9JyDiiz/nm57X8MnLQFjya
ooyX4m76h6aSJzhhFDYwsCjIGoVr43d9C6f/UKlq6QQdOoOMPDQZWBYXSNW9LWbRHA7pg240xJGv
q7eB71vB5mQyWazVMAwNh3XuwxVGlzqGnX92TE6qyHiJ/qYSIqKUYbPHVZKYzjpRI0LPUGxtKW56
DhzjrZDZV3YM1Dn5r4P8s1i9Pb9Nmjj5kkbwzhtKfUlmSSEkZ21oJy/i03orYQQrH1/k2eOLWoX3
jbanohkBn9TzkjuNlq7C3iLa3gBQvxRKJgm//RGF7s9Vjjcq6BVsCYqigp/uB12oy3kOsPqs1xwa
3r0bdXln+qYah3q26St+4yTJGtAFf1maPk3WnCoe0d9NlTEPx4d6xwgFbmIaMdgdzVJ7a+SYYwAU
c4B8w4PhZW9B9DUFuQAgXI45XUfY+zx4a51r7ukBNQFAsmjNScRnvUAykB0dM2r8Z8VOrATiFZMw
l/eXs6uN1r7Mm9JE5vt5FJBQ1abgpzFjqT0b4/uk1fQ+VJC39Gtu5ggKrjM8zSIH5eiejcfHvqOf
35xCZBzLXgnDx+jCXCYmJ71RB6wDbdiNB3h94DAOek5MnVF2YC556vtdRYF8TdGpCYJriB6+86Eu
KhL0+2e6gbwYcrsh9Q8n7bjWlSGUHvOAPoO9nJGWAd3Ks0AqNORvMNOMbEgMw4n1eJTUsbfa1VW9
pXoQ9Bt/Ime8PASCuCDoP6WUsMH4+9X55Ju3A+jbO7XfDCoDFBn0fMV2w9uLeqXVSIsAkkcAzaK6
0Q76sBjfitC6zWWFn40I+ui/Pllh4uI7YVinpUDlapKjIL5RSlh6haio9jIE+D6lH4+6ckdaSN2p
FeHbh6UMM3S27OQrdbTFCgs0N83sMScjGoeuqfwmbEd6rDO6Kouw+qBGHoNbuF7pG76dgtdRph/i
g/nMhPRu/vEmTTR8Qn75ZggkJGx7bcsamNri2nYrCZ+gomTMagHs+s20t5E2ZfF0wYhzhuRxEbqB
03Inlthqwg0CTaP0I25h1QDOTz06mEBpOd75Zxws9H9vChuwgtq2AXHNOCWdXAXiB4NApZKiAzcs
eJdOWmnsa6LEPFlqaK1HqGW1JhGCJz5xuRJTISxM/hVpAbYYbh1UjTvZ0JdAzWSKHH7RPa9JngzJ
PSwpNwCxYVN3gz+wltQbSf4nu7ayVR4i8PQyz6xoDPg9WKXId6SqdFHrRyjQSgvCJ8u6STz17uA7
L5IFXSsZl4/gn7zzLbPk1B5fFQ2uFxriLgMThhWJgmMBn+HIIjjtubk6P3U5cLUeb6WLFFUgBj1m
tCcCpeKYbDLQnT+xJgrAJhT7teTVhZdlxsXRQ2B9d6VGqqHRPPFBlp6S1NYNEDwrjrCwMp6QK5Dw
0WQG9ovTcVkCtfKmc4ROEcl7z0cEGrSt6qAeBJhAHPnUuYsNB46ijR3O7hI31B0sVzqKdD/e8sWy
GgTok3v81zH9wo7elMA3+B3hOQAY9EYxgP77qhszId0MIWgfp7Y9zePlMeN5PKRGvwXzx793R1aF
0tobqOlf4+zsGRyWsA9k6hU8Bw536UI6eEofGmMxcI0uL2gke+h4FWbEz0jNa98DK5dofq0C46wF
N3ko8m6ic/hrKIe3hG0UU6PjXdcGx/iZC2uBqgNwr1TN8pJkOUJmUsgf4usoxzQbG6x6olMdQntA
0EKnzzzuELmgy4SA1W0Fo+07v+D+lbZMBl6nPMWuVK3ufpjDI3BOVLDQu1ykDyhyu+AiH4WZG2l1
gGiZsM+UZ/twhIB2UPVIznUshzIwqS4RdUlnAbr9smqCrGcnTCrn7ucVfDWv7PzvVsy6wZGrwANo
wA00d8298L2oaIypR9bqpKHgVBhaCtp4qXDPdm++zdHum8Zqcg+NYSUv8ShshmlTS/GlHd+n8+zp
v92vRT9VUUCnDLG+1n+s6h5cHjdqE0dw1EsKifrgZFUOAQ23L5wea23rCzyPf/KFpCBnjj93IL7c
d79wQwKvjXoKvihLxi9kBVCf6+rh0hCFafNyYJWdmsWIqgcXdwuOMrxC0hq//QagZRKU+yBz4oQ1
6itWMCi7e8PFFkGWBDol8jBGyLe9hguQLTGhxMEXJoc6pD9CkcBnTCm+GQ79Qg8X0v9M/WA4K/KI
+ocNkXgNHOQjvDHXSdr3hzABJR7CxSlNtcBSNeIC3tGvzzsQ78QhuZoxM8KVQ90H+bepQrwIWu7L
GysL4BhEICP6DEFrtmC+O8pW/sHmdKdFMRLtMCHW37Va4nsQT/3nBUXhkvzZEoYy+DVYYAobVLhG
Omybd+EbHPR3uFnto2PN/84hxToEZwrPruU3KkbarDn49Q82xy0MNItMv5fSINxMR2xi+/15rFxE
e4iRM2FLz16tQKRpsjkUg4LpFY7bocyaXuAJD98gjL5zNeEMuq34WYsL6OE/4ivdqWJGl7mhdfxP
PqGJsyS2Bvpalq9MJK5iiMa+J1FpQOrchaonE0L/LMSd5maeaBg0V0zniF4mjaMZ6r3nR0ziUaaD
Z5RzVHscNxoZdG75jZcXeRNsIbG5TGcN5uu8ZWhGuywn14528gAlbychWSyAJixVNI1OvsPgDpa+
Ft/I4NU95MjGdrHfyyTKXT+x/JEmRWDG6NY00MDay6n/j+7589wiVDWXKmb0gBlppwsxXEisZEPs
n9UqIdutvzW6ovMwS+oqCnRSDuJZ6D9CxCRXRTzqpTecyvvpq6Rg5CBIbwhXmL7ZJynm/zzFOX8X
M7WsoB5dtcp6rYgqxjXk9sV1PscIHPn0zLSnjYO5u5Y44EqO21YXbLeMeDa6lp7sfcM2oiHVMRWq
Ngd9EcmQxZ6RgfDSjsp0l9V5D7B1q4Z0civlcSNUngCOCBlOA15QbCjN6MEqqw/lZhbjQ1rmmjDF
fdFYz/d1zevlTKBvKW5qo9kwjjABbUDhP2eAVJwFpPVW7URWDYlbNp+7Q6sU+FW0dBpS2m2Yd5tx
ENPK4EIU31sr+gAlBgcdMJJbC8+2e+zLFtCyiI3mgCLF5m1Tra0nMUehF4vyRpQeSi5S3icPy6Q2
AeF9OjwcAntHEtv6WNOXzFnH4/5DCTAPnBrGJ5SKj0WFcOYtAJSCYfGOwnqF/sHNQ9OrCRndfSQF
3c0ljczOyliQDIjJm+5WQVVEfsH7CsGAeLj19P3uZlYc/1xhYrnSjvEbi05vTEkLHOJ1m7qZyUi6
nTAF+R72PDreS7mI6w4KyCCaVTGfiMm29gEyd/u/iK49kAxr4hjMtxBABcFgkTBQXJ+7MZzdD6ss
sCtgy8Y/C0zG49KrpzDXfM8rN3tyw0DoQwLNYuLJcn45O/iaQaaed0K7NOk7maiF8G2+PybFOWoh
06UfyyYhu6ACW+wR5D1H6hxJrZGdIKqk8/3F4oarp+z/ITjsYLepRJM8eflWa7l/cMOcUVYko/rT
iBkGYgteRprtHku1/MM/3uLX5u2O/1mrOLJvDVIt54U4wDUX9niMSGuSdRMWLWVo3pgxeVTzdvD4
ZQtiFizGp5QnH0I/TE3ExlcoSvCi3arb0jisE85HYlEZ5TcFTrRdVBl44l8K2XmuZEI8bfr6b41V
mNjWDdlbF+LQ1NPC7jsggvIr4YkdpdcElORTbOXjgiTSCxXh/hX2HpT3pZWwK7rKYwZjoUV/ojFJ
/WXRefwDlD+wfGvevTy0ONekzGM/T97XJft4CRNy5PJHXpT4mmv3cv7pv91QS3rEvgDJzn0fDhHc
B60saKXUsBzVSBMsGXlCeeq41vofyFYGNJjQqTxnAk5gdArvUokf8IDQ4LGkAhgRKj6jnq6WAZOG
i5P88ZdLOPGsrIfSVQ6zUNT/dEFuBR8mFXt+2JulEvurNDpU0kcKB3GHczbcswjGTA2/K0T9UrTq
ihAicwE70/X1rgY5SpJmtU0u9pAnmMIdRJnO2yyuzOxZKy7kRhNgoc/nuRtgc8wC4KfXPRxZ8EEu
LYWByLzwn4Zgl9807otLbTm9sNMc0xoUNFqZ/eZLRLd+V5SwCSxHSJk2soY3eeRfR7ie9iGmzF3D
gdrweoNQxSN9ixhxpR3QNe+w+f6fFkPRA6+A0eaRE7EK2a2eDeoBrM7ZtXZSTD4QEub03nrJAXJB
Fi/P884k4LdzfLhL3THsXAZAUe376jqrD3JBbKBbJ+KyNTn/V5mW+PDsNlfDihHCPN+h+TmaYrLn
e6gLFVwtJhwLVXYqKv/Gbp3YiNqLZwR9M1HO0SmSgNtlf4KDB4cnmSLMH9kLE0n8DKJnB26cdzUN
yiMuDEsQYJN6sq156YgOxc6MFhD2e1ileNAiXXWc689Anmx/eDE+jrr/soHpJH85OFIX6p6dO8vH
Urt4O7S8UmubfRtZJSpjOmwMY8692pOKktF/obE26H5vewa9Qd57HdZOwKynM2PsvbixNleg7nm7
4Aju7IXMkzWpQvYFKQvF39ko2BrNgz2rlhg7JYOqn7KXjIJ3nujenPP2LrGaPf0fdKHnTjNADoTG
nG9mdVx9HkdaF1fYvdkuuw1TMQUpv0pvha54UAivd0S7iTxnFjmFQJSAXAnis3db6j/tjB6JcQWZ
nwjvt/JGBtZip7XBkSgh0XZu6gi9Rchuj8wPqmcPgstiMuqdXnAOFc71ONc76XuG3wRACgIyCfsF
IhTuPeBGT0mOn1T1W+WFumaVVoYuiPRM3XymWMOltQW1Bj7H6JEMNIjc/abPWnsEH6m1G2YiNBAw
Bd83hd+E3zASgXWIOJUeavLZrfjSmxgW1+BBAHnFWQrlWeTwyXq+cAa8mHDZTA1TArDRHp8PvPeX
ihokwgpz7WUbJXjAthVwYAiVCM4aJvpCjX0a40unuFS977kmPhhqaW977K/ASfK/sNjmIVyuHSFc
vnF/hbjiV3ncJUTzMulFIbz93yeCr1G34WtgGHZlwZxXlzePXw7avUb8iJbESbi4xA65jpKIWasj
9ZBor8hLhgJrJUuvzpfJr5rMCrUVTvOgYUvEa8nmDo0bZv1qJ6PqpAXLYizEZEMdvpUxzUd37q5j
XNljgfqgDveFXdw3+QnXYZ2gsYlnpsOyNWSI+LtoXwJS2HNDKQuWxNlp1642DSDTpw6fu2nz9XlG
Rj0h/0WeXuGCQD0MF4hQ7H4O4YD0oUFUeIGvL8n1+UbOM8QFDRjdJRipH7Ij9L4Ka+bLYvWx/cOB
PhzHh8bs0I+lBaegwiCNVtNHMiYThNvWCeDFZQcqMc3BFoOX70OkV6nD2R7Foa71IbAJXO+nBR33
/Iwmlul0UjE8m0TChHE3XwDf9BkBv6bpwyQxyg+ISNP3ToETXDzt4RzGVwRnq4jNkADXwwNHuNFn
7EnKYe1brhe4LaSc4aIjBsDZEcW69x/ZSuWMyRfXOXz/tQjgv8sC0A9poYMkKv62G/z1rbhdTBX7
7wWmgvBchnMM2OcJ597sk3ZezP5X1fWiCMwiGmgMoYlaIhzvPNFggoIzN23HwQtTxmcrPrA+EOcG
7Bx7FdVRMfE5KG9DfGS+HOi79GBecLa/q/JGmddeDNYWvzEVz6fnIRLLYhQwqwOsnWXabmKwtcH7
maCuV3HDqqAnXtSu4HZUBhcI0vDtJF9ADh47lqHCzL3LMVe4r3sIfdn09+71ByXtgltyANQOxsiE
InOPtGzsHV5NVGY2cXcFSs6MsqQ1vIO6sLosFEycSbJeojOECoBQZtSxGcmWN9paA4sgGDpZYONn
Q5BIGBcUHUJoo4tSzHPlJyVzOdBYlW73enyLXM2Zwd3R84ntTIw/zv6gLdlNR8Y1fs7yWjp7YjAP
vRo2NAncpch+Bg34UYimg9u+Vl0h2cX0dtL+9fNEhgPeacqtZeXtIp2uunvtYn7P3nvaoYcU479V
VpgV1QFGjzU5YJqdEAZjO1bsZIq1jF8oD2sOEf3N3pWb5eWvLWzfqyGF3o6vd8LrPUUEL1psU2i2
iM1jm9MR7ULZHTZB9SP6lG7HvPgqjUNPKv7c++4hZkLd/Zy7peiSxifofP7hprTRveSNsyEV4rvO
WT5mkGAmf2Ydk9u7C2TLKIDsmqEOh3TXPxTReGSS70R9+5RNthT07sMjw4NZt1pmHXaOE+PHbkzq
MerOyAq7KfJQY7qQIf+M/F53QkbAuE138CHfK3OTYeDHQ7ow0RVB+dhRTAtmYPLx1kwBMlpxzYKF
kibg5u743wE1JXO3UyJWnTeyGCTAR46IUaFqILH95JZiBGDNoIdI32gguKGKMRuoMgA8ajegRWrU
D14MDNoq3B3FSNDuzJwzgr1oRf9HfGxVtQl8wlSn//SpjcQuW7FGG0kgc+cpmgOF4v8FEnAHZkKv
IZa8S/VcY0gzv6a7yaNdVfxDERItE6CovQHoTgHmUtIqa04Zq2WElR7bMszpKZ56npxb2/XKfKLd
4J0aZIsrjnwswvcFJvsVGmBu2WxUYseaP167xJNeX8vy6LB5WBrTMjN2jl4uZwZJsIjTD2aJFOEM
mJqgYxmDWftwUYpmWjTRijPSLL9sF7TLps9Jq7+aP2NJPQVT4TCrVhL4yAbJ22YCKkKp+ImWxzZw
rWNx5EYz+ZnaVUMvhvGkKoGkhmde1cYzG6Su/6wc3/tu+yy7D01GZBOVws667dhlTr/6hPQnx/Gh
jzxWGIltYD5xoMZdenASTTZuoCEPOrp6zDnxzbaefrHGf5SJD9A1mmD5LMO6RhuUA7nEfpA1Eo95
z5NtHmYoK36Zv6x+xQ81DxafEzwyLbjJDffbRBg2yZb+OUdc3La9y4XxioFBsdkre63rAFxqltjV
hzLVscZIt9qfZ0vYWRCI5v9DPD7ilsiGj+H4ECwZsRaKM6KZZG03JWWJMXRqOK4S0L2vRdLoMudJ
K/AHfdIVROb0vretMz7Zj04yki1mxpIQxJ3RUfOLwo+w429gfKSWKX+1AzsIabp71YqHcf+uDgnE
8dUHc2sPvcDkjm0cJdrYd4tNgJAkvh86e5OjMa1Fl/Y8hFd3CxAYwDS8TRJpLstIp07eDThGWQOt
n3gAb0eAptg7XrFUMvqwIJXghPX5z7z69Sn4Okh3UwUsmJSf0iAw2Jd1FZhGtfCjS0VKFsQA6St8
NUp0hNhgAd3fclAEDf/2uN5j4w1h1qRB3jsu/SsTwS2voxr9WKtj9/OlB4THK88adUQ9K3wRZHtk
+EC6lXB7mKeAweMz2pAZkh5cYWHhHPapAcKqhTok5E6HPG5e1bzum02brrq2Hxeh3qPY1Jgne7ZU
fuc66Tdx0XdUCtmU/mExkrI9YxzCag2B8BdbUEyqPkyc5YVulkzxOIL/1tO5x8GXCxhfysdg0um7
aTx2wXYe5iK1bqLa1iE+sk3/Njy8+ARuacwm16o02BFIuw4O6DbFpcJkbxfD0puWXgE08LZaDa08
CtY9eXQBQush9kv4gAGiXj43X2Zl0XWD0mVMzmCUdLu773A7REdQkRPgUYPGLVXe/G9VoHXGr1wS
bSuFmYRduOTA9iK2jXn+87vbOJ5s9k3eM2yjr+cVqMFqfUKJIQ6omZ1/tHiZnwUy/GJhHBIXyvBZ
bHAHaZjsQUFkI3rHHUJh/7suWOEj1D6jw08fk1bkBAZ4Ys4/vcVnJAIOKyevEfQ0kxGEowxi4myc
iilIBvK89ABs4MDnpumBKLFpmQ0jadC9WfJimyugtOvKb0jNnkbMQxZZQsbIZVdM+GZbVKpQ9aIW
gdb9utG47tKe4nX8UknVQ0Nt3DPjUkAv4ntfA/Yad1zFaSlh2bO8FQRLdQKr86FZThYZfjrbC102
Nae6hsQNEQWV4lc6lJXs7hEHoUkL7RmTzOdlXXpiORchm1VGavRKl7/UWM7pnI31O/syQZ78/VLw
ku1nXQ4vAI9W/J7slPCh41wIDiamsluZ4aVGwvoR9D3WrDtsMgpphX6s1pignoUs8xWnm2ZE6sez
E9FLwVTRN/PnDWKDI5fasEwiWLud4WCblPDbhSmhu85NUHKiyNJZ5TuAFIj06C69ygPB9sEp+z72
I3Jz4TvPAtHHB02a0NmxVKiYsY2GTHOwY2eHNvHuINdKdngc1nzv2rrEwM3Run+5NzlfKQ8TZwVa
U0xnZDA14RsbApx0qYrRzCUQon4bqBij0dOnumyVoDYGXiJZOgTvK0aUvT2Ob7mFMUUVmRbwFQzs
Pvtve+L9x+h1yoi1IMlZk0fw/dJ1BCdZX8ZfP5h+tVxdQ99aORkfwGAvYdxBXDRcpT9eI/fIhUCV
awtDMC+7P0E4IIitSYvmsb9u9uKWd5C631xprnb94bJ87EFYmQYucjOETNTBXSpm0iLZEZxe7JGb
cvnl0ijxb1N7fgDjNXFSdWhe+OlwzaCN9c8ZAaFXPRvr0z/l5D1oV2xaX2+ezkUXl0zjE3XlTqJr
okC/Gw7PfvqfkAX4eRKqzMGX5RUHz6NGc0/M7ffeOXRsUNCp7j4O8MbD60wPTO8NHBgGEjPx29yj
IW8wpUYTY3PrMzClv0tuC6ivspSjhOcJNAUMkPqv/3GPrIknZAg1Plc5Z6hfQ9YAjkfCqx6xExGY
C87+zvU20VkPh+4Ao5jsJBzsel4WnhQ+far7pmOAX5diya1SZBuTgquIJNeD4KBqKzeS1LSN8vO0
RNomlFuz/My/+16mSalzOq6nB8Qx9NcR6/EmuGKAnDEM/exCNoXwP2wEUvpkDOWzLzn/lGP8o1TN
Kl7Z5apK8n5Kk8ziFbraGlL3n/lX5G6vYkte+IdXuxIxgo92bRp19hfyYe7e7yiwYCcu6vS14WR7
UBQHClo9zzezvfd7GU4kCXRsdngiPBju2VujhhVAVOkNPbKNyMTyz7wpIqWCA/uVOhnsr98Z/C4r
elEG1F9OHyV4birSMxEdqzvYCwT3TjwB/228BL2E3osBeWctLo+gDRWSI1hC+ineyj+GsyjyPkn4
ZORJJHsFUEyz+DdbdO/GWmLTNcix3PnHJIFyPUcGzk/U2tnIGJ6iLT/HRMvSHooPiyTn94KoL0US
+ND5OYlNjvuNQNZR+uOC7PjRRdr7mCIQAetPz/KFYem4sYeN424TWqJt9lAblnmdjuTTLsPzLCPa
spSdC9AtKNWkbh2NbWOhMUfmeOKIveo2U3LMC7QCeoJX1a5AMVnasxCMXHjXzuIJI/+BAI+dR4dG
iS9seMgqZwk+5Hf6zVzyv3lm9C6uPwVkuXphB+bt6DvGJ1J4g2/X+7f553WiArOw1uZEkKoTr62r
U00ZXExrlRnqasFve+ZXuDZYFOVSAI7fjCWYavH33e8u+kA8ibsTbUangcNx7EadI9vqZD7s+UnR
y0mYgN6/Wyt27E4FmCgNWQcTsFtEwWvwNhtgT4LmIA/r8o1zTKMP/s3DivtlsCr78yHCNVuDsxV/
uzGk48lUwBGmsn7WlY8ISgFuPKEUPkBY5nyw8vsyyXbPF/bxOmkWTQNuly1VjZwul2qPgXq2SZHJ
Gij/N7m5ZIF6+CzTiUgMZeMXPmoNo7wcmBYem+Ve3XzbBmxcfK8er3hP/5HXAucf4AC4op3YF/gK
Gs3ZJjK/hol/Yd7FDoSzIX6WuJj3N0X+QM7E/yF15pmM1Edn34b6RSOE3YLFqbfW5FEHLMV2H4xC
GMhdUz9fHR0e3mUwI5wueWCRJLWd6p9Vxm6aD1Buy+XfLfhIVUa1ppRnzi4EgdwSQpHbxWf2cRAZ
AGycL6q9GCU34kxwxhFf7wpr54yjmoAL2muSCetKTOsId8uv0rowYt8fSkv87qbR5dD1GTJRMoua
bjamseKTK2mTTImtLWuSq0ZRV9G1t4UQdndPlApWr7K2Eiij0447Ct/3Um+S7vPfwYS5aJ8C9Bao
pREZwxIHUjySSv7Xyg/fBlqPDgJpvXkHJxMFsP8k+RXY7Po2Reo3iZj7XzXQr2QWKPDnV1o/EMKS
hUyn58ScNpabjRKdh8o0wgTbG0pmCPp6vcO7cPvSV8B/EOWkZt7FerAt94mrxXKFn6y73AWnjUJo
6ADMnWhpPl6k9BSOkGlfwUvkcQ+GosJqKysP4tROPEdQ9xE9tUsQL3Ch5w7Z4P6lIPIWTq9clctM
LYlZhiOlbCAGaZVAWKiv5WkDnvCAiYlJG8bcc3IzN+kcDJNCTD9SbpC1TkYiRJ5e91KpY6acLoVY
hQY6slFNsovqCOY4CYDTr0nC8lrQZq7mmjRl4SQ5zbjrGmWzTIFrP8n/YQOzB6/XBqXR1xFY6q+N
BiKP8uNRSU9zz0sQhXo+LO00WFz1HG9djm/pGCvHY++lXP3P/GrXk94YEg8up31+mU01JcNEwuet
lVSS4QTgp4+kVNuptRaNWpEfnUnw9VPQMDcL0lglsLGh1Fa+5odfs5kAsZgIeMPEl+DdDJPGXC4y
/HvgOghCF653lYGrUubc2s1Twkk+hLnv7MfPAKTTxDAxY7laJlBDBin1VoS4wYfMCIi4f5hotxsI
K+eH1qYhX/RSjDYfqKj5N78KRFeSkriLJRPXCJUHDF+GBb1/qczSYukLFfVOjzqX9EZ5JQY0nk3r
3zFzVW7pFMQPpXRr+nfF+e3nyYIVugBPsu6w2pEbDzwi+jOQ7/4o0PS1zEmuGDXmFBPq/l4pheb0
zBvq655m3Kuk7LA7dj3syQRt+zaisYa5hYMKRaiRuMHRS3caXO7nHQMIz1g4uiJwFoeXEs3bjUaM
h17qu7CgYgbD4t23Etpq7sSmZKgqsJh1oJBFYWq52LiZ8+GUKNoZ5K2/IFRCcyDdjvh3GxSsBHj2
IsMors/I3MV5p3FluoBZ6GhL8UT2ovpwg/sFGNg3EJb7X6Q3S3P9gsd2VMrgaskekF0adrvLXnzg
VOn4gmY5W3pcBxYep5jP/xjBIeqBhh+vOosD83rg123zWrjj9zYIzOEbMF75Yyo0VAOq91E+Bqih
oE5nQPpRdxPqOfhHa4VdOwktk0Aq1liS4Hhnc7zRQCdOs/hBb0aWHAUDD6dLSXdyO2MSAIIINE5b
0Co0uP4DcJDr5RfOFSJBKKPTJwdpE5ky5LU47KHgAaADRt60cLRjPFXyz5GwKJYD3TmAwZ/4bq9+
UE3ky6R5leJb3q13uB8iIHx6WEiPcoSdP94KXs/v+iGJ2eHFWJKN2HNuMLZX76lShLG4vnhHyD3h
04pF+mKNEeH3d6laxnEnN/LtLdjoiUUoEKnEJaThFcdVi1Uu8QaNNKtKWovxsOKLT1jVeKdhomD4
G14C+E5xSuee/hd3anpdes7mEa3va33qJVtXY3Tqm/l8fdlgurFR96PFz8pnOJIDDELADyAa4oJX
cY6Tb9Ic+n1rLYIhoPf2sBfkQz+nZDdCM2Ccq9hute6fav+oL4QSG2yF05dj6bVJy7uI+DctxI00
8WD+ypFHtKijPZWi+dhqbvjukTzyIx6mYcgJXH6aQ6hcTpxqQiLLDQubHCuRofOSeMemSD+9NxVx
avUnprPgBvpbsKztWJZgQzlGRXOdZv6ZtVCLr8QdOC2SRCoJXXdTCE/nxWFVu7crF4NGusReYXy3
WxzfzbfqaSkQcWufR6oCT0PB3lPvmLEj8s93AhoAythXf6GnDrA/x7+fW9FTu6uhRlniMKUyetBA
xwwWkwPe7VPRUusNM8d14v27y91G8dO7pb2XiiGDEBaHyq5PjBgN+8eLUVrMgbOoYuLyYWGCjBt9
noTzljwKWadNccKrcDrmkJWiE7U77CbJ5Cu8IZqG/XvvEAnuH6QDS7KLHE12cDUeoiLYAmhZzkiR
Fna0DCrqkt33JUN8gp7JYOdfCthss4doJR7BCiDRpKmZxKuimHj98rJiHBcg3bOUP00g2gqHHjUZ
gSy4mSryF1UvxNKTnlQVXlRYwQBG13mL4tjGHUHQ7yV6IhKmwowZ2fweGZIQXNLLk7RSvsJJ8/3u
nNdwdwnHAUYsFWa7TcgrOvxvNxga3CRdKO1EHfMO+wDi1WfPcCCtSLx+Hjm9LDMaeczSXAV11t27
u1QjIB9drcBE8z5ZbllUr4bFSDHnNgw4ZRHBRgXU1OYiJNy4oFsqUATlgxu/IE7XccFoRZAfxJ0u
wl4QlBI8+JaHKfFBZ7pIY9hieaHjPl5ohoJjw7q3Kj/oPLfiQzeu3etjCXjSvE5cMjKqHfiYiiGN
IR8kTxxJT7HXDtse2R+LXUUuNXOxmp5IgMyKgZhcQ4ybjvbnJrPfZjACwcfXMwrfQFcNlUgdU8ZY
1dBdoxCUvAIsDJkxMKWPi2XNwSPhhHGkTZl+oO5Cpukz9f0R261coUrdloTQQxZm2vPGG7zuC2WH
nt9kAZvm2kNBWC3olud3RP8bivlpalS/WqtsexXYY5RNk43QjbAIhpsBfnQVLpKBDq2RbhwB1ui2
VJdyn4AFkCgkepdhG07ka/7bywhigV9d1nLYyfVLHmt1iQji65Rnx1L3cFI7t1GeaDnLjF0A+ovK
SYCAvIDq9/XP/8dTECEqbPF2j3jTzyUPL+HVb6IClcIrDxwPsQfrD/s0FjTWwbtI1OplwCa78J0j
8L5HAnYJGsmssCMqlNN6Iv+DCQaNqHEfU6qYFEILDQE4WFFFI1ceg+MlXP96muKcjPa4j4JFVq3q
vZMeVft4k1kge8gRiGe5Kmli+kB4f5xXiNW9GD0lTKWYaGADjsK4WsN/XMMJ+hba8Lz0t68MsPlu
aGovXLZ7ADzqHoM3TEbaEORQAeIxKn7Gb7XCMIWX/Rz8yEr3NclhX7RrN99cZbHRqFl+hjJmFTNW
4lrq9GHZH/63AJkkvsYqzHczHICKCZRE8u4hvRj7IiIy03LOB1uqw4Ks5cIv4MCjz2ao8jtkwN+i
3Ih+hbFJJf+dpesxsjpusAwDwZCTw1i2yh8Xtu2wbVWl8QwbwdFn5EK6AuqhNVWRvYCjWmiI68lm
LYyonSeMQAOj4I0zd/fFkepAb+doy7oLfIOev5npr94OtfATBEGEZAMfwpwyHzJRhJMCETFateeG
lpyN41EKy/z1tsZaQMKWML71oCkHGiEGfVDkHM2VIo2Pm3p8e9JqyoKSAfmT7CoONH8e3iKpoUds
nWPFhHk8cCQQ+R9AXAznvKsE3dsM6SOy3Yd50UWgfXO3kBHfJas1ueyj5lYOGUJj6c7hg99zVy1B
M4Gn7SYClx+w/M5cnYH6tap/VCgQMmzeF/IOSsMVekggkBr6oQtw3qk4EX3HiCmGCpdbJMhz4isZ
N9cefaEADyBKWjwyuLGntfTNA7UbIFNd3So3KAkG2o4V1Z8r9G3gzG2oFZMikNZo4kQ0Vm7z4xdP
GWiNcv8HBnirI0V5jNm2Ahej9zzq/7lRAG9N7UNMj7N3HS4+0ZxxXL6evCb58B8lbErnVFgFqFp+
8SI96vVwLRmadsrOWCOcwvcXFZssU5OAJDRPk77/zdDwYCsxbhBwnynCTJLGcH9lzY2iVdS6wCmB
Eie+6QyQRyVfOqY3oOzjJGSoGWOquZ1IKKWcVlx76/Bwjwhr/XhjQGYSUk8m7tA3bLmcKUtTKikK
Arx6sTxdmhOutVr6AXsGEGF1PeQ4wfu75bedlsyDpG1gnoejulZdA+reCz8VStjDB9DtQcIB4QFm
YSJ9r586pDJ6+cylexWb1zjysKoP4ooMp21zslMDxqXvAO4UlpwAV4e38HprUOh1SFi8Vg0xLMqD
0DC0i9Z+YmI0fTAnqCa79Cnont1i5PH7J+buW+zWbK0OwfA+7Dxj9MIj0oUI5nYcuaUAlcFVGGU5
4vDEllpMaBQPg/Yt+bns7OqzoZC/YypFXrDUkv5o4D533GXPbLl1GemY1H6xZi7SOOrpoKlic3EL
N9GbTDG3954GfImX96cJ6d+LhcwKfwp2+PacZgWmeSxi0Rt6V9R0rj0XnlPEA0cJ4lCt55r0dFNj
ksjlaYZhDDNA3RQ6EgN/tA+QUv9Uy8KGcSbC7K7LvOhZnEIy77Hb1mTjoecvVr+3zHqBKS8f0UVz
kf1W/DmTguhBtV3K/qFLIzU2TcwDO8TjXNnYcpnCG5lR2ypzZ/YyEenA1aRJmv3gwQS2rY8+xIP2
+gz0JB3bUrZrWllj4UQJHIK0PjYLUuTz7DDktlh2Gg2iUXe9FZ+gSsV5OvVQN1yseJPM4CImHuRA
5opdLMh2FNzAPDOzBlVqCEM59PCG2h2YFr53sCMBJnH+Boqqb09/A2sbNL3Z43QVPSo/7j8qZlsC
QmK1CGKaXH99XXNilHVI9b/HMpJF8FYLD97JBN/RZ7wqdWXAzNHLXK9zKQv9ZimdM31seG+02QvZ
/ljknQU1uAnCTNvEYqhu54KiSqhzkpQrX+s6YZLD59JmjmHvTQD8re+A7ZzHHGBAaqvQgxMH2M8j
R7ytSBgFGHdJt1O7CuBUpgcNYyvF+1o68E6SnMYU4lV8Iy13vyyIwBn61/VCcuydHc9nXEW/YmaW
mUMNWTC78mg56PtYrjtlCTuOiGNLHjEQvdSqWpsiWL6w67mGc4jLYZLav7QBXIH3Mok+nKNJb8BM
02WBIjKd8dRgG0X+HlROuR5fUf51qxOBxk0IZNwbB2XLT9c6RakbMu/sxQMgTjLx4FKFKY5RguHF
Fq/n0/LGcDnt3yhnzXpeuLPic/yERWTnJffpJIqQqBqywykTIwEQiq4Nr8lEJ+Z+AqG+usJblclu
daHFCUoPWMXVinVACe5UYi9we4aVCcNNAaI4Mphr5Zf20VuUimDbQytXpgNOOjEAY2pn23ZMVQ1U
76MbGPfAR2YOSJNnZic1bEKSgck1Wsiq7Y0U4TlMV627vdGxvfdcgIc+qmcYZEU6tIuObBjnOkvE
iTMEk3qyPLupxSNrW3MkWnSqLCSa7qKnwYvZ4CwqPDfdCJm69ppEHmp8fgljZ7f0IQ0GlnGcWroD
W5Uw7HokacZH+AqC6xe8cynt3opU+QO7XcYWqpVvzGPPnuCP9Cgmkrj02P7f1hQmQ7M2VA9oJTfV
fx5xBygwKeLdeVhx2FOF6/0ew4UdjuiplBdEEQsXn8RU8l9ENYkcxrZNZGgNNNRgzBUQ4iyaA+5o
VMiyzvcnMTrD0YEE5KQoibMujRDsUWQgLht0uxq2diqEAiq4enew1agWS+vfI38kWV+843q0AxTJ
H+kTZkG+U2de2kcku+hd972h9imeRHFqctKY4X0uSIkGBgsfyIc401/v5z5pEJBtu+1s3mlZXMBv
CFIwx3g6gxqem0/uW0mfx7GW1/PcyrwHpyMcZ02dPoJvXRSCxRiI4JeLqv1f8lRJOjzbfQkpNEUP
Era6WHrpwgFVTIpjl5q3mYBqKXLZQf8tdp/xTFjHB0Ik2PZRrHqfeXLl6jz/JJ9R6S+SSuh4F59q
g/MA6hzohjS6nntcdFlX2eo+I1N9yZrya/KYxJ72xsYM4hHN2DJZHYkDMX1Vi5ZyR0Vu1YSRvKhh
iiDM/s8yZxR+mPkFoHGypOlPfWpfVMCOjUSAO+07Sa20Pt6zYxCzziHOnqcSoCojpgW4uIGCCP0E
XGbO6YNrioEBW4x8Wt5mFWNKiCcs0+VQ+0tk/W52lGEUWriX5/xyDDaZgGeCPaOjRGoS6LV4FLiM
ia2MmqcQenE5DFLH6w5KfrR/AOcNYdq4oHjf6lWDYzlRdehmqr/e+9zifQ0U82JV+jXVZc1+ev6/
i6jjrcc4qKonUhzN9RElz96L/vUpxLA1T0DAea7jkAD1F+/koN7kc1ehoriP2YlY3BSrNdgyua9D
gdA/CjcTxdJrvwAzuIclum+TwcPbCUAUo1uJpYIjqzJz+1L8k7+wIoveWcHnlv43ent1Ag1z/85f
+ns53ZBBR12se52I+g6pC90xQ0fdLZ3kHtQQUcSwqQFfPhNVSMmBLgp7unqZD/nQ+Vkw+ySLqo7z
XObc+cAbpq/9TOHO6QG7SgnkHCTGLEsipvUzh4mcGPb5zgSImOQpoNoiUT3dvAObaMUbtYd8GAGQ
tRYTd2ey2rEd7csX9syqZKou5duZyN3X1yDu9/LzbuFV/zV3DKhatZbq2RJ3N9dcLKkMyltj1lXC
uCa+njlOuFKXVVL94MoS7gzTcT6vcw7DwSjur1HSqbWoWHU6820/Em13OKyQ4yKneE2E9iV3ZeAB
gSASoxqhPmuruk/Zi9NJr0unqRUjgSg50TGOFgvy9V8OsoF09mh9akdLvks7Op+S/aNX6cLncDKX
nNiVPLL9uC3wXirHH9UJxoF6L2I98MXpARUgLqMBzw2+sZRWYdDGcorV3M0RYdjWEQFrq6A/JCOq
D/YTHPqdCm2m064vsamtVcYwRDJ/d6m9Qvr7CuUsZvrDvb7j2KFrYv0Oy9EDdbOwZA2iM9arJr6R
5/PvVwlKminJRGYBJYk0OnF6xA61z7Poma0g+aJ/m/7ikeVOaZRSEtGX3ReRiko7D3T2mQfw9E6F
IKq526aT9tsY5p7qpbvFXtvs/bYD5OcEWAjp5eFaRWdtQIkwlkTmXd59aRD41le29e8ykRZGeZzV
cgtc5Hx/uJ7rKwQ7KDfGtcIpMa0ztF0CG1x/KFIPASo6cbN7JjmrI77+6Ue2guKls3D4fPDvqecM
ndNNLQ4Zy3haiPkWdql8rSTvf66ZP9w2p9k0LezCghST0Ty4yZv0jcAwtI/GQrBtgDwz8WUSPGEm
lVd0YrClbuSDTjkl7eWH1/SIrFFvJ5qJ5h+QGcTFmnqVdOnrIhMJAQ+4kpraJOxWKHagVV9RDbaN
O77VBuNdz82CfuMAZ8IdZpPSXb4JmQv74PXqBFH7pfh9tAi29B2Wt956akMlspZQ65NddHeosqA/
lNz6fsNRC+qofXDZEyDFzPt1AYv32xYJjOUTa1LznGml6AErSAVRH7wyPOjZ8+0vqOCBEzaDmz08
S+V0uM3jpn1WbwvCOiXPdqx5DlC+kIy8+toPbgJC9heBjOFPtYW9RAyrucxijaAUVdSyi45fHzDG
bDvffy8qB4t67XPh49+HVqWLZQeKsLobzOdTV9sSo/g4Wh194Q+8WT+ovPDrmPKqmnMk/eKaVrVD
sgyxoqbrrPs+xitV4BQ0yXubiwgFYBXrmlhzP9T4LYvEJW+RNGXMvRmRx7lwBrva0EYB5WmiD/Jo
dYGSjGae9TGvn6ZKMw/0WTqpEzXhorRz8Eh2ukKuFgMV7plTxy29mRwqEjwl1mMeh1cxOc20YWcs
wzpy49VqkFpYalsp/J8dPU5o5b/4NnKhS4UoB8F+LCyqoOtFMrw4wdkvEeByY6cQ9Zsy0/ExIUwb
6fxwWex0NsTDcbcrp3NgbGZh4oNyr03C4V6cmx6myOUzzmWMAdlG3U6MUaEdqEmvdOSvzRPY20du
DCEXAm0/N1foGzxkejYvuOL00pgu+W4b5NuOMOHIpGQs/D+rHn3CLpfBvz24iFfN9Zs2lFMi6L2g
KdSWWej4GglgOHiqm9wzSGdggDi0NzbqtCH7BLx25s1j8KTCU+X6Fu/Ja031Zp9tq5XpeUr522Fk
sWI4ROnSCZ6uATcA5cjw6mSZ9RqBk4CZigZbCZCDk2S8sF0++DwBDmOlWW4yJLLf8ipkMPEZs0ri
afrjGNM51oDY/TVE+x3G/aQDmycswtJvBsozOR0YwIrVrIDZvuHf6ViAhK7gMmTwHkGNfxz+/5Fe
DTOObZ3iFcs3I84wwz5oqf7RgWu2oo3PvQzCV5+R5b051feufZr60dHvkX+IcmksmhcJeZwdfpHl
g0F9a7CY4L0XplhGKtdIiHNbGhGqDID9uIJ8kLfkktybTLwVSv6B9efHOJHv3+lP16b+HiOZ94MR
+tV9JZ6ORCiP91pfh/fGELoZNa3C2/CiqoZpgBS5/s5vY8m0vmtjlze/2J9KSvbzyAs2apX1JGzl
C1W/he5Z0m3VQGKYgFGZrTqY+WCMdNtTJG7izAf8LAYJ/TAfD4HB7jgg2jjOrMDviAZEozHMhRU3
tSjP+RsizHpGiQtpqBiqwpGNr8uZYGAMXmh6UfF3SfC4aO/Y5y+mUPZBOLjg1B42hufJ8u6P3SUa
lyJ/hEIh84u9PPs4/oz9JvoeC2mOZ9Ftxmh6xONWFG0v9AMU9SSDiYPDzbt+Y5HilhsEL/MspdhF
NxHFaoY7Q1zvU9nYWStPSLQ0nGCVSoTxFdIaMQcFXJbzVrFLprrKCStQv1wfawYmN7ucZL5WB0x7
c2etacbLrHzsY14hash9llSQrbMTZXu/k3shFO1jRrl8T8xRFxjJUVYw7VYPKqTr4iU7vr42gIHK
aEA9oZT+dl2RsafdEFXJOHMprPhYrfzom5U5mJZ2tIn4dznTdY5NFLiszeZqK95gSt8lrHiU2m4u
1ND3vnD/bvfmRh4zEqB/3yq4U6XOeKNK1VkERRtnc5qjWXAwVbMSTXEkELFLqDDcVNh7eS/sRZS1
WkAS3zgc4LmrmjlLr8ZZfRCxO3gaLB1/zRRa0ow/iurcWAnRjNmrHu+YFhQ0k+93SLSXI7KLKJGW
sW+NFLjDBL5wuCxJx0Qx5juRf+voqKTYStzClTOiyoQ7KxtjJRplFUNqs4PHKPK1LZagthvfD4iw
9SQIr9rCCQyFBQki+g/Lv3yDDrkFGFbq6OFYiaAwrdLE7mPO/IisZa0F1ldShzX0vREPHkb8aEFe
t2UNEGFp8xUE3DsBIPIGoKacazWZK12oDH5OAviWW+YlqO5HWeeglx3mD/M8saahiO2eyIWk2EMi
+GR9jIORBL8UldjJj90Lue7iFitJ1Bq6w2MgKGOudrN7+em07g1xB5ogQx2YS1em9nevkztUI9fs
Lk6Lb0D7fVfyFelryxmEsm2cdxkXrguiROiXN0pZyOCHf1x06NqaOETJp+1UFNvEy7KFO1FGHRxl
Qq9eGzsWs/Dzy9WqvOZzyJQDYIlEUS64h3hgXlhodZQcL8WrbaqomjQSHvaQ7A1h4Zu2gX32IXyd
IKLTjXUOyLARFFmBMeV1D7UqanjjvH5o2y3RUd4TowE+//XJj0QZCjBTqghwFHmLxvjIcRtL8yDi
i2jBtTM2feGaTHZk9RsBqY6257GzIr2wNBkgaiRBtKafGgsVMf9DPIsW+DFLsh3L+cpRV3d1OtE4
gj2aaP65tJmfDhtHJXJAO/+NCuPGNKp2MLxasoU46CnfaSMUQ7sQDG6m2n3UNUvkphvWszQ2PHmu
cQsbAzDtV44BdCeYhjP5F/yPVPvUr9+PlsrY6eSB+b3GMsZm8RGKvhF94UJMOJTXRVVtXjWoLWcV
rY4vcXiInC2uSZrVX63edYQNbZO8Bmcb8qOopNty1qWIO1eZezRi6oylG/ny8vAfm1R2IQWtMtWZ
trl+fz74sQ0BsiFHK/Ykn/r0KVCUTJidDtN4IeT5JWgvcviGt/quK97Xanvs5ilJ7r6iFeEvPxrK
GXg8bG7NlIgB5Eh+l993AKopjdvCAiZRLr9gdeUp/tn/v/TVaV6bvYEq1jPOW9ewh42fQYpCJYOY
3vajmPTBT59DX1CGTzdr4LGpWGDhN4/KpjZi2rdQucCGteQHeyjdyRVdgF6gafDPuuSAwyHc/BWx
ZNbJkn688ATxAIsAuWxkdfOmhBzNAC9losY7RsLSdt/pbuqYB1JW0oRhmco91R+ZlbuMrxR93hWj
AibyDJ57GbauWFGkDmYe1hesf5mPa0TL9C7pzw3veUQqVD2bDgKMLmLX7kbki/xr+obn0DnD302G
APJ1sMDQi3Z6EcjF0k2qiVqXg8DRvuhYCr9N2tWwaiSO7WYyW5qZha2QEI1mMEX9Sg8Jqno5Sdwy
7vwu08gcrvGQaXN8jExPMbBKQTLzAc6XB2mzveXKmy93F+o3U12LmS//+2YF9RqUWac/ZXoWwJn8
ULlxT8K6EGi7IbnGrL5McfBA/gZds/puZPB6l7UnjB9HKo22VSnrBO3KPZMu2GvSfAHz60SaARcO
hmLrZhh9QX4yu626jXKlSbedWwTTgtiCaB4OGmk73KgYJF8soQ1bsH6jNZ9TZmSPddRhUvoEt9eu
FO++mRY45KwlbpPJ/Fx3T755AoAjSCYtSsOOhw+vbn+tOJ67viERnpp1byfptwypTqKOJT/OfHzl
NfH+6elS+Un3Bvo8A6TIPyyBZM32UyA9iJUyCC6jt1F3pglXNNm/JlYFuPtcTfRRCAoKY/DKUkd6
l698+USu5c5qGlM1p1ShGmHhzZkb1BQXVK6z1LRxee9Qc7E7HQPe+CCz2UvM3Yy0S5BAx2dDtqAG
tQY5HOS2xG7nYpCFQTXukc54nsQzump7qiKItpF6IAy2VEzUlmM7eC3Bi8/mvmusgAzt5ZsZE7RS
8SDhtQD42XTiD8P9gyGcyzBUk8a5Yrpm/eH1lskhYn+48tGCZQLdm6U4dsukm5lFIxHW+AVo4hnu
9+aDE0tBxvkdKTqHJ/HXfO0mYPEYVuQXowG5gxmcTjB1O2ypfHn2pj1t1OWnqxQIVDi5rfz+4JGt
jarkQXk7oHhwzymOxpOUF3ia45wv4MUod4oe/rBbf+zmO3tnw3HVKpjNaOalz2+HfhSTM8a2qUXd
hX6DreEhx8g3gbFtseEU0P2oR6tJYxMda6NCtJ3ilFlVu8jk7uEvK3ZfeOQXrSBGPPKPDO33569c
97oMh/ONAJoVISqMZdVfgZ58jyOYoLHQBB2dh0B2fJyJUip+ktS678T9EYK8wckeqwRQt9UaOer9
5igQ2yVAGa95VrrV9yfiiHhAA2fOCJkv2GKjcTe22hf1UaqNPxEdS6ZfOYoZTKJKgh1iLC1A56Us
0JSHkF1psVkZK3wB8ZvdcclkSX7sfm/PsjcoGjb4s1U5XSxpT+JRKXtVWnu//aJbGsZ9IEwTHeD4
EabCQzGugcZIwki1ELs/4vCFPa2VRMiJladzzDGOGLb5WGuD41vE+Z+bQjcHW8yzID7BlxCFd4WI
tFulSxVJjZ4iQpt4Rs/jO4hUoLkIQumiArKfSwUFoubWV41S4WScL3WbwJWmHPBT8I6WUmELoPyc
gDJ353jVswejedxgb0XxQxJZ/gSTvHZ9xYcOJ0t0hGQx2soU0Tb8ZisxaMq1WtTKUgYZjQDPGvkp
gDnDF2pZAV6AocnjC95g1qn3A37koHusV/TBDFVrwrsEDVHLiMLbxPd0SMgaTuqThm9AmN5mlXXO
Gbm1w8L4J1iDhB/mFfYDYwXsMIZOIWNRxq1LoDVwdA9Tsbf8Qx6X0vHrwehpkibhZXZ5p85icKKO
tcaE2DUcIxIlBNv0O4vpivGZ0b8OOrsooqVqysVxprKqF0b7bhjF6zb+uWT2mLzaBCjImlanC3Ok
6xtytlpaAEKD+PmDgzEgz3wzH77MuEj3juojOvgzioar/lnCwKB0oQ9KMTD8viib4/jTlJYaIuue
ntPT7ckAH7mwHBOh7q2I7VZixCo9Y4Qnv7L4Q2H5ZoxHVPj5MyoAseeLtoeI4WYDFgrcQrJ3oL7B
kUid9mvdfmY6x3WbdFyAfkDJm7qKqqYUMJHDw6dT0KPIPvhfCnaEHY/Toks0XHBDZkvlLsBbUbpu
B5pdJ6CnnCpCusEKMg3KTFHsl2BLoA58rR8c4vUbCNLKaPQpqmMvGfWRYIJT8fPaDfiJ8V7aIDxr
dTA59KZAWXUGqegDnTx6vBjbPa97JYspiltx9NbfdZpnx9bG9jNVeprsJPYcFYSjZsyLxIuVUkTZ
xOoOkvSZ40K3070tUjWngRERJvF31zj8/7850u7UxnnDdqu3qwttI+++Ci/jlBer8mQQgGtUvr9k
MApiolgvQOgCr51SIzMMin2uNZI1WiucGdq7koNkTWirdqUpfIl/MV7zT8Rrit6ZudUM1QZC0KZ1
2IvGjwQxEtKAHWs74tIuU8Kj0tZXnuStbK/2dtVvZ1HAqx3nkAcddl8TpT4k5TSaMIX5+beHhq6E
IT9UzrS/8pJhWeasCdyMvd/5RewtCoQjSFzoh7JkLYzKUfwsHWMy04eDsnNpBh/Ba4FtqKmzGRwX
0nTMcJ111lGfgaLs/ijVZ9unWNHcfN/0eYHa76MzvLmBR++GoMkbmGG85QFRueUA23ejfd34kq47
auGSOD6DQGyjzH2xzaJAePbf0WrYT6CbC9ISy1NIhXV4Nt4JSdIbIxxgiCUFaRkhl8hYL6/Ed6xj
UlUnqHCMxi6S3ZzTx+H0rgKv272/k3XnEjXOi32FnmIQvKR162tBQR2OO+fN38GnbQauwwrZtg32
xd4MzDD3tlDq+Hiym7eG00hBjBFP9cienuWZOHVio9/es5mfGlDa2wLV5JqNIh2HVmBMkiLwLzqo
NjN3JHxQUs2eoKBYTgbvvuOHLbc0Lly7wQGhfVZQWYfXUiuHZQA9UCVZMZM7PrSW1h6JXvxZe3sf
prJcXUrl7gIfij2gh9mdHZUKsTXy+LcM0yzsO1/YUTNq399/vFCwrkJ7stO+jZ065O5A3rl8hA2g
WYzAe/LgxpUEHlPCBEuk7vo2yVDnWrGGTfzqiIyzZrW17C0GgO73gVskZ6X101rNqa6j8s/o63zf
Hbc+eatUCkt/Zn3ZRyPG0C7i06e0/z2Vjg/f9LmnXjw2WBXdKCExQ1xgrGWZNA/JSqDoIg02Iv0x
k84cjgcGpE7YB830k0gXkdGcIVA2rPCKJFV9hXTEAXbY1iu9juXpD4EwwV+6fSxMMDC/aIO18yo2
hXUASE5FZBeDAXGAD/FackNj/MhR5tA9GceGupJ/Gi0LTb0tkalfyu2MOVJGSKxkUrZ+yPm9zZPP
7c6SqT+EYhOO+jGAeHt8NbaKS3c+ovO/2Z38pOJnfZrAMTCvaNx5zZvtgxIkr9fNt/+3kZyKH33x
o7aEpPKaQqwR9F+bDLabtUSQxxSWqtDnl6Jud3Qf1ZbuLF1pBpHQRtLCdqJ0ryvTBaUerVJ5weCs
rrUo4u3sMt3NKVOqqwb5/SrnSlNgQIG4IeR69NZeUX5LTIdI2gQdqPxnxkD3zrVTuDDvLj7ZJMdx
r+cxDo0LfYtuUUvnb+1HPpgivBfxUjTEAMxymbzR9i4cwBHp9xXChIt48Df0oHUbtqJra+mpBuRt
OV3n79b/WWcANSERcq4v9mGrKsuWIiaorujHgINbWAEjMwocBHhum02PsaxqhFWa7BNhkbef/DgE
SxldpwsZBbEXn9ltORh2rDwmSQOb/ALM8MX50EF/oQqJrWiqbSYbvOj6J1aRNNm1mvvorkE2O9En
q0u4OiLh9I2b13HqlSeE26jKM8tkwd34wkbiTFfFX1WIFC5Iat2HlgIBfQxui+nnCAwuYEJe8zY+
VRrTrPf4o3Zsu4rOtp8QD0Ek4hdqc3tg6C8+lePi0DNFSze11088oHo5xksCd45LcuOm88t7MAgx
7VvrDO5YTikH9N4mXE0eHry92TrKTfv9S8lVTQfm1Mpbz++k9u1ylemVCJLmKgItaiYjSpi3qKx7
hk7IfPIoHvhEfAPrahAk6XoIzaFGT7fFqB8Lx2TfjG9Nr/v75emAB0OXqDKcueswOyU/yce3UkUz
1MERwHIayGuDzjbWEGLw56itzLmlhXgHmXBJ9AD9DLX9otS0gbzIMOJNtwrwkv0bzr6wt16Folt7
LdSRwLruM1I8+VNXKTHgAu12zPugjvS5dnKLvBTKWKgAaSVJRpRNJDeFySyJ/L3Zc7hiAqwltyIV
FCVAtWefT9l2jZaVmaxUavKnCmh4A4BYZVA/icgmtuD9Kc/FNiDm9mteX35HT+l3vpGHhrClRgBo
9DZfzXizjqBQfRE1uo7S4LnCeEn8klFmA2ktZFp3jw5wYiFXrQIRNTPpVDt47BPSBcPT0xB5yAQK
/AXiWOlo+6l0yV9XAxkquN5B+/eWF5pa41lNKOJKl6G5SVnTlokr9W4TG0V7dN+5PQHCfnQ9XZnB
rhiWUqfcDNmxzjkL8worm15sXP1+lM/d6ifvx0F6pt9qGYs98j8+SWvKWwwSe+NufQYA/W/g8IuT
mpwq7yw3i8zVSk8IE7+doZQjucLwgzJ6ET8DlqPaHQmG+KyFiWGp4QyNiqLXJipPhUfYIkWmgiXZ
GtQLD/Vd7hgUV4YMV4lPchDcIJkQUspxAsjnHGErR2x5hXD0P/qqEcLn+gSnCwpfEtpHviFn2xsK
vGuS8pmoaZuznDQvdvaanUetxL9SJbEmK/Ond+hpEds+yAK9C9AyL/UZvLBW2UicGo6lkLwiLAQ5
Mq+gPzf2v+o/P2EoQC6qk354ETSrfMkEHAYlOc7hQk6CCXCw8M5W0a/AaqFb9Acmava3D0jUih9a
QgDaVa885wqk1E0q9CB8+Gj+0c4xnMVYHXLhHhiKPLKMS2UI+1qAL8mfrb3C8kD8jzJ/b8w52Q4e
0ZiL9RALAqbA94SKRJaeMKVSFddHmqmrmWeG2t8CUJfce42cBu0N4SKbGZ9WvryPxd28bcbVj15e
2NMOjBWliadfpdUSQ4sDZLFD2Gyqcjk2WmcyDGmFTFuD4GFsvl8G2OM4T9RXUYrfuphIl4JBAhXI
eRlhZ1lemuyL04j+4VSpxC4zphghK/aLsJNg+Z0pPzKS/pyYiNbw8tXas2JBMmjwb+b3Ez6mYxLT
Aqq4yX6zJglt0XOQ+VN88l8/aGwvTN8nElOJFksI7CJ9JZfa5WrUCwwel/xOQkXfU25xNzbS1scv
PJ3nskL33bqCvqCqJwnoS003EqFNFWRkEWYlEnRTwEUNFtr7OAlK2BQmq3ec3BuHuk6EPaIUj4xq
VU0UEMla63Gl+vIY2v3XamvyR63mEWEa/BDHbWyaaVH3PU9zG7JIjENP0Xw4Sp/K2N8CC5KjQJ4J
lAMgWbKysBZKLadvnMX++lPFkPaUY1pODd48XgDb+PaBKw2F1rh93vLTlIsRVj8jUvkaX3N3ySfb
aKIrVmY3R+gYN5QAh98HDFa+c9u1rcxQqYcWXxoHJsH/C+epBmTzDSKWsPTpd1XC2PVYoCx5M3X9
OlUIqdMW8avuo7tP+sYdI7GzHF10VCIlCgun2WxJAV/zsb2BhDlaRJVTnjrbNeMrHtZAmaO292S8
qlvEaksXR0Eo9J+ddoPVppwE33Hg6xOuIn/4jMb3UtkwZ8Dw/a7cpOOCSOAx2GNgw44L3/RGe+AD
m9/ZRvgT3e9x5PHyd5xGjC+7uB/rflikmCV0Ma2nWcrM0vs2jlOEbZNpeTsD+LOEZirTcLyXHGjE
AnHi5nLVRfLZTpaSuQNOIgaGVOnFiR2xczyL8NpF0guVPMVL0qnwsMm4/dP9OtRT9YJG3laYR+yZ
8nYUs5CZDnL3cAZ9N3Gd6eS3HRVYvj2OBkQXMonZ5nKtBG3AsTZkXmhHk3IH+d7HRZ4QANL+U8ff
1OgNRZ+eM2bGUXlvEey8zJ0Og4bzNX7lKO+bql6VZ9jSjsxj3jSGxvr+Lr68X/xj4XIM9Cap/Fqg
WS+melMqkN7YnfgOq0sF6Ndhp7cuJHfqus1gz/5Yp4cOmZJX7UiCbgGojXJFZ9JFkdIdyOJQhPxa
pyMhjf7xG61GPR9S97tCObILjGFcwNfNPtK82+j4e4EoUtmpxW+ErZW7VXi29hnyFYZ1OwmCmioi
6RJNNT+tLPby+N/PEmcc1Dz1G0muqWnvuGBsVLmy7yyPKpBakumV2mzyWgegPjLGiVyDfCnOB7vK
SDu/eqOs7uVakO+nhR65wvhIqwI7QSz+H2SZJsi9OAF/8VJZY+6dHGEOods6iiyMoyStpP+UGqZX
5coe8mofhGLmKxDAHPkuq5BoojbJ9OUZiBuSjGiDY/z3VVwcwArvIcFp7fdit8mq7g7a8mjoLwJQ
MPNQbltNm4rRLosCRiaVMVimNFoYvF6URtM+7AK4In+xFOwI07SAaCzEu0rZ/OATjsV4iFE624Y3
d7oDfLYCMu97w1JetL4T0Mr+oXilOcwaPOb4U879nmRa3CX5LL1yEb/PjGLyNS2zM73hZ/ItQygF
YtZJkZtHzkvTh13SuwTx7ZX6q8StoBV7fua4VjKZBUqv3iCxJOhsb6mZLCozwP8LEeWe2RVsSDkq
UYzD9RDaqD9ErEcBYcZEh8xLZD0as78OXHylDx+P8yjRCmeW6EAi/pvakCxVZ1cs7M/snFUbepGj
dduzUR5TT4qB2z4PBuwH3ZRY+f3mS0de/i30YBYgxbvp+E+uhiX4jMGLxNXtvPOlzp16lTbrO5lP
BahQljtLouXf/PN9vg9++ZZ9jK1PfgdvzDQ++x68J8zNrqhAtClovxsfaWb2X1nehTQEu4/uUnZ6
QRl2a8kjDTDlepnJ7+JsbefHKjyrYQ8AdTy49Vs2OFVVG1tLL5RzWwWvCtvcDM6Q7cfGzVdQwkMn
RkSXT0Zo/lLEeWsM3ohYMVxqNAFrqgxWYNv8pWi0USrU8uCozOpijdkF9w9wd3pYCDzlgQ33eInw
iyJ9bEvMCxa1f6X4P1yo54Q4pZTVGpBCfNUFjaEGEnNCnUhEio5nB2ImDfhOkKaZKh9PkDlgOtcv
kDE1SORPa2Arr3XieKPIoFDo4y03kkuukWsmKiOULdq0OrUHoxmjLCRHaADe9klfRQ2CwMlhhJrn
HGmgMgL6/92IMpzHoqNJYZnRYrM0F5MuhTU2FjCDtJzuTAcdkmlGBZ6VHHxr/d1WbGsjvhcIS+5Y
rro3RtRMQGIHmjc9FeJYFzNwLXLc70EtLIDgWKRX18bCrjChpLyQwmIDgedlZff5/Auuc8ZCM9OR
4jrNa5H/eWk7ychvbvWl902LtNXcJquVebl4U0BUstwJkD5Vb+wFSfrECQe0eM1xXiXqG35n6GAw
nD/pcPiFrqIgKIdex5CzFVc5/qmEw1+Itrh46CHSnJmHYJw8/ERmbIRytWWgx1eLjgJvDbvUuVBj
2VjscWdZXrRJJqtVvyU07wsWGjfeANol1w34jLoa/1bvjv6RB1i57bCRE42OwWaRs74n7wBuD4R0
mqakYiFsEfZcd2sjXVGwTQBTwW8mEOzWXDzy3ATfL4butv4NEc57TIAFHj/RUk4IjxCZWzTEYUzt
pzC5+8ZVTO+gt77Y1ug3RFh1NBD9h1uWeeZAyWJihbT5N049GKfZ/fpf/GZwPy2LXKIOTscBQhiJ
01ojs3JDGcey4kmO2MuKIDvh+P4LB+MPwHwbaua6/dEHosNPP4S7LGVUPzBAWEnI+VbMUSC7PnRj
9I2Dd6mB/LUpU2VLXL1DsyQm9Too4nDFKfsjbrQTx7STIYXk6NLqfg5t96/o07HeJLCxrR4dH0z6
Doic7KQVdMFBdONHajPS+Q21y1UScglhv3HaBXbleCnsWumGTtfhphtiUi8XvRpwX7yXaXQo4rcW
v+b9o6Z3Ks5AWiHfl5Ow8o5vFvdZP22V04mpygG77qsE/57xJJt4r0jbIMeDmuudkurZ0AQX1Lgy
8fzkgHYc0IYkiil05s+rQlaM/dXpGIboP4O3lCWoYgocA5VO1WpeM5IGA1Rwo8m/A3c7h27GLGL4
YmcDeVC3GyxXJT5w+CACjY8yz7+R8q3LEmrptxn1qoKVjChxmDSyGyfQFBq9HclTWvXYrVR96HOE
UCJdxoWNHTxDoweOJch0dg2l43PLDI1BSNQWa7Nq6bBPWzEL86Lf4zTO70bbxL3VxV2rd1fBx0Fe
I01L0+6IY2dUNNr4T7FmCqmT0xiUT1aGLNfaBkfNhuP8jpsTzQCtxFpYqrOBj+rdOK/6FyZTNZ27
uOhegCwqQh7z6YGsNVdHnezqKVM7fcZYWsLk8DMqYQeM3rQc+kpTOguQTOcbg+GwtJbWOkMPceo5
6hlOmbx0qdcCnDa5CuIKb7KXVFRGrXLIEe4rxFXM2yA6dVPeLiskIw1SD0fHjYt5HQA5bskfupH9
LtlQPhVqVt1xkREvUM6sEuEKD3FYLCTdfCWfdyQo36JZgZs2hj+2juh6lnCGLRTCJX9Vch2MpH0n
HEcsrtqDh+xg/WppVLKf4K4osG7XKhd6pyLbW3X1CxdKGRjdGjxbgTS/Ymh6ykNdja66HLCVnDcv
mgJCK2rRpOMU41aM8mJBiBj6g5rWRgrC9Vd3ONf3fBxO/0ooVILA5ukbrRxMkb5DTNwFiO3zMbtJ
sBN7H9JRqThb8NbBooSLQnrmlwrh/Fv/s0eCCzieN91t1XVjiGcM1FtD/HLaCWgRouR4o36GKNhe
IOEFVUVh42W6sTmiGBeJxLg3sjJVFJUrSYBxEYg9HIcxj6GUdSvPG8xRkXbPoSM8CMV0vp2nqMzN
G1kNdkYDEjVUGa1X/Ww/DQtkPJ3KawnONDH4Vv2XFDJfXGxo0e2o2gKvCAQxqeM6qFPBcyg20bF/
PEd8FKQGGDi0Z6JsCc18LmMCBPcTB9NeJKTvJf0PHIslTSacDcOewv6vvejyvxkNheVYr9fnk2tw
/EdUhFK96BJxwUlxuKjb+dh1FfHSBWCLSfyRveGp0tbYRMmYxFKP+h6F5p0cRlaUdg2Cg21dv0I4
sBwf1LcVLWKQgaJ56Hdf5scnmLlxTvnG8QIyVe/EIE2RVwdo5JxgZHQH7F+3U1mLC1tR2ycoUde4
qH/IXegCH6j/yFK0KAom/dZ2PWpw3jQlOdnpvV5b817Lz7gWXtpdN0UXpH7ZF8IZA0wA3afjBVTO
RVIiJUx65mKwapWnEXzjbFysAopzhNtqD72B94mbtgCya/FdqNVsYu2MZVyobf3l7aJte2V+z9SP
1cvnlL3pl5BF0DUAMIo8VBzh3vw3AtwFw8r3zzYTJbtkggw+cXPLTgsf1FJjHx2ySQIQUs0wVRKr
hhCBc8yuZYsvCxnuNKjuKtaG1mYe98nqwNkSDJoWIdsZkMGki1cR9UeAguj3O0uXJ590AVKB1Yni
4yRZm9W9WBwNNNWeUHSoDfQFKcdj2JVTIZLWp0tmf0J7PUnOqfot9wdghsLMhrrgzytUtD8/Dh2d
90TL/9dJjZQ4z7LjJksJ5/ad4M0CM3YStaZGADQWEyVSavfrClAuy1wIzvjoNvjVZCVJwkyj7En4
Da+pbsKJDo2l57BnAZUd6B95tARQE0pw25CozsBIfgyiln1BlukRsn/45MC2eZ6pWff/KosvzTbb
xrp30e3t1oxqjmr3jXlCQqqM0jaOsNWedyEaYRG9HIrrZhIJ8Bs4gaAZfxQsb8gYf0OdhibrW4Vh
56Kad00cgqmWC8PMJsroROKHxf6i11cgnCbE1F+krGpKGF6b5IfLTH08a8RxQFTLeZ6fBSXgl9WZ
JKMlLV59y5Nm5PHeMaMhiTkyGFf+X8WwSoDvtVHDT/zwaoxZ/DeJR7gV7NlOOtwfIQd0wXYidzJD
hToUIRpjQzSYHp4nBGyfEt36WD3CAo+XBQtGOw5FDJn7OLJ0C7Rce5UMxWA71qc8wys348iciuDY
BlAA2b4TfyWIDIgoHXGc91tU4gGJWmH4NNPZZXxBx8+sUVdguLiH+C38M3QWnt+bGGUXmWeb4wWj
W7h+xxJoluo9Xx+JWPea1bOhAbPZu6DN8f4OmYHekVpJE4VrJmV5/SiufPbzkb2HozdknwIE4xWh
yu2b58CpWr2ZRKSMy4NqFwjIW/IH/6MvL/YRxnCeBL/PWKnkIidHf+WEuH4JzErCNJh8kaYGi9UD
+9QNvzINes+CFQdA44Cpi5YrvtWVq2Nsgu/+/9Q7u1keCIYQGrPWav75GHBpWsxZHbss8FJFWxko
jD+T53KngwZVJEbK1fReGlNMNM1D+U/86X7Zlt6SrNHMJChxyEORgeheU80R9pNzn3LHTGQ4cKMI
qgCVJjfLcEMMtQrr7WAkLJJrCPdla4lBN5jVJCKyHsU5rQFo5zgZ4vHPOO0Wdz8ziKCnfMd1zIf+
LEOiSxrHRi3AtCqRDr7YEjIjTlBGYwRrOHVeM+JQinkRW2S/6p0GTbsGIPjmxBjOet/vSnUXshYp
ckijYxX1U0o/h7faLO2M7VyMBNyNTQ0Ug99TY5++4RVKjzqwvkDsXjrRo4lYSgmOrKMQpLI6Vd/I
NRvIfoykh++w6tzKH+fPyuS1Yb0lecw9gPcsTs/6aYWWWsKcPQxXWv2lEN1KK/eGQzYig3E6g7Es
RoguS9LYF4EmxzihnF+cStyxDLNgEoMkIFGcF1z3QB+Cq1mEo0IkmOOBzr6ZCBTZpmydZ5oElDbW
Yv4+bk9LFc9Lxz6yJuHcbiPr28PycxlMA/yyAv2XyJortDJDozwnbnrzJRViIIQD5XbkmhPZiXKw
2y92EkkiBAryu7pmzXvtKQPPnyIP+qgJKlo8MdGQ7+Fr7oaV3ssTCZqtbHb6kqPoka/Q4W+UVeHh
fLCE4AjwGdrEhjqrOSaJE12WHMjlct2QpBzxNy/M6UqtmTOrH67QpQQBUhUfroCSaPDoPOZdrVks
3qqfoQd0CnHWteitfywnbodf1rMOhaiug1lmX4LS4GQJDtyuEk5/tLOsyiJXNVDSn9XROkpBvvTq
ZrZKz+V3V7QATXNV6awyUHynckIJqBY1jRM5eZT97Gah6yyb6H1nUmUTVy493ADmsBdkGC0Xglqa
r897dWuOXwTgrUjiRwv4rwWxqbNa8MLBL6Y7itavibHm5+FHbnRd+2F+DAikWHMwMYpw2DBf45Dn
YplhY/JIPv+CLJuTLtsaKCgbppvd+qstUg/3ihgwJpckgO9L/sYVmfLxDttNQQlx3qgI5Ur1juc/
5X/0SL8OTLTJ7RI/i2voS3vcAUNni3Eh4EkY9hSQuU0E+9ocTYaGzY+EHys2UeMmzXkTHvNG2oFs
Xgre4xFptZVmfrxPBFWJ1MOx+SVOcjm2i1y/yhXCtYCvlb8akip6TVdjz4A6B4kTi5a5G11GczzH
ByzX8L4gngKYwFJNBHQSHMprNcu5WwvRjJU+7S9ffF+jmAMhed8Xm7Te5FRTw4KjRKHshpeaNw5Y
CNnm/ZmYuM7S48jl/JgWkrIZO5YUHvGRM/2qt1xaqcRo/1Qibe7bhnmwWgz62fb3M35Yn4+2I6/U
BH/DakDfoexCrh2Yeh4yhJP1KwiZTRGt2e6lqj3oxwbCFk5BXIVGWHJBkVSYygDotlwv9of/jeVB
0jcdPUPUVc8irLk5U1iPTl4pDaReUQzNp51cIw9RIS8XaSjfS/uHF1yvAasiM/fo/Z0sCdbeSK9J
upEJYYOWjnOWP3O5vOAok8ePicIUu68IrejS2GFew7AdsVzZLniPxAHM7ci+iOeHiYEc47H0U2oB
Wrr70lYHGJphXZZdvKJ5wQYAUjvuH4ub+ld7C6P3Ijdt2oxuj4p6TaA4eP/qyi6eAU6VB8Y7GXJ3
78wNQsAMfm43oqFAWqS38RxWrQ85GCmJDgrzLn2eKixhwZ95bW/CYyrhKmVvpbED9QEGmMBmlJk6
Ljgm/htLbqgHJYeEqKodyfPmrzZ2ADy2z4nTUSWVHvjoN219AtgsnTFso36zIye7TSi+ylji55g8
R8CFjBCVYVsyhINi46f2ijA7xy4aOHvA9eyt+2Ftbo2SCLVpjO37h0ruzsfIO7Y5mCfAcM+zh+zS
T6CaSQuPci92Y/CKbofAKAorVPMB4RkuPkxodWy2fLquWmx2im63M83cwvUED4Ej9qdFpsCxIuHf
+WTkCnowOXLianShvD3Ev2vgDHWXSF0lbebBNilPKKuOVnLXJbimWNz6QSQrib0EpkQR6t/eZWZg
GMTHlKscEJW4iIfeqEetOYuaXAcAzbOBjPX3JiSto7iYEFJQblMqX3VqKC90Ks4nr5p5VSQL21qd
nMHww2DlaDs8bfJjNjzaCyfQUVfF17bzLhvYCtHhYayyucpvjslVzZtIBT1hUTQDD/1752N4FI4P
ixXLbLG+tgrZOcL255Fv5VZ6JxgvMFbCrh0ydvHpDWJ6UjKxy6oNcbDrvEJSuRUyIt+yq2MqA+GY
7YyTd7ZGLSP1de4tmTvp7j9DjxItdBL295DRf0/b1KAsgzK0NZXH8em08f5RcA38mAedmG0dfIp9
J6XlTcPRXpAqoEDJ/rOD44bQqxFcjH6TV3guA9uLMjTVywBgPi3Txhy5OFeNmJwZCV/ORQuHbrIJ
jiYcaO8iCCj/dj5Jq+GnYGJJOpN6dHwKnNDn/efSfCS2YqjCOZZi6yU9FmjznMHbFoV2ZCgNsKIT
zGp9O+YVsAwEAf0IWqEqgAlVbb573ieVaFyqrb2wp+Sx+K5VHmMDYalJ7+va0lW0i5NcakqUIAj7
ry04q2IVy3xnFFUTCAZ/zrg0npirLdlb9Hkp7BtvEeos04m9mtBdZ44IBesIPqeHkGiyjh4coDva
pNk/ELNyMGEmMp+4poV8PVnwWEKU4Ne9osrqgF4tlJoIAxJoxsSz3tpBMRt5EZTtDBMdRzxk2Ws2
KjeYYpNL6Vhx2ZSIE8AQFoUo/6mhhd1WduhRMozV4Bg8JzcaZpVVap+CT9JALOtV8wweG0BiT3Ih
3UXD2drxOwK3KDIlMX6qssrjnjIssXIfpKJ9AhiIrCx+KdcFI0RuqsGGd6h2ShF3c59KRbBBxXNC
/Qx+2jGgTEqchzhE26MR+u1ehat4MLmpphL4G6Y+5jDb2tRkgYwQtmXOkq1nhMTsWEjGjuzuYhSS
SMHgSL2uM1RhuRj6u06nV4XffcGsY+559wtrumJeZjQXXfKIDVg33Tn8bIdUetRiLOKMz4H0eY0K
tO8z4gvx85N6zN4sfXE52oBlFTZWXr7W01VsPxo+o1p3mLTVCqn2D2oOcAvEK5+DLOOo9MbtzB3Q
QTlwq0PyXRBx3NC1r6c5zthWomxjMbupR2SKEWmlW1+onCIbFJBLShIZzH3tzDiApUkYwXYAhlE4
ojV782eCk882YPCvRmumcidjs8NEd6iGNhaM7V76BkvmS36oBDku16uDIXo8yqEfPwIMqwEU3YC7
c2lJ7iBymjaW5CatwXE6cGCAGTRD+RdC2Lpx0HkOs/5NiMXnkOSRlBccQtR6qLTu9YK9RNrOg33/
aHALarRP7Py9scprMmQqf0ngu7HFmFMVBdmE3gdAAPdhSdZhZO4LNvZ4ozqJWfd1hTWFdcdynk91
CZX7RYOmorRy+/9zxDcH8Pq+q6CrFC64lhs/CXOY2UgcxwVKN+npaU1qaepVpjFlGP8NK2M4P9W9
u9FpX0+hgXReP1+RNLCc62azsldT2geujg9+i5UDDbjEyfNIYcPJiiQYc/XyNRMoZOg1FRJHNua1
CECE2NSOU/rHBpDldU66+Oo2perwKnBh2LwwMJ1RQIPKsO6aqwBB3PpIXwBkXmYC5ybfpEyvw5Z1
BYfcUKAcwU5N5cgcTdpJFiaeVnnMyUuwH+cvtDCegksEy/h78P9pnZgwzQkvv+rFQzx+PPMWb796
7pIMYM3CpeecBgPvb0LUIaHx1ccehlrhVu5plct6I/XwhUlF1OpZO8HPaRFSow0utSxBhzhMCUWk
Krs9BB9zhP005KhKUBQex93ykgId5h9FFN29WLCZ3ogEQf0b6rpvktLGkf+EadfkeuyO8zoN2CGa
dastryAnzOURFk6hjSs7auqoOwixXE6wHb+igmUxOoz9Qib0Xuello9fMh6lkXD/QQaRKmNzjfPH
AknSfZfl9UlYgkqvPybd1t4vHvy2jyQ9JFIQ9peXH1eZ/iBLB7l6apGqY/5LDW6GgnF1Lm/8O74s
OHr3iCS/RCOt1HtURiBS9ST3xOXngvLu1TRYXZHeesZkN+xiTiJ2KlW4HPDEGhgSg67nkg3YO1cW
qx2uRKtRsCk96bedHum3NAP9W4e2prk28nMaxRuYADt7HSrIAkRg9TRKIIajayudX3a/VwPM2dCK
OqxLihUx+2GRzEqnFsL7LkjU81qw/iMl4UxBwEF3mpDMBzGhHRtY1khWZ6KLLzNT/T5r49wfVPuZ
uBgTWOiIEUEhkDjAQ4Uihp+rAfr4rJbKxnAOoxtxYkaAX+JviRruRW7C2WUOU9GS0xzWvGx8pcuG
J0HV/rdj9m7SQcjybsrgAOlN1lGFcS9gsW5OKDhf49ksvnKKbpzQsuFUfg8kbeiM6gmaH/olKy6d
CYIMGeklAFqu0xn0oFkNneOkT+Iotafvf0bVOBs2kP8gxk2ID8R/g+qfFNXe2wHF9CYA/9z/KHP2
4CEvEUhmhAb2PRTuFgFpW9orlim62Opt5ypx3qUxJJuUKnmUHloxDjm4d35HTJOmFK0HZKZQaGWQ
5rj+8VH/un5RFmk0meP9pLaC0kfC4zXVYwIeAlD2HEB5XjHkIHGU2SvcILQDX+Gqlc7rDrA5Vg1E
tmTWsPG79azWa2DFXfeOTRwwc7/8wnsKUQe8qUU9pvyZMbmMy/YvjyrF2iHQN/ZWP0rBgIm85bKH
GNoZCV/ktNc7EG4H0QOHufDTv4lL2R96CgOCb+qvdpJKjNV96WP+jeOsSpkF+M6vcUAtp2X2u1oI
QMgZYiMZPwCXZgMnn4sjabNIfJXZQfUIByCGVbNjCW8QP3YAlEMRZyuqoC+VwUt3kEYkvY1Apj0N
SAD0m+2j5LdKpzJJXvwejkjWOdZr8+AsuT+7B6jLjWEobLIIzMfaeodHfXDfDOWli1BcokzvEnm2
/ZZIvjvOB5fS1+DHnVB4DWszzkr8fTZka/6lGXbgxzJICysPyApXcm1cTaxbY6/gYNmUCpfd4paP
MUYzroROM4o1XaI1VTVD9sS2ZyvnQcxmYvkxPFEFKZk7rHc8VMFa3Q+VWEr4v4zM17gH9ysBJHKG
N1TwmeQPAu1jBbAcZN6bBv+fFKk1H1tp+kj14WUYi+6fIv0iMKtRRDVMr+LsvoNUlHcCR2NkqcIo
TTPRCBgJ68iqSseSQWGmPgVpgI2CK+lHQLdU7NSIk1iRLuhel9G8xY1CQhs+Huo1XcZeWCI+C2th
lIRpeXPGWmLb01J/w6+oxB6wBaMEK9rzZYIZr9b2DNjuG4wCdVf1i9YjuibznuGJdcjZFqG0/jua
qpYg7OvQ5Gs6anoFlhhWZg4wfIKte6zEPSmgdTNn3zfP14TMui/iS4ZgsBEqJjaz2OkcVDasi4Tp
2J8pwID20Bv6f6/t5qNMK2iiAA76VV/tsXU1C7i2gfBFKLdHTLO58OIt5IsqPnmUuKU3Bq+n/vL/
x9tgEkRv+J9zd13F+OjC/AP9s/Eng4mWo+0hGZAwUpxKNscoVVWcWTOS/xoGU6wWagLNmXetEdHM
r1VJW7AMBVZDPOgSrb+yup/x9q8pMv3ljG/Qx8uk7QUXL0SXAsMXf9ytpkRTHErA49ZqTtZGMllN
T7KNby/87l5S1CyLY9jVUeAbkwVstMVB8Ks2jj8yEoXkq0wbM+0ghjezXlEIgbqtA03lNBc46ad3
gXI5izXjQNmhRSi1YZl4nPiCM/djPAUAmfL5aJajp93O3jsNwp9SXE2EFzkeMQynboaG6KQ/qwLs
49gXjL5ePkLHFJ0MRO4wNG/vlTYVnY5Yadkp+IwX+cpKahFP3Mko80XPQ8FM9qx2ogRq/dIuwau5
k2veWcs+/5UtwTy8GtLT1HyKFGusuBm7tRdQt5buNMwWnpuxCSx3TvbbQ+5vmCW6yre53sM0tdpe
xam4enNoVxdrJm3yiS9LcnQko/c9b+qxHCp0HQX7BR+q8Jr+t76jd/d5PiohVPnNBpUDsejoJKyd
BXwksPIC79kfBOpiPl0aAb0uB7NOsdzCKWkxHzBwESAvTrBkDPX39fiJu+9PuI5hVEIx/qOvfAao
yDdMYr0cXj1qmIZEjmdrEUK8zQ2ccli5M0lvPbwnkpYrI2dJ4oym8ZOwllByNtKdinOpafRA1pny
0dOVXl1UBA5uH+Oi9Lpw5yeMWbdgNn4iidSlRQLjaOjiCX1w1SEaiODvY0De+uyPaHDSKFak4qsi
j4EXc98P+d3BtsuDWc9pIES+V96mDZ+d9UKkL/2jeaKNPWx9WK0XHGDdPYJyrwW87uU8CxvyOuCf
f5iMtmWqyPPk2KCIzlG4dt9P2qYy7AoAnKpiSKk3vKeWMuXoX8dcFS1a5LpEgbLdoQxKZoyF/yTI
TKoEQXhHhJuM9uK0pXpbeIK7ipMoC0Y0N7jkHSGatJgbiY7rkkPKkEE3LMSh04vgqpviGfH7BII+
0jzsVSk6x7QhxKKcpFyqHH4FJRU1Ftj9tZZKd1kX89iYqAGwtUtyiK3/8B8mx+wPdH3mT+sTH+hJ
yCz8lKeTt+lZFZ+TC9exaLylYR2RTmSq1pMaM1YjFE3ipb/FfTcr0Me1YpZd1LP1+Fa9xaLt0wNG
6juiwtsL3kdNNpomQgj63YpVVqPhlfzv2OgVETexlGikZ8BX9DyPI61MLMXohONtIzh3tN3E/dI/
aJlj130gsfACZpp0v5yYE/qCALnX2/JgUOa6dKO0mkKFsTcpU4sAUsG4fc+TOhDMnkjPxno0u9Uy
hflWVYRnVu67YyDx+THH9UF1LdV5UF3LseCc5OXlAu1yrK8RE841cMWaMt+lFNJt9Y6kT+uz1mvJ
3ti/vV6ZAXjQ8IFz9fNKslx7JnnVSChNOAXNs54TerrN06/Bv3EU3Y4MIEj0/PHS127jNZjCRvbe
pV8oxALw6IHUZ0q51y7sfrmB9ZfawfHAfg+8Qhz2dQ7DP0mdCrQN3Byv6WcI58o9I8L9Pm4i1mTg
jZqt+5u7kCuFHQZZP/2824iGg+xtuad3KhpK3x4kEgY71Ny4Nm8gyHz99eK7kfaaMi+LNIzBBybD
PkNMNDfHdgq+UWLg9mvH0UC7u1/Ysztttmku6g/+1/2M9UtFz8iUX7tRwQN4Q2LaFTmAQNG/x5/9
hmoq1cOS1dEjiHXUXLx8IRlWknVsTs42t/M0wSpeTsgZB/SHbYUY1k9O4zzIRjVnDbFFMoYhByNI
2E+tcrZwgO9juk5zuK+ayRhf7DgmIfjAfGXvvMqNk7lr8PhwkDSOD6A3uymCHsoa7x1zMxTxTkWD
y95OXOCcf1rziQDtnt1rJTRjgHHMfScCgHRC//BgltePUpFpxj248Rm0rBE3p3DQKZkdLepffhgM
BLd233J7MNs8BUEVIoChIDxgo0okxYgh98l8kuLEAOCS3MPSNoG8qCxzAtSbMx/VF910rOUED+Ny
QDk1KFFIgH5Ad4J/ZHd4Z9KRVZWZdoMcuiGEUMtMhbu5lrNuF3i4x9C3UxCtKEf9DgJT4+kjbq4Q
lCaaiB+hrkMQnV/38Zk6jn9GmBH1aakxHXb1bCA+GT0nVt8X1HxBrZjofEZQRfS6GeRL1iDwt8Hg
NEV1UQBhtO8hlelT0GP23KxU12aPxkyS16/0OD278i8+Z551/AD2EgIebtiOCBYXFhOQ/VyGTVfG
DmlvXx1vxCv8AQAaNO2grAaX8xZTQRL3zmyKiP03SANCF/7dXnf/e0+8ClxLXE+NrukG//wEan6v
jS9uwT8SNmdASu4P1Hu1OakiMnrgirg+RWJUGQhUWXmH6eboemaHo28ds6N6hPG/OVOH3xGsI1be
DtWt84C6GvbHWivJlblIxncOn+pc/aX0Q/gtUH0Glt9znP3aV4vEes3F1QB+pb8eSJ7xftrgc6jL
Pl/R1C8dorpRF/hTYKIjlrF4MqGaQDqYOgIU7FxyT8He7ukWXHxxeZ9s33T4EPxmNMwUu1FNK0oY
+yJCwWbCuA/jyorAafaaY++DKHi2UftvtdvlewoQX4Y28ypjGR9PyaMYoel/79P+ql+K1q1mjgV1
v+GBFo1z3+gA/IR0ZYtfgLPdwA5jesQF9yYQosRPbu6f+jzaoDEjmYhS84ntZTswuaqS83/gAFN+
Kcp7+7ED65/8enfQdHGTLdwTglFw4KEzclM21wEOQzGlRarsBluwsjMo+W2/OGj3YouZLwjR99Dz
1sDgHZ/+m+dCIQkfzny2Jhdy64Z0NmwxhCciJ7DJDqZI3UFMU343vkLuh/xvCuFUbTyWPCegdMeo
jG6+lWJqCudKLCrsvevSmNpjeqzlO4IjxPkJOUml2Mtbm2wR/5rZC2b8oieurs9Sh8P/7zU2Anmw
boxEFChZZu2tvYQRqupsUKVURAwEo+M2FhV4UJQR9K7d70V2eObf+R6lt4TDlMk674w879x2svfI
YF8+SKw/kN6S5+N/DOWfa53FV0SEbQ6u7R83VpYjtRLAOApxCcSvGVFoSdpX1eztCGefzsMSBl7a
GW+YrcO1LRyEeLGEdJ7ssblU8ZIBKElbxjPop7H1y4gcwS0Dj3ACu/6Uf85FK9+3aSh5e9wIpPnQ
V4K1zybuBHXLwQE/hKJtIcrnlOXk4wOiYHTcfCP423RLCueP+Fz8MKvOl7Y28bsvKhFV13vd58M+
CQ4/ve3K0XzbNIVJUhpcBPnt1w8jgu9aYoU+fJMSl82B7BRKIFNhvxRHypuU29jkuy19id5uYEdN
v6orFxJwE5PYj8zvYXdGqp5GDPjTtlEZgBcXie/ashgFCu4VKcKQW+h2NhCURFeXwcavtNR6s+NW
AOED8NAd/FKOtzUsgJuzwFQ1jtSLyJ7ZY40BTwSghyfepG6nvgCsddturgGvyfrOlum77goyKX2E
NKGkbUpi+8I/bbhuE0hgTrsiCcUjFr9mjws1MaymFHC6VLJZJe0rs4BfnFmoT/YgQyKVVbkwPGtr
MPnJUwfhlTl/kXcvfGW6FV1K6rx9ZteMQny3USBgRQaMEQpqLT8+8APt66RwG2HVyKBI8q4qDWEq
KNc5ku0iOMX5OReC+2p2hqYvizGd4fGyBUqytF2QlD3zZdVcfawdus3B8sEqup/MMpdhFMbgcaxw
/fvgKrIlIHs2vk991KL7yiBAMieLcpsT3nszE8Vvf8yt5yhi+6TC/T8G3XLFFjW6nEieI4mBwgOv
45WpU7fUAJoqyvUCWb3FQuhceNrgWVKg9T+J7pkEGd2/5zrRNV172wALZBXajD1/87boeRJGIUXS
py695gRIGj0ul/KSe2q+vOBzXCyLQUxFFA2IFQ+3WZlxgFA3q9oS2ITIrHSOPWQsVbf14F8Fgkxl
0XlgcZdh4mB0xIZhVb9anZ9O8GmIVYLTv7CkqWBQTy88GzLrgkp5eUOwNvwrhnfSA+MeqMNAde7R
i83rCq1bzA8lN2Xw+Wll0EO7faxu2b0BRrCMUp0EJf+H+buMwl+IuYbTXj3rJ1D8rAt2CIHoDs5w
tZizchPcZDrIm05P/zI3brtfWroyz1enD5l3YctJxCbj+P6Dzv3ZWGX/E06N+V7EpPuclSsHnP3J
D5LWfcyDvjfizYcdfu0BaAm8/6EC2IyoIdeYfQ2J+UYYBqRrbzkI571mG2SwyLssMqoHTD9lToLE
JDYH1PlnAMZonvbXVTn+4NjAY2D6XfOUHVcvRAvVm39yd7LE7/s7GES11tUm6gWkkume0BHCi6b5
BVpRV5jWFO/+7S1ZJ/HVimYOAV8I80qxNZK5VU7IFhPAtExXX7NE37WM8e8vjc0blsiMpgAywtUJ
i1euAjjdw2HlvqGd5ab1n1RGwyNcT7FnFFbMyHfoMO1qCAMYbMtSgRygcwUP45xoO/YLc0kZv7Qe
czJWQewVBMgbv6pIukBPQEsA6jYYLSq1cVJ7CmY1GBsyBLb5PZrUipxnSMd86YknpqwBv4IUEzHx
/gB2nYrzqwqhyIbNDieF4x6uy0IQt6u54PxCz0loMctadLVBR38mB3EyRjuydONd1KSKox3niaba
DOfH+svW3Gjitgxg4lebUjWR4++q88y+rT/bLqt+KkLyLJVn21Bm2wAZ8aKRt6rK5GPq4SdTZvO9
NgkjIMTuul6I3ildteOaSfGRs+DedhEfsMPntxa/9biu3II7cqT93uvE5VP2JxAa4wS3LRjASOnh
mcg5aUX7NkwUNECFZSZzenaEzqxJoj1s4TStimd3c6akrL/AJtUTgU53BFxJCmH++LwvG6hQq5Yi
h0DS43wguD9e6P3D/mhuC7DuQ5H6upjlh27azKXW21O89nPNmv1xdM9QJIKLKWftNzT/WtMD1r0G
HaGelz7whev734AzhrhCp7qfPF2AdshltxcKywfJ9gx0BlDSu5ajTHYCvE2n62mFoBZtlcTdyxCY
1XF2Lh7QOdEbX2uk9slmg79faaQpDIAC1fbw9wRsh8fMt0XaW14tAKdxqYECl+tsResiID315dEL
+jE7zO8LT0rf0D0gmAzkGeLab5GXLvq4LAwSWgorytd6MkTVZ1g2r6FLAgGr5F5u+7DohC2oIu8u
Q32YFnAPsMa9SPXlB0zMb6rSldrr/NjIgTs5aq3F4EM0Xc5LzGTpnNZvlV7iYjrBohTeqhqCDNON
+ZWyYjbsFMFRxyQMWFyq4KU5oGN0uPB0A4ctTXYMoijV5/f4Oj8qiR6R5FcI+XDgkz+/9q5XjZPb
RUWFr+IAiYdBX4Yek9UEW2TqZCtIxbTHFiBuA1gmgvb2D/1kUEEQ5vI4UZprnF63xXlzi2zMAMCg
QFAXte/6VL7nfDTUOCMSVJXzPRTdZYtWOKP9ZwrOeoKAfKPS2PJIXoCZItuRqC8kbYXSCuduMwoq
EZvJjiLjDgiZm00UZVDYfnOeeKaelB+11bUhdkDb23oSY+DMot1b2nhyzhRyx5g8cDdaPH7gtL85
R+H5Pt2SsVd3CBI9f/w/IMvmTFOystnA5csBCsvj1K5bL5xC7Cv168H6Y+0HA42H4zc2kcrdzg2C
quSC/U0M8D5vQR5I9KceuEJHwUwiMCOGhykbCM+7Fowh19fkbbKATBKm6j7DrJn8WLvaKcdcKyFu
TBHpIJW8ELivQ3+xOXGSFMGW80V5Rh490ZvnTSDvH2rRooEGiiR4t+cao7QaXcjD+iHiyaGGIYoZ
8HZMUrZMVpEEaXOafrJLWp0zD8tbCiA1FzUgvamg8HPLbOlj+MqjiWYe87GD2q+9QF+Ct6LjMHZU
1ij5ecClOWw0PKZ7HmDDPxicq8MtmI0ItGQj3kcTpNicXvG6ZsnpInOw/vrEgvEqoDpJPGBU53Yl
U5XpCknW+QoxkY1PkFtPXh/Q4BRogSqGBugmlHaIGnzkU1V2rx5jIShqdWuRlJMscOzcs1tH/aLz
h8zUxGBKZEKSTe2IZTWIWykB49Cu8krBBE733wZr0T2OY4i/I6iSwuYzAjIWx6LQsLYZo/vE/ImV
VJwvfTEwNXmRZpPsk0EemN8W9yjAU/UPawzJOuTOfUfV8pHbGguLu1camnuLy+4bng3waUBxcyT6
RksCGeu1Opa5Oir9HbPGqSUofwNRuzyC2sKrlbPBsOJDBkJaazXg5gaLkUI5EHb+vKyMq1RyVp5J
N8GLGpVJ9HqOI76PIfyllk7SqjZWWI+9DSQzsdvMDlRp4y9POhiyYwJ9MBhnlStEqILhw4KLemdm
8/g9EnqySqFr3nQrKFFpxPOUssTf0srakZH264taxAnID3CzXSF42YHYzM4i9qH3nbDKNpSI1CkM
56x36MzGSucOacBAfACuJyW8rbyZA0J4nZkogooOKVPcUHfHvQ/FL94+ATScjLf3Mg/xO4KgqhYj
B65DHQUEuQyFQsQzobYSPUwKlApbKnNptM0ex4vZ0wHK60khuYS1+iQAjdFm2Nky4SwOWD6dRAcL
v0ad54MOGcGfc6T+HrJKnrJsHnEL8uWv8aw4OyjssOlL4KpH8FHLXHd/I1iy+Rzn/OUFz+pcMkts
UC5cv3mPSn/j7POcGPEb3kN58hGgBWAUy4tEfT+aHxaGjiPqDaySex3PEThucAWH5ck0vSRbJM9K
I1XfQxIVhsNX4l1LwOFGKbQ9zWea5uEGahFQXLKnlWuaZHK/ghCywdhZ2sah5sE4hrmBMaV7nGKX
6jGqemp4akzPrhqVz2JOInOTwQfOd7wbwIS0q8S5nnzz9a7ebnI80JogSHNrCRCOZizo8/GfOaIs
rqaHTl6tV4dJXv07i0vm25Jhy24+kmyem4ImimH1BM5AYV4AB4vY4yIsUCB2PKP+SF8cZPl3I0EF
EjcgT0uiPwqXR4aXq4I5kFz0uGnynHvCvNmF5aFHAIcVRvetzcQ8lQFIFrJL8f8Xkhd6ef+Nsgvk
Cx3GpcSLfoYtbQSeezEFq86rM/Xg++7UtWJyb+vPfK4h4r+E42nibxECobqDpY0tpNhYoH8HFxQj
cImBF7w0D3AU3W09RvTNflNjFiw1Qk+OL2gGb9dcDlqO2vvNc4JLPD8rKPDGi5X1y0/PzQvJuiqf
CP7WGV/F/upvDrgJu46xRj0NwEGqdGN8nK2UZstKUeKO9vvX4k/8lYI5Ll35FFeHThoA9WVv1GmY
ZxqFLTnFYQr37ZOaoKdp+lkWrRsrKuC6NQPRBVESS+8DVXehG+PzS2HFqrdOc4vMxXiVjy5JTMnB
puKbYPXl48GjRWSx5FvBDrQEERLNDso7En/J4j4O1l9oX2Hw5SxiKtSLOzkEjxmhplY8YYAe4U6D
H9dhq6KOi0fk9ASON5mfpw89ewjk66olF42CdZ7MC77zfci0CXnIMpiidbsKwnEzzffmPFgCtDSa
lgEg8fi11JMTtfQyovI2sGOZtpV0sIH0NzbU+7cf/kd+VoMk5mt9Nzv/BVu0gdWc+gxJzESM+DJ6
iOxRMB9OgJ6PklY3ATNS858yDWqm8yDYLcv27uCvVS+kAxBvQAKJiLX6riscircLSQb1vpPlp7ss
qNUfcrF566Flt5LswfHJ+8MqyNuipcwhbGgP+RJc9du7bHnt+z1qfZfkSpX9TsOsmDYjYxHXbxF4
Y3EcLSxZ2qdsMZfgGlf7YotXhupQVT4aMlzv8XVvxePe+Hko49xns+kankEODwCdX5tt2I09Zt40
BVn4/YxxLsWDGR/HKwRCC6zPvLXpLiSkeVxNbgcfzY1MxcwhDXV4307sJ5X1+K6K5UJGxcoPuGsI
SVW5YVnN7XpXrBugIInTHh43Nn4GOQ7FdPFmcD5W9qjPl7gH8zAn52ylnZZGRzCqsrVX/elqMfGe
o6Dvbm7lklJGs0qRLaHPxJV8cc+7UDohjHzV6I8gXt7O1mxtlmbmzwshmROvm+E0/ZTEpRDILKsr
yqh3rCnfi8K/kbtdF7MN9pdWJjAUvCrrJjKzRNrZ4+Vpc/V9/zzKj9DMiJE3sDiZCR88V5tH61RH
qyXB2Y82kxC4Y2vWM0Sc4cgvdgtjYpYoZyi1iPNQjHB3zWPxjz6cUsAjsy7pr6614ThAKe/aIJnm
skbzIFRdgiWzEk86m1sBtmIYQ1vcg4y0oaKD3I7QLBsLvRNac6YsV/tvRpLZAO9QN45KDEYqXO+/
m2K07xRxRqobw4eXoi+p8qtwwTn+wmujOKbYBZUSnCsNAeEaY5MKX8zBw/LwulKvWBg3Tnit4CAZ
ffne1Y66Y7w7k0wPijO1V+ax6pssgHQYQTgLaVRu8Ts+LZTYOD0XDU6oDV2XPDyfYvQFTC8Br0pj
jN5hmgxJI+wFwx6NikxxEarwy0tCE+QmzoJo8CiG8/hNS62amYvNVXY4PK1DkEFfU3htiPjZmI39
TxMwg4F9NcqeqUyKH0CC40OizXoJCcYmeibpX0JK751ZQu3/n4mI2QjWTynNL5HRBm77rhxzeGMA
/vg8P9R1cSd3Pj1/FWMx5YJ9DxN35yCSCuxI690BaDGmL637RsKW6ormXAbe4JQYPe6J/WrHbEfn
FzkMUBx/wo3zIX/DIeNMbd5O8dAO4/BgS3MA56BRTyrqYw0f4IGZTAy+a3Dj8MLcXvwUWaTAAOJB
YoIWVlnDjPbKmOEvjgP2/2ysqIMH+rf3OxyI3vq6FmtQb2CJNcS4RPNga4aeY94HWFi0BV+m6klW
y7P7QSP10kkJPSVxevl+6dmcVSXpW5WqL4e8eV8cHDBdorVHWuS8jeVexhYf6VyL0PA35nBdf/nN
ZUUwEfYCzw9luNArLtcU6DWeMf3ztmnuV+E08YBzA0eG5thdQwQxfARRh4cAatLa/aE3DgfTct3N
bjZPdymcrjE4gupng88DBrTbYV9qzseDxw1qnY+4jELh8xDDY/zdDpjtwjIoyh0cQB5kW/aDIF8X
Vwu4FzLlVj8s4z0IBO7DWC/Uyhzo3oN0hwnkq6ApLYMt4oeyJKIIaxkaBdmGfesL3TuWLCTgqBqX
4paWTpmoxDHTv79t83PDk6PsIvazDIJAgZaXWXMNyryMeEJ02dxQm5LMvbdkz9bKDlBZRD/9/6Zo
gMejLIz1+Nf7gcixRkHhuhMKqU0encuh1DA7AuPY+eILFyrCetnPFm641a59SEnpGBR1zlU91p1d
Y50y6UnndmTn7y4Spgf/qM1OPbWmBl1mXw88oU3C2NY81m9FUFqIojZn/A8XmHMB91HI/vbR8EDm
BNgQBYKjqffMmYEZcwx+1T8KCK4lR9kDYmqzuJvxWxsYBSKeuXxrMVSAyJXTEMTHhC07fWuk/CmO
L/H4JuGJcqIRGBkxOGVn60DUksyuQBjZSGf/hUSSA4KsVhogJLf5jR99hqJOnTbSCEvbq/Qs0/hk
920h9xO7JGInMXk5VmPPEjy3aec7rWnOKEaL+6evtBJGXiaFhQaov5VLHyjpOagJsmLD0cMdxzXm
UJ/f9a18LzOBRvRKUFZetJyciwC8OqkIxj1U0xCN7bAcGjhVyFKffbn2UeACOpXOS5YX3yi00/nk
e6cBEDt3w7CukEVfrJFHJ7fpzF5OSyi3KQcscd8bxEIIbZqOLIecqEBSqiF72MwAldqfIyb3bPLn
M/NEmLpCR+fXWImcZujipy5985byIMM+tLjul2dz0xdkeHYJ6oGLeEuCA9M6fe1KYbTABxC/cOxV
rFad3LOhUTopCoRwxuseBlnJZac/I5MuQlRsUFyoU44jU38n9jgbZYyv/Z0oS9QOwH3ovxE+tMMo
wYMBDJWaeIgWsbH9u94HDvgBwckjXj00r1ynrbyVHRh50yI8Pgq+HUvJ2OxU54GxJ45eUiIQS+Rv
Jubj3tLkJkyXA9q1q1A9v4Q34Vsa8D+BdV47syQQG4BaaKwhVqBOqgM3izRAgveibIgY/0mmPz/V
l2jNEf+sT1W9Pw782Ec6HJZ+t4u9zupdSa23JCeKWkMzgBMBuHe6JhMBgvtTcu0YETqI7w9+ckYE
Q6YYgOqlmPPexT2Zb96XSvnvrN/35N4t4iZUmutsFcoVBxC3iqhKYmI+pPeBpGhAon2Np0ajnwd1
D8IlJFLvHPrSOe+hz9Eod0xBTY43X9eXwvQX6CSwQRSQ5dfV8sLd51yH8nWUmV55dGMFkHt4NSD9
VWVUUOlbv1NKCRxJsbAKx2JqE1/14ckfwd506x/Q6bwpHAro+n8K3sXnoXvB2DwBE/+gqyxEFMOa
h+a7yAMwaswCGBOAttyyD9RdExgb2VWYulKZSY03FOtcHrNELzWD5opadX1o/ZSlkAZPpeDBTlg5
DPky5g+R4NVO9/wrqaKd1561janLl8u9cjzrhxuvIIGwQqPjiroyIIJwI7byhkdb6b0VFaoz6s5l
lD6zrcyMhooGv3N6INdQKMuwjQ+2bg3U1/jQIlt4FlBmLZ4FijqzSp4z2up5IiwEg0qU6RzY3+Kv
lEOZJFf8JiuII9HkmcS+Z8PQtqVmAges1tE12Fayy1+ARymN+JcjRL1O8Xa8BP/Bf1P8VmZQeQ2Q
466oHKF2DSTI1SUhdZRwvXBr/Z4jlKP72f57tmu0Zpmk47fo6CnWWkHxcgHKQDzKYxiAelH5gis6
Q3B05OHPSmy+G4IyCYf3+0wHPpeCfUbUeXxyNorkJz2YgsjsjhegjZD8kV2sMj0wGuZLF5O+4qs6
CavkKr6xgIOrfF+QKOoN2gxzGel6yuHeKp8b9YDxWyMUZovPYNRfvrtzVCMGyc2xiSihhfgeNF/K
4/FB9iz/LL89UWWPlleCeibeUzot9MIHsgEkKA3fBYVJq5cNJ6x6lAuikMRTXp2N4ZNzWi+lWhUP
C80T+fJAXMugYkVv2p88q0aUtMC5G4BFhxcoaH01qYeY5TOZrb/HT8ywnq60uOCWbSBN5VRv56Np
vm8TEulQ/ExdlFKl5PL/gcqA4BND2qv4rryh9SfeneZb2qhGnD1e6FMu9/uiF346UaR+YDQBEbk8
XEWv10HyxUAuRnZDkydOXW3c5a7vrSVapU9lGviKKNz6idEeyrmB+ThL3mlex9wovkm1LVEdI5Cc
fDRacZQR9Sp/DaI8OSEPzAbVKM2Xqz4w5xTORMDq1SIxefWANHskLl2Uf/6epNAxPT9Kq49uULmL
S7Kv45rOpzBBPjiWK3Zx279HrVpvMtEndu8aBr1KZ7lwfpqWZcgrMfBqaC5YQCF/6aCj2w2UaAST
hxIDNh7uCbgAyW/KRfjBf9SO31oI2HdP8Et9iyoYGZOy5regAOahARi795zAx2fDRuy9uMfb785+
bz83807CvQZ/sMpeOJDVoVI1SEit7N8RWmI2NZ0T94ETBPgN267+50BsHHTW7GwKgn/to6ytyxiX
yuXCTEKJOgXBmg48xwr0dBY421JGOnY/TZy9xlowy8i19altBx9FJPEG+dlHk4lZksTQhPd/9BqD
/1Ix/+yslu9p8i057U4GvsTk0enqcL7DTxY166djyTDSj+hCXsexoLsY5I8op/VmlWnF4Tt38ZB5
AtMLCHwBiJsNs36rHxUE7iZLzhttD/rOvZVOZxqYt5RTajS5aB0lWUBKs1W64XazMOu8C2wcgut1
RQvpoxqwdxS8hRZMK5x56IF/Rb9WUuQI2sf/QC7xCsEVXsjX1/MJ/HtJTY0wIJPnUHELJURf9+dG
MHYTwos6OLXrWFQYPQgRiOBkOuQb+OzVANgqWQI41VtExFYC4x72dUNa23QDC9FIV/sddXiQSPH7
fknJOfnPW3fWUiz0QY4SdIwPkKLW0Hu51QSr8i+jcqil4E9uozXY/TC2TJQxJ03WWKqv4UmJKi+d
41GLZJcoTewg90V8JNG0wCbKa52xZOHSsZME1VkIhMAU6XuFPd0YxZWbvKrMxURLOjZdRInYujT9
siQSiMHE79LP7bP6pzE3ag3h+gG9g4b5XdcDqOXGIR3cLJ9grMBFf/B2LpO42jhNqBjWXcDXQ269
Doq8esdNkZ9+7s5JNV2wK5eBuJehy4ASKJSxfjhEoukd4ooyGPdLxuOonhCDFz6Gbst6J/hCXNUl
oxgNpeIdMybW1PbRMDHdhJ9fGY3kAVcqaFPAqKjf9GbIjVbrxWL/M6FiZ+cJcsC1AW3h2TgWpJn0
XTsGL0+TnyZGFJ3XM4WzUpQAEcnOtEdQ1tE9xrUyMlSehYIj6LSfX3VAdFL/hgpMvykGritNKS3X
mDaxcThQFzfMi/L2ll5NemIjQwiY/1h/KZvtAqoKneJ4/NWa/8f6bPRU6/7LIhXlWpKRs1F5Cg4b
b6CQYM6m1QxGF9CNxz3HELBZSGqhftghx9eI/x9C2LSq+TvKy4RAfpbP60rhn0tD/KSsciuJ5LAN
/EfRCs5AeBN5uSAACVcRgIedT9MIiuoI3lxqKDgUSMyDqOid1GozbL4dC3mQFKvreziZjAXgtI/T
3AB8VSNEyfzWe0ZHD2fldIhraoJWV8Ndq6C34sdCRpgkCZ6jY1OOZqicNVk5jzHB+GUZl7ta9KIw
0RQJKaXl+pFSWOBTmpjwB0BmVSjeY+Twp9LsBtpDHPJouwaepxSumN94iQ89i2T/x5Iu3FXcTXz3
nf7Zm9Cq31NDJELn0hjumWH/u9R/80BO6Btuh/L6T29X7VEAFXi9c/kgUUGGqSPY8j6WxbK48qNG
JX7EekzNr6TjH5snB5Ep80weFNo/CxLxKi19UHP19ChapQrW4iStxofei2C9TTLjWfou5zb/vuvN
MEI0su1QCZ7SbwuMvQe7QU7ra2azSZx//+z7o3JD1zE0s7Qg86vJOQJdo2ZB435iLZJws9xjtmjQ
/fCsHQQoZ24aRF10LUPgZdhcONsJ/b9bbSDGJYEVHr+MsS1d80tjrWycZ19Brx99yjKf8/tfBySR
KnpKuFn9MvS2lPaYhYasg27aCxwaVUGlpPzCqVEyQBzjN7dJRovvcWcuT8uRcxL8AYDNPrv/VtZy
jVc2CFfeG8i6PiOuY1CvEGLsI/e8a15/NYaDwGTNUXYKyOuxN/019tyfAOMDQrxQ505VrI7/hUUW
/4Q+ojX671+8w4IdSV/PEd/UwmWBsmY83bVXjZyGcpfyXXbXK+GezZJgVZWCHFPjo0enw3VzuBLJ
d20FGnuj8uaT8pGXLZ4ZU0bNPM45uAANHSMDcWeuVJ7jIC3qrTF16OgKMVPJUfaWOpbv523uHMvT
Ju1Pc2PExIBpE73kHEr58rWv5EGTFj30sdu9madV+dQr80z2xuK1eivyn7RUinZynRhgXfEuguhP
vt3zzT88bVufuzLJ1MeA5lyc+pxVwKL+TRedKEvMbrWdBDvgk5W7LiJKHqrlhoI4BMMHCdZj3nn+
W29OUzkeiBHxdTzm9siqBQeZCbr9rm4O/+8pOq64TmwtCzeHPjyGT6J501zQo1mQAo/71MRik9ah
h6CpTWbcXNSNYQz9ddUkh3onUkifm+bZHOCXFXdj33ychT86tFeHdfARddNBiWFGoZE857PhBqfi
6BjCqn7YmPIurMvpZ1u3OE2eacUiZPjjJ43tjtWQZt+x2Nd4SReaVpmVDbt89mR85foFxDXnHceD
Z44aT09hEnEJ40+Lhw2h/4A2Ni8K/gdyQ6a8q8f3WAPDUmd8hrQa8Jxu0p1nsiw4fhGep9IGGL3m
yuxqyb0oDMU7s0X1H0tWqLSbkNlwTIiu4r6th4fTYr40ct5DMJxHJumg1JtCAV2RBpeK5O+X77Kq
XN+9kznbgGEgWt+7xqWvK+lJbe7CZywMkyRU2esORDzxlejPO7XyQ79EnzwUqZOVyUEdGFXqP4RY
9thrbEC3zc4eEzX52+Ny3u6W2vCpod2A6kPN8hwoiRPUK3T6Lm2elCxxu9Cn4udhmIvYBs+NgWNx
wWFBip0zBxYYs0T0Ec8pPZWx8hWSuC0tvcMc2gFVsitv4EY/tGq9leR//e7gZPbXnYsliCx9Z9iE
hIw305fp3qSeyUx9ayU7ywoyQlyTUvxg9Vm1iIsQx/FN/+oOOmpCHrdTVy2ouduSyQ/DR0oNMxuW
hmNRaX/1wOQ1cGQworWZqrsb+qFKK1MGfUP3+2Qsvp/BcWvzVmipo5kd+ucSeYNRkt8sS1PL3t9r
y163Bj3/YcYcFan9MS+Pl2yPahEt6znLgVR4CvPtucXX1w951acL1pCQnUT9wbwf5GcIeS8bcrt+
Bk4M6LSTxoPpUDPclP/B2gt+ywsyfEXBxprvFpOhN629nJ5+DG8xflyCKS0VcYWN5uQ/01ODCM8V
XQhC10OJhZxOayvRcOe2Qf0a+zJ4hYK22DT1tMI1hEXhvVLKZqciukHu+1YK2qr+7JBXu3gTEk7U
CbL9N/Fs+XunA63fLx+1McIXv1a2gOxuYQqI6pMmAzmOaCTXTOWQbgrn69dv+ZnI6Wq8dqaoa2a9
2TA3q3rzFX6sEihPKcuUH7SdPn1k4RPzHRKC//4JvhH30ahi5NhOBJQO/LvNLc/MZwHB2GuDGSsc
hvmKKQEQYselEjLAg7VcEeEw/gQyNxxhlR+hkeiJTp0Sd6yN76mo4rKY9VPO4EixN5n+8aG9y7hr
AE6bV8NYjnVI3ncPzpyXXMLGaz/7mvUrGWMIL1QlodLWOXmw9g/aDWW4+FwhW4SAY7X109+tx2d9
9gv/FilIH/k/wfinittCc+iQYjlkquYQ/EWUaNXAYVNNXGF+wfkRNdfOze0dGTGqTnmDJ6f8/oh2
q9u10fdU4VDmuzkxtPZAnZN6eYw5kOdUaigkO/D2xj2VkPS/YBY4ebDL+NRgR71QK9OzjQ/JYyUM
WtC6nHSMvDoUYQ3UzCN59MIxplApIAm0IdvjljsCD8wdgIHNvcKGd/vJaYlDxW+J31/RHAgO+Rh4
ylPjMQ8/MSMGgILbgLu5vrLIAE+zVOPI+ubNzXiLkGW5XCS4vtgJjRW1fsPg7i91pNN02MxJFZzg
WEGNPuSIpSiiBjqgn4leHref7hPMSQ/YCRU6yeYfPaVsidJ5x7V/d0jZtsAwQzW5+gSPggUgnhK4
nNUmTMCFVVUGxx+eIznlbo0dCDaLiHnkaobaahr+lEwQPs6cCq8eW1Td/hH+9ciwQO6ES+uK4tHl
PA0qOupGwD6lYexKN64TB9xQDjOzAlvs5qSKk0ZSNNkvCsl7z/Zn/I4i3+v3540GKu2BqzDG/1R1
CInyqf0R3IoakL4mnwklUIQpHPzAS1qw/uMe3Z7gQ5Bsg8UqfZXW7A4sJHPMoDiowTLcI6uU0oXg
oEYhgCvhUdXywrI6X+m0k2MP/p3wr3O0PiiqR/Cn3S9pqV7QetOTZsE6C7UmP3PZfrQjvI9rHqfh
CZZKbiTsM4Pnd/PuUsY3ZaN3qrW8Zavcnl6hRWsEyIi84ijIV/p+m5l3YSfYX+HC57w6SpwDOY43
9UHrR9lSTa2Jfwn6aaTlSOjVUN8Rgb5Ho5/XoWkiSgxejvZ/pmDKkM3q8cI05qvx6caFygqT3DSk
xJ6oDUsS3baJx/cnoOcjkxgJ8cP7ewwPqGHSA8nHGGNnCEzecOu9eVHdeQ0vlBV0pIFN32xQUfIR
3yZQIhEdoWhDMlNC/70N3k1PgMtKCzxJUgp4qbp/SGcpLUFoPxrE1VGMW7Zj7U46DNF+1FCImNSI
ulK8wrisnt+5ynXW76w6sOy/wLCZm/Rckk9pZ+QdndcLWiDSQ85Oy5G+ldMdhF6MC6Jdsh31d2SV
OAthN8fALZqIroxrno7wJbHMbHNH9vOe7RnyQHFMmw+l6u/Xyl2ZV71UIi1vylexUKj0tWNIyB19
P5qh38ZA5x/MNVcbEoC+MNsijeM49440lHrbfry2uDzJUqHNTG8/BdNaeadPnGMMXSnW54bkgk4W
O+1hBiYyMf3pAK3nY/U7ZzFzNPE57y/audUJwmnqKr/Gd6feNbtsTXBL6xUYCmhQ7Ga7Eg0MrGO0
HNtetTZjXbKfyYkpy4zUsQB3K+lXQ3JE6+EYRRvAIfXII206tUDpvjW2pbQdLkpX18PnDi8Wet2e
rzCJ8+nj/MZAe3gOLRtj+JvAoF1T9HJpfxvrSHADOq0RjLC09oAJ2BjkMDMcezdNGc6PmDKpFyJC
FqlZ0+NKwKugqhSpkX5nKQqxiKJs+pEG38WEuH6ZqK6lNT7G4ZYjpLEgd89gLofi94uaJIIFzZYH
rzmIUkKfYve5jS37uHpecrpnBPcmBXLk67VKpjL/voxWLT3H5KRIsy6hp7kCfYhh9GcTQ4x787fi
oZ6yAPX8D8Zw1XAcxSbeGc7RSzK7axqvH1+Sce3msZdTO6ReGCGf8YQhmZZ+YKUGI3aUfiL5D1/E
sPJ8AHYzJ8NpkWRgTMj+/hlOoeqMzu2iGgZiEtdfmxDNE0AUKihB+uO3Hodowu7aIukDnSvdvfJM
+1FSLrGCki0g3wrUltRCYPVQOjd7wMyHxqaMMz8KZ3yhc+LHcr2KsuH/mQQJ5VLny0nYt9RmHoEC
0OAjEGPbMW2mTh2OeDIz/zt0J9G+Vke3KMyJDABQYkJq7epu02oem6V2et4hfUzNzVnKiOKucUsS
t7qKyLyjPpQKKk8sPOKj2ggYkW31tR20H7csqFkNvJ34pUaMUJTSl1NWWR1cDEHJzVGDOXUQWfi9
ZVQ4t4J9JwE/0J9khvmWJw9Yl9kzLjnbsP6y30zaHReRVlUlGc6fj7aPhp9Tu4aqh5qEuhDM/DAI
RCrvFmqEuXO2f7UwWua6l/5K9wrV6R+iOhTGT/svs2OhaAokSM0NCdmAWOS+MnsUjVbTW72A+bJY
3f3EMjqSBW1+hP8ul22EQZnS60FjhPLzfK6emRtl52ssh33bEDlDNF2gsYqlwlFncVb6hz1mb2B2
1e9dgEFtyNEaoY0xws+xwMpag/i5AAsA+2SZw4KRyGFcOr/95kZFwMDlTX8E5sOT/ydT6fV8LuGj
I6CuZHQu3r0drvMuJtYt0AMt26vRKsVz8Fh9J0qq9oUTV+gRT2+HfQBlSeDynSd5+Zegx/+qM5qE
0Bdlx50biXvn+PKwoJex0p1XhlQ2KlUnM85RJ1qgxZTdqMGVzgChf8SflVfT2m/T1go+tZo8yu4/
ApVxQuTgCwfqMBBQmAEYwQfovq2A2n7mPS5KZBvSV6vqhxu/hBB5hFgUU5Kfj1ihGH5Ir2xqcIj3
PB1P5jwan5R73oo1RtDH87E0vDR0OhNH1/BeMJ7NW3WWF1K0dLyxBFRZBj1RW0G/S1/nEvUGuqY7
Aw6q119LUaasMf9DKpOYr4JHLmFaxqQsqli+hAVuSL6dzSfStlKBoQ01fSWrMpwl6xmkBl5BUUTT
OzDW3mUL92+vjCT3vqvMQOuO11KiTWyMJNqw0lJH+QIqpnmDPQJ0CK3oSK4RvV4yqzmfojH8qNYT
ewDbzZpWd5Gjol5JvqcoMoxtkO+tEqJr/7+S1HBPkY16WoOhnlib+Qs8oSY1UVT0YbwMhKADBjvG
0GehX0gUQl/W4du35ynLGmQd5AtsV5OyMlAgXJhmuaJMrE/xXs5qpdpJtXu15MuYOSTmqLk+NOZX
uS8LWrWnaKkXQbZdfND6647AiuNZHy7kQthjUe9ru7PUU+M9wlv9+IHW14GNXnqk8eG2PoMzY0kO
X0VoqWpgSKk4gm8gjrYNjRkBB6ApS715xpBvW9qjHXFUX9RPc8qyhJ7sATkab6j/NGHKqEicXXoi
jyLp2nBe1rxbWIXtPUAI6i+ss78XFR0iODTtZW2P+YQoTNrea6enXyJMzXD+On1e4DTY3tEx8KYZ
TSthXUSvEFc6aszKW7lHtVl0RB4KaTbUJv/GDzQxeOTBIXIG2KC4XFx8VXzyao+RFpQOFMLm9fzb
2AxvGG+UU7jP7wICW9BAASYqa0y6CgxrNcLr6AVkrfwSJAob2Lon93LFeav+/21YHF080C1MswDK
jmoSM/Oudpc10/ahQy9/jOG0P5j4dvyyaEbiPyzKW6seT2ffgdxm6zQCGj2km7V9Efd/btSEToVb
N2fj2oEmZlyx1N2ttfEz3eSeh4BUpF2n+KMjKsdOmC+fVvZJxT+MUTy8GfZtEiI+g42a3dvHWDr4
ZjmF6NNrYiab6Z0eL/+G7AJaNZPTWGoeBnVJZ+5tUjRmJqVN2EGoN9v5sfPXV6z/SgkRatoUCS4l
Ow+DbNWr7Bmnpe61WTs0kJN8bzkp1IUpzsSgKqSXXb1UDHd+PzqPfD3IAkHlTGQrp2FeqLQZaDoT
mwunrp0LE7waW6oAfDqBIPVRyA50j6vNv1mNL1g+jQFB2qZ+IurgMHJo4Jch1cEaJOkjT7OYX13u
4T/2JI2wzLnDgUh1Z27/bctVrnvlxl2sgnsNPaI5NIngb6oG0lr0eZ/gse0O/cTQiYcGA/n+EUL0
AJp/zMlu35KQdnztX+PNbDtJJP1+rKg00AGDhIQqya47oMn9d45ACOFFXbixXNEy8+eGDxpvQv0R
MRyUtoIoYDCb17QoOpsg4k+NBG/gVAni7RkyjVrGXwv95yN6YkALuTrYU2bQxHgx3bZDB2VvEqFX
Qrfigw2fgvBuEFecsInRuTNzHuUWMfTj0xOnD4QzddHkTKic3momWSz3pv4sOz+QMUPx3ulpmFHC
lxp9Zm6Yp0R0ECv93f+b80qOr+dodxXfthQ9wcOiCXZwBqJwbyBL71zWTMzFCAYITyOnsgYtMZJ8
p100UbGmDPMnpzAn70X7bkbX9knGC1bIcqsHUeqsb6fB+XiGxwdDwslwTleqGUbMgSi1dVRi779D
Rw1zBxLqS+jnUGj4+JwOI08YDfJFpXcgknTjATrO4Np4qZrCaq/cAwoe3AKNdby7O3jLgc9BUo9a
bepGC3+b2+cZwgrHM2UCp9ooO29kYL9jhqHXRDrhA1mXbxU6Fi5H3LVOxkRkMcQxgsBLmQTA8uJ9
5EoVrWwdowlQPXDp3DliXI1NCMHud3nJ+PEVt2Shosnww60edBYoVb1mONuHJ2XSNTWz2Unr/ZFz
aZeBD/Y90C9Ox7wfKfuyPXbBAqyOfpfbkLmBNX/N58Q2v+sfBD0CQCSSn5MIoQfDhqGnjwqspPxS
z0jcNIkcvd1w8IU4ehA4tQbIJh2NSSDwrLcKEY7p/6v9Wnd4TflPpK2Ic+xTC7EgfOy7VExjIa/z
8HsqweQYgMBqXpBOt3ZHvL2sRMDg0GhoCLz0LgpztVjIW+RgHzZLrI5ILcWe1x2e6qBeJxD4h5Iw
BERCR10PBAPdTWo8/FrEa9Wt/AbXWdu/GPfEi4ebD0dSQPWFlc8l/1Y8lhfVTqBbAOOvbrLz61kN
IDSbAtZiVKuf37/8LgqBIo6TK2TirvUgdjWG4fuICP9fCqmmiqVEM0M5WeYKr3J77m/JSY2vSSYj
L89gucLDCFq6VLc14zEH9VUuNX5MTurqu5Uo/f0Bp620scf0cwq5/4P//vHMscPnjvLoYmw2CNmw
p2TbFcRjdmv0r+hIzNhX+tLxX81tvjJq64rDC8FNCb3O9kSKOjmuArtL6tzXUgT4I2eeToHORnV8
8nRq4S4cejul4AyO8DUAwX+JTs3VbKbB4QkJR7npZMdyXlVcdPlC29lh80shByst8CHSQH54yp0t
WjYXJJQfJxYpS8rInHnPh4uefFLnn0j6wHSp9TUQmLgQVZBuSgg5xJdDi0Qq+2LeLoGijwo8mgs3
W62QHHJNS5mFLUk9LsB2EC1wZuywlJc7YVDLZJfCFvM71TZw9OVK7m2mpIiYxVONEnxz0uRPmpvB
Q9amRCZoT6EwCNy3CKTB3dXSQp5LDvPzJDHOOPVuyDpdiOsNxLn9+E4sOI5kITSdj2+uXeAsmZu1
RXIEKnItbuodOHpQClWZrSCUvaP3aME2wl8qX0WbPABNsSDFkRvxKCpugFB3k1h6F9eB6l/+w1YG
+NxkPyakHAuArx7pVgRkiYXg0UJpcQzoz9m6I3lChf2uQNMbzsYNEf0TLoH6oVRc/hcXS0o35NqV
jQ4BJxKhPlxyhtZKP5AWvgkxhj2MhN83OMtPaGKBpZD7PP7U0HIYMUofApEAuQ02iQZNHODNuKm5
YaPDxUhwAaFy5IsNtvRte5b5pg1WtApmIjB3JVBAvFN32cQprgR260uUU+zz95g9H7QSltIA4tuV
UYw4gFatpXlmRdxwHCQDk6/rMbC8hz9pttqUL+WNTHYgINp7y1pRkUtp//aaRHdAZ+HRdDX9jaCr
gl9ampC7FLpGMWQH3ZUEsQ0vFqBA/X6jx+cyAolb/SAUdfFb77hG/A4pzIgIZx81jOvS5EhL/2u1
hfUcSU7jiMsOQJZYEEcjhtr9xuR0oV65xtgPrOkFlA4zfVyQvddDI7IwEDMRnK4w1mmIsyRIgkXz
Gfcsz0euazXarMfzRlm4peZpv0K7+78NlKDzhgI78c1kauC2duMfl2H8W28QZtw5TrzMEKlykPnr
bpFmqYCKy8ChPRjoBNR/+wnsPG1xCkRtfU2NHSjq3ii9wNEhA1YiqSS/Zu8eJGs9su/LYl6W3c9N
itd+W8ddmvpD1OAqd4aH3V6Fy6ve1jnZsdAcWQMA0el1UfEOmWk2n0kPg+kQrBujq83EcO1CSDIo
402/wPCFrGgSG6PKNH70LZhXZiiK0/v9CMm/shJcHfLZbluoH5eBkWgA55y+04J2nQFvGWJ2cq5L
9Ma+vl63lxenvGdA0WdwUcF6Yo//nPOeOXHj/9aEf3fCOKa3hD2wNRt3fSaCN7uAl3lkSkE+DRwe
sumMD1ZCw80Ds/d60ZLb1nUgvrAvofq0m96n1kzC3rPrZTkL8F//B2XrEuTJVeonfy/RsqJl1oIs
QR0wZO19ypxBGTpjdwtg7H6Salp7oylQ/YGzTgqTHe92CPrmu9CW6O9ejpGEgL6YSJcILLBAr2Wf
BDdt1ONYaYxSlX1jX2p92VdgyGr62qyI93ZF4et188sCJrpDT2NphPyYbSSMeXzYD7WYuFp5PcZQ
CSTIzNhqpOSHnLU4XBJxNjhHzsVk0IpVoibnOpX4qaMEW9VOB6gwx/1XYoHppX8GyyOYWx0yhfal
2NSVpr8o9sEqGPrN9/tczjvyX+ZVovDBNHySTtTgDD+7oRXe1vC+ln3qiRw+fLmMxCj5BQ+6lH09
bECf7+sFkPthfn+NeWS03tp0PeHFDiT8VT/yApvZTNwQGTf55cgSlVdZLqlyNe/csWeSh20MEyfK
9LU3GO+rX0NNQlJ5YHHP7UpUAOer1OLl3+qnL9+K40/TFhQBcvp8ZPp9SnwRsAnJ0S+8ADXfFt5V
b2z1HDYNgwpN7g7EtVQ3YEqAAFQrXJEkC/8FO3e677en5pSnjoJ5AcoiH6V04kh1BsRbMNzGI8gS
uDqHMpHYiRtQIrqM7DGdTei3Nqcep9L0SgRwUNj8w8r18X7k5usenPGeD17BcjIOGKRLYJDYiUSZ
O+IH+5Y0P98MlOiyXNTOf76a3Klp8KnI7J67Dle6kJ9Ws86zblIa5DEQcjXqEfPGJJQp/Wj1+VrE
Oqek2yKNGalSdVJo2KPFj8EzJkU8+3w9ZafjJ0plv0Jnyvzsm7pwjBzPg4CncTxeryoPmn4YPHYj
KdTmQRZeIDY9Yw9jvnxLAjNHXqQ19j1aP5m8Z9Gfri28c/7mQUr5UGtE95RdF3EljS5Oec/QPuoE
OpbH7mcF094pqCiXLPoolGc+TGtZf19qL470MjtwiqQZ/GWNl4IzP4qhh/V1VvXO/y6jV/1ikq9V
ah8s88YFshuwaboWrUeiIaf6sXJABA0B8U+I5KY/GRNHBGxyvPi2MlCyGJtIfn8+Uw7YtfEnXfYr
XeNOYJ+L+NzcVJ/7BWjtur3VEudm+KaU2RvWaWUaJSlQYGVR6Nr7WptSAvw1ZdwcrNSmPDCIAG9A
1N6dISqY87RQpdCuR9Wd4yIS+aYPA6iUSfg7XWjzglbGqou/LUNgAujL1yZ0E409Tp5i329q55J+
EC+m4vtaU2CcKGmusxFUxIcaOUC+gFux8kwC2zl22FHaNx4veIm+FqgaoPstRGPxVb/kJHP2Ops2
6RUXeSEYir6lF5dKAIWDiEwsU4NVqrzKRBLP04ohAtGvlCxvy/sSLmrgb9CDNwjhGthvyWueoQwH
LZj50LtxVgRPoIx9Fk/Wp2xYivNXZL6PI13WLxLxiEESgcOBdpVTER9bh01GnYq74R4zhgPCIPB5
NtiZi3zfHNT8B+/DFNKTbVjsfqOggGrDIbm9KZSigdfu5Rxqs4DQOPwZJdHQaAcxkErNXVHcEW2p
HPBo0xLlWT7akJtUWHkMmBi6XHJ4o1MloWSxyiENe6WH4DEAF9/PqBV14XZ9t3xih8Kq5czYRCSr
9C4cktoBeQAuZEL76h4kywQ5AhDpcCZrI3ts0GGgSmTu2qGVlobTnClGV0u2DZKJy6nXIKAab22O
qSIT58FLJtgsZ5veM53UB77O6jMKuOmx4kEb2WH7i1SIL5k8NkUM+ENx4C/Vp4RdD9MEKPvZiGch
pZZHl6+wmIKb0r0x7egL569iEffGjUXk6391158dx9hx9+S46eA/fJsQYRIMiUVFRNRIHYwlEu9Q
kcRpYjnbtz3qBs8lIvXev/sC1JNx3ZQSOr2x8K4sNtSCT+mxO+8IeKYNlMHTFIwBMCIK6hBdUqVH
YnYaGyFtPrhsy3Ll+OzCUEzszRf6ijVJpqaRFy2jNZL0xA/lGi7QGEY0PWCwTVL/xstyIxt+jQC9
9YJKJq150Y8R3vwRjSMX6hsXu2C90vS9ea2bXjPg6StHV2GEFQLYXjh+AWkoizaCynJJNpspZkex
JbBcG2TZ87Ah1ZNKK2wHixNDPwdhfmVyBR9tcVaUNKYVzB7t+fHuck5e1p1epP0VOt5pl3d+p7PO
r5us4/1VK2mom2KhIyw9/ho7QjzFMw4ESCp8XER987/mv5dRzBxWqbMZcBA1MPMLxQlufOCyKZFE
Ps2H13JHQbDGXHpnfr6WEbUkz5NPKP99dXUzY1mXhH6aCAefc8L42FCyYhvt4uXnJEE/39Co1DSP
tsqOPlHDeJAXMpJx4MIiuMcWiieSVk1x4d0g1njZVidVFr7ufZPHK+PEEf3CuUJlbpOROoSgsPH6
jH/Q2YysctJvCczIxcrPssKKfWTztjtv5cWj7Nz1WkZ9KyCkT4kVdgl6mhKjt27dD1s9HBWd1Rxg
l9Q7lkWbSfeTTAFNcDWUZUNadvbeP7/MaJoJTRccyV6NF5ka/QuVFBdSX17mYOoowOFCWIobx5et
9Atyq05bQeOoLDcNNfXYqcb8NnIjGXX4KkHd3C+TGyaw1BuTvtJHRYcwh92A24d+se+udRa0CbMs
CF/iRvTpOY2GRFyKKpMyq8q/vSn9YIgC12qw+h9VMycB7iJADPAkcaM3gXFbeC/jj0/d3S8pBQZa
N/j/oXC9iILNNEsVkKZ3/GNQlniPA/Z5jMPpf5Yc5pwGR+zQ0ISM+YuLElj4t+owoW/VEgjiEXPj
zEn+1rRcFpZkw6WeJZBn21K23RG2pG7W0pgmKdNhWy4oCjSFJkA8Lhcr1C2b7OfiAMtB3EiVlQGC
CTvxvyIfJ8w5snd+L8iAVH4H+82ZctCx/evrTbc5N+Gxa5xVG+Ck5Kln9zYh8/fklVBh5vf/FloH
9uMVKMvW95cIfq/eeLLiu6vBYm+nmC5gwoTeu1zrMAgOKO6MXrUIrsjCOCnzpFoa6xnr6COJuimP
agIj/fOcwOVMQZoq4AZDa0DKkgazU9BjwHvZweI3pEFkzK+tL9LR8lIxdkrsp5NMgG0ik6RlEGnr
wHR8EudTiaZDGRhJrLoD+hF2rlWoWGV+kJLrZYumIQSQHeDoKd3KejB4zusSZNmPR6L7Y3n03Ogm
8ZlyaPjnoVS8klhocl8BOYqfPCSbXsOVwNHMc326xXg7xQjR+nwDZ3Vlh15/pR2r9EjFMuTmEbJO
+xk8UeQelTrXuAsb2f6UDLO4Qca29+lbEHh2tB0I8s/8DJsmlEwCNArot0x0MeTKaK7zrYP3K4bl
2MVEp59q+D3QmlhUk24NFqjYSak2iWmecW8rs5Mu4VU27i5xA5M6F7gtJRORRkI+Dtk12By5AMcN
rRVJz4zpMHGKC56UvZ54b3cLzBdWUoabfzr+CWHDN+GsDrSMDPLBpIL1uqnpTtjmTR37A+UvV1bu
ww2cRjULrlQ75nlXhlVK1hc8KFZjVzBBveK7eU++4kHcblZmCZ8xsglQEUXh2sqq1I4xT1N4Zd1z
tVrmVApx5bWK0mLKfBd6Igz1P0VWp2ljN3D8R7PRjLS3hlhhjQqqj3xogQc1sKzcqlhiXtm5gOPk
2IZxfJvt8u8wS4JezN1hy7mnHZTBsFgcxLniKsdqBRu0C0XUBr5wZ5tDZ9J+h6oBIaXn+50jif4A
lXVojPrYc0kvC8ePmBJsRz03qh1rKBhSO5kucBbJeKdyqBnWZ9X9NUOIjvty6OS6nh2I2kP9qIC7
lpd/9Rg6iJki9sW7Vj6FJhLlEwoCkIBm7V6u3QKENOiMKxX4Rj4J0BynaraNQ9e9bLYC2RtYSzur
yRuFh+23PgCdsdg1EeZlbr3Mj04WwTsC1WJpAmxwTLr0SBC+Hc17APly6KN2rQ1wewBtYD+ghmof
ctZ8+tAhg2MiPr3+5L2GWetxXw7bsa5IXqksvVgudzkNzeGp06tG4tqgsY3h1izUJ3JyROFAzg+D
avbFxNHiJfmb1JO1IaEuaRJ7rdOqDvZx+p61rKLBEgYlbCWcs6iPag2FUZi31JJypL+jY112prAW
ZXDVP6dKLn5ho9d+l3nT4kcXYq0OFQQRyeALBxKBYJBqp3DlH9Lh0ZVVreCJZhHL3QPD0uslFQXK
iEqcqv3BOG9EM347y9or3ZUE035InvMPk8RDHRnQB7ShSLucyRyzZHj9DX8WJmQR4CDXadzY/Mzq
w95tKD7cVDE4qNmPAD0lspD10/tEq9dM5WbMXz++XqTMFNsP4hWObANAPkYNSwZSxTVl6OH7Asqh
xHsNNjRdLST0vE1meai8qqd0xJA+dzF/z96cNskCfQKaBYa79Fu3LY5qpU4ob0gYgt6ceN9P6qjQ
gcm/K8jB4nUPnE0O8ljogxx2+R+bsqJB1Lld6ax8ceNlgz2emetc4VdXZ1c7C0gjUiQAyoVxTd20
Tp+XUB6PNBt4JKL4evbudAeK/4evRzBLoe/jTXB5oC1ABT+vL5TJHA3buV2kcEIRJIdpvlUANLkE
dNvNzrSJlIi8tn+ufC3Ef5ygHH0J/2qutvq7F0Gju8i8Oeal5AiG7XSme1Jj90PpeWIfC7CdKylt
QAzRNh/j+VAbVISi9KLaAZdq+xtk4+/YKTBKr4cns9ZQvsjCaBN8d17RciRrxJ1/TjUMYhUae7jR
AtojPMa5or7CoRDYgChk6xyIdVNO5USdJavsVJzOPHM162V4q2aDvONPa3D9K2rUvyp3kFbGquud
ZmhOqx9iQZSyfU50iaoYqjjGiL8OM1FewNQlInctyLhvrnt7Mge9l+A7I0zPvR52zsW3bvdqZc3u
bOu6l7SH2imQCYmtmpPdQaBJsWKr1EnDRc0Z6sVFsc7lbscjRAHO2eAphnuu0tfmksEahO74JMPT
tpsQEHl+pV+SDVbkYpMv+TsOMneuoCaURdAomhviib2JpbliH0ohNBaLtJvWX1hng0tyrLsORoHk
2Ilv/QBswOqS/z7r6893w8VOLOPJxwDj7VVmJ05vceWulJF3Ezq63wNq5YfwdKaDEAQuVfywXOrb
l0pNereSDnrR9RmUWzgiM9o2y6JYmm66KXchk2m+PbrtS76KBzI/J6BiYUnS0XXjz66ga+Xzipfi
QARRnu0BcGhOhV7R9EBnWrW12LcaP0vsndqzaeruR7KHfEIYvsFHgqgro6rSrQktnrCQmATo5A8N
m1aeHixPMRnKgpXcCDb7sLyteFjxCB2L9mKhQMdtuEvlFVuZvKnkiZjpY7Du2sqG6BHZB/C1kaUb
gt2KZzXtSdGg6/A6JLnavpLvQL4xmSp4U8Nw42kFLLLUWpiWDENyfLrJESH4FYbwhtPvV64eN5+4
ods0T+FBmobeeJ2GsOsKABv4ST88a0eiiTZJeTodr1EzDDbUUyxfZeG1utlUz5wrVueQG+j9oMMn
VLUOROB4ZyEDGOhv8xJSJ7r8OhSsFERpFvhdE3Ni0fWaQ+lmYPDC4ZWsGdkWOLspkWY4f9A5CUDR
sqADHdR079gcphhNPZ34Z6DPsoMnaX1Gx3GMeiFDSAilNc/nSKFQcdMgXtA2K5T8xpwKlGf86SPY
0QS1rABDYzVzME7z79+bBMVQISAe+gSEcirKXiOybrZgYDS9Pti/+s9pvRAbKTf3t/oFCzO+4RNA
Z6VcZOCEV3OmhS7u8CmTflEvqqiS+dPYES1ym7fGWQoV8Ezn6WupcIFhB7Dm6/verq1w1tkUwhzp
m7HCkG/S0lpCplI2Lx9IP3rcRrev1IQKOUdwNoGk5mOO6TU+JgLhOGyRlRkTmJZebwYQZiPuKN/8
Qiz//22x/Vt4lgf9Bh0ELjYoY87CsshugIIAitx5eeXbj7flJkRnzcmReVShntnF9rx/89b7ge+d
cjJzneh24Q5x4hypXnoDFR6CTJpFBAOJCnARnx+U/VHf+jKhogkBlZ+dJNshVw7CiyUU3UDi4o9i
HNf4MzS3x1va+sYy+uH9SKGw/zI+s+k3PcBlQUMyjP0ao25V5tkXAhOBiBPEnCWwsHO3MLHdCwwV
UM50XJcThAv5ib0DgOQQXT1mmh2O4jCDXRhQoWz3WjCCM1X/1zL03P8LonJwfn0i1fLqy8fm8Iq0
+8/HpkmZKJ5zBm9fswQ35roEGTT5h1sR1mO0gDzRxYpHR1eTuxP7YpylkPUVR1UHGVMIxEsvrHZT
FrmrPAj/AMnbu48nasik984wZIsD+qeltLCQ/R1Mexdwy6WaIyg69LJCfDegQn7o6VPXNFgRlCLQ
BrE8+x24t23+ARZMX2SnM50RG3DnKYkBAWjzvmgK1CHzYKKxxNxET7deSQUj0UqTemOwX9Ilud4V
M+9UsdqdTfi5C5zX3JONagicjTpIwNs8rezO1uZYk3sPgMOFeRYS8vp+MAp2MfPIJwtUnSL1sxZM
uTCThDcA0gAPNptoPTm0M+n03q6JMS6mnugGFXQXW18O/KDPCTuh1B6mQPTqqxyW1xf5zw6SaWkU
+xmB8962cNVhDw6VxhTLVC0XAvKxS963kWgmWLB6o+OCdKLMfpKfOW5FV/ebTIGGEuaL0rynZz6T
6WNJ1TehcfRk9X528D4drrX+Qc8V0OOELZ6Qhb6FdXMi0AmCvZiKr25aA5MBNDNYW4yCHDjNGKqt
RcWPnW1icQO+6qTD37A2PJRfj+FciapCMeSAA5BtH5Amjk9rySNoljyP788MG8I4rW4d59LoKFq4
e4hPImkNTfac5CufDWQEnsz5Dt39A5JSFxGjeAWzzRTfQtc7McatEBytciMqopSL3KkHNSRO2CyZ
MK8ff/lpHTf7B/vhaJWySqfGj54Enhfvb2ncH9M5LbkZY5ZvICRgzSpqnmMn6KyPDre2CTA1zmrh
+GNggnBRKqRrf+wP3oc952lacKrFdIUGoPNecU6BUrKXkMkKB8SezKOKsH5TS4J+qANrTqGw+OOb
f8pW+T0RYTHJ3wQtSZR97I8Bm/BsobeuaY/stQZzmJe9YdzadkNCfgXDJ+8/K2/tI7NxPmCBfn6c
L33UXz67Ib8duN3iTVH6vXESnRViZPFZh1WZGCMEphz5ETNPCg6ntEDEM8cF1aFuiQ7OPUf06ePV
8NrvJZGJhH6xLef69RL/bK5xCUW8Q4CTxP5TzFE0ym1pc9F0mwg89Ku9+DdrPQCeKJi3ruOXefzT
6o6oBtM33V8X8Lro6GDKTckjhAOaj8OZ/FJKWNXyd3O613yqJJFMTbaoc7260DeztysTvVdiopsu
SXycWi4YEMrZ3eH0uoxvdiaWBjf42sGQ5+9SZADIkhrrby0cI0FZoRZB2MFbTU3O4oRamZHao6bF
oX6lAJrVlO2QAe8om3R8PInHuK/jrrBg8L2EmgWgUVQBuhkZUYz4V2FV4d10906yXySOOlbViCPv
ingdcytypqOHRKkQ8J+gv9T7ToUQTEJOXqHOqTERWgYSds8h+Vj79iVDiJ1/tWqOIipVuTHyxvlI
+VF3fZ386w1cBVdKOdmEjtm3Yyc6NyO1ucimqmXvjHQzvRqTVkKFpMInQODt731NSm0B54w3DnlU
w4S6pYDVirKJe1XO5xAQVHd8r8ZrJxatoG1OHC8SIJGUHxZsDGSjjoSY7UMW/Nrv5WBVQM42Oqby
3v/9PCYJAzXqq8IVYATapHfg8D5vvcOA/R82GOAvrTJJo1muW2sTpyn6dC58AyBPjBIdgSBLtFAy
NPHccXY4D3zGcT4R0acVL91C5IlCaN0+wWPbJ2QpmYv22P/EDxblz8AxsLsbAwIvhIu3eAGmaXk/
GcBYefXyGjVRaS8GQs+LNV5h/Ywknw8gXw7+b9t9reRMl08/F8BS4esbn+YOleHiUyV9Tnq/4m05
lI8DYVOyu68lbdeixixpL95QDRs77wuixg7M2RCdAC3V1BhwxGeOfP41rWxWEGyhKdNvUwZWOmtR
4gf8HOq7F9dBiLcoGs8oN/ElVhAi+WvtAZmCDMftxkOm/c3+P+xLTP32TsIkKywV+nKioB9i4Phc
vKJ6XiNYy0boQ7SLFFKYq7qhlTs238m+SkmZobIxFMt8eGGYdhnWOUovMdz94hIk4PguwIJST9Ej
sf2Z1ubmT8pZ/9riuKKg5jEYESO+/MQfP/hcsMMKvPz8HVWMsD0Lv0rZp7TJzsSnCPI2Kn1LR0Cl
Ww7kVIlAAFLO9Yg9pF7n+jhTBzmWpHi5OOa4NRu2A6+Yp4yKT+Yxol8HphB1IM18jtfp/ck1FSCO
UKAZlHIwuyj/K8STY12pWiTsWK428v7bW9gC/6AnzWEHqy4dgZS1xLBnIBGj7pY2A9hGZ0Ucqcnm
ili6crzYVNbSbxV5axwJFUJGsCtfHuNJmGfZzDYSYwoX7+01gdqtVWkdtuz3pC29jaaAvQryYRb1
28GxFXdKewt5Wgj6SJSaz95UpSiWwqhX94GdCtHARw9e3NFAdgdSUNvLp3T4aFG6U/8JAz4XYYxC
xaKzqyZH5snb688brqPBwjnLDcMHfQkEZffVwrfA77jqElj7UOhx6xx7dkUEIcybzdikopeyU0Uq
quumZLlFtoYeF3fbgi4MZuZ4pzi4KIGftqMaAbdXBPcOKar0+NnHSthPCV1kY+MX632Q78vqinFT
Xdk50GTsZCeITl+70YoNNb4gfOdaIS0QL9YV1nQ+zWgoV/2nzLwsfgzsp0DXE1ZxkyQsQD4b231B
jYQWBXflkpPBWyr8v8SDNnoLOmLM3v5Oou0TKqwHTdh1JCVj3pc4C4PK6p+HF6gFQEFgIwrGdEe5
qU9+G+mwk87TTNNvwUUCGidRKW2TS7egTl9SX3h8enACfwaXkZ1uIKGRXxmAZJFG4XFYk6CrRybS
TQHAjKLLhfgm+GUz7R/Cp3GUR3k+ur8COdhv8PdImlndnNe6P6GMJjmxS6US7VptFcv79bSgc0yP
DwIL5ok9IvrjsmIHA0sKZkdYnDNa3c70jh/RwmEStUvf/1VYAKU4ClkpPgQ3H8HJMwfxmZ8sbhVW
QSOwODfdOzdmewkA6dRlf5Y2VkgfXVtDXGjyLbzYA2jZ99SdsbdnqHkaA7p2x74cTOCiBaUDWGGa
3u4Hg/jX7ATH96NQ2+HoSORstOTr1xne+/p/3jXVgwXhuXbIMbO3oo7cK01oR2bNdSADTjTqTzhZ
xjl9dixr6SOwqHYe3obbRE2EKyBEUmAfNYQoc+Nws/3roK5i5M1+QUEtabPj1/tdvnR6luscZjU9
QK0OMEKfKjdPb2c7pDGZ7XKyDjKP/f0e8GUrto+6C6ZpGGpOK93hLXM5NTxsgd8WZwhsrY6c21of
dogcdExTLTeaG5pPo7zKf1lBIhVyxqEFnQn+ok5FUxOKRZ9k851YCMm073vJAsI7sG5tnRHUBYP2
JYsXbDGkHxKrHEQ8ojZ4m0KZIIpquGvxA5WJ6qVcH1GQae0BKHX6WXz6s5XDjdIHZ1lBx0rUJ0pt
yx8mnwhbix2JjacfkWS9Y0NrgOmpJ6/XF7KhdtXk9ioAy+DVirO2YU589cHpYrIY+YYbS57nCVcH
vtJfI77427akbgfOckWB1n+4DjHaW2z7M+J5T2xsnO/puwbC5AGZLxdRqkqCgXcx4ajDjc9u+GXs
lXlJtsHQRU0BNPJeoThLwJxoKdfz4WLELPuULXsT1MohFhq/NbFFXtQpRRf+OtZ16j5wWFWuzg5W
FtQvEcViooXLADoDYnwn8svrLmA4VVye6BZkb5GLVbkAFXKl9GCJ9e+2mOo+dQlYUtJH+BVGbeos
2cec1ec5CxmlUek+5u8NdWL4qxLqIy4LMIwXUWulDCDxoIeCDJqUJzPtiz+PG8oNbbr8zmVlCPEc
+51LeAhqoiUOeZ6jDH6VIaua/ynvQ9Qq5/ca7vyEMpAD6dADYksu+lRS1AdPAlmbnHlQ4iyOVOLQ
t9bY/21vp5WmCzlh9+h3HJiXznyRuKyhrq+/ln4/Hey6T3kYCAdCfXHl1Yt5pxO1JpvyxVB0IzpG
L87qudsnKrS1hRQ4TEmu72UatCt7RYhCiUHiRbaj6Dkh1fA/ITYfP8i5cNqjQwYD1X1gK8+mbVyr
E03GOoFJLZfWR7LsXQ1CggDvmNzqfsVzjVTVdZrBa0nXcbxk5ojsOAlg/r4/5vpkPLRmGBjqxbJA
iZCj1cG5j33EtSI82hl1atZFadIHNodcusYy5ngCU1o2GJEYG7mTK6Rylk2e150w1IHy/edQNy8N
eyvBZAKz/ZBfe8+pSV88bOAPAkSk4NijpeAveDBOxvtDozctwniWHD6mftonqKc2oTJOd15hTvlA
cVEUuqBTacZRXlmYoMdN7hrYMAswoBEd9nRcHQ2lAM4ohRwHUdxLnyTpECK1qyOWgjQPvYCFTpjG
Olou77dtLHvo4n/2gDF5R/3L17LSoa/Rkr5FBmf2Aw8sXGNdNPsn6hfNxzYvc3pVPfsK9pTxYCYZ
AJvSwWk1xG/jV3eDKmmmCHKgrM+9wwVRqCMgrYuQ+2ICthooFBcnNa9PJxY3hWNjnkP6j2+tva09
uAqPazyaAekXRH+N5zqzq6guHgTgTO7DV+loShUGt3W4k9aIRyiMWhJO7ENfL+jgkcoDqbLxCG1b
CeTl+sLsiF8hGNbU9REPW9o4jnnqtw2l23YTNMXtH6mbIk+DqzipI3ZDUZX4JeWwdbIbW3oLqk7Z
4lR3q9G2Pfs6BSRpeSG1lj+pQCzBpd6fn+49pmc17IxOwur2Mfk8rCNlPdxSdDKutml+xnnTWwyW
M5lODHH6ZyGIcZIokp7LlCfDGJtVXZIJgPCwtMRE1dTMequXfnVT5o7NoNBbXoM/9eYLi7OLZht9
Abddq5v7WAUD1sthP3Q44hQjwYsOyH81F9p+TykHJ8XmwmNAvEj+/TCLrt9/0YKZoURds4EUVva3
fu7MIsvzFuobwI/7dfdr4n0zTCD5UymS19G8TYyZP0R6OQXCiyxcfwK+XdUcGA+Jn5eJ1OSzCAKj
xI16bZ9Q/hW4YTRRxqNwbHz0ingizl6aW8yBrlMBiROfVitwz9ih2pfh21qVpJyewP1dtzJnC9kN
Lm6I8aFHPhYWDzbrS2uOIs6Yk7P3mSKbYJj78Sj6SFNn+dJ6ui1vuzt6HeyjqpNvPS0pIDPkWShI
RQDl0TC5FNv3csCtHXx3DnI3hoN2JbvPDPW32OixcpVDrUk+y7YZPx56j7UA14b0u5SyJ33lV3wt
VXw71A9MVa3MfTUX7EN1fWp+nEgtRSLtkKl7YO8Y30t2cjIuFLjniHyqf0/vyqWNhO9p+lISfEsc
rfWANMu8RuMan8LHyvK7UV3PBiQzNO+9rDe+r0ulOLr5QA/77z+Cw33HBMCicAQ2DCYZLTCu6Z+Z
R7cajNpGBSRLA9x0j9k4ZfY9VWmTh5EuN+fPCfdEbvII35cWISxkRHDjQBVf0hs81LKC6OWZLjll
neS8EeEpBHcGEwm9MhPw3+gF2yp4T+18ddrR3kWkmGzNUoY6ESB9vNJFcqjvOiFhCYz5CbCb4YsF
nRdJfwWDd9pD6UsHMShaMV+7E07+Q+Gd0p4rJlRvqCvjxILN3znDaUJFp1Fj9Mj1fyVFZ9JiIZn1
9QAd1drfs/cseP4nBzv4Efbri/3FzSlOlPREtjLagh8lVxn27JGkZQS4vh2eVjR9QnXj4Vm0IlH3
wTNCUaXyGKXOGHDKyd+FtbcslHexf+2tsIQgXSCW2u6bVLfAfwauFlCTaXjEcG5taqKHR36+ksxV
KIxxPg79UC80ZDK5m+kMtZJLDp0N6hdjcjGhWeqrMFdLbFlKdPKLSr48N4QMI6rrb7uQVVSdl5HO
2fkVIlmF2LzMKG0YB+p/hIeyTlEwMJLKI5yJZ85KoHmvwEJeddKJhAbRuv+uZQ9paSu8ulVyPnrk
tl2WKsQi/HNMf+WiTSyxlsHlQgZGCP8kreBBFOc7Vo6jogDrjN6jMFV11/ir1i3ieEG7sKU6pfFZ
FD7No8uvmH0cHdScubEj13qselXJFx2ij321uEJtj9AGio+c3ALyiwktXzqgyInb7vMD+cxazRBk
6u5KorYdEu7gmq5sj4pqCUw9CB4iBqJZAlHhqtEkHB6gFVpyn60bx6sl9fY0IsE7YeDXdEmgQelX
MTuPczmpoAZG2pkQNtuo40w3KhkaiSb4TxnhFjJPpAbg7mSvVyVKlzYsISgYy6iO9Zs9P2Otvql4
9xDNRrJgKzM3C36t/Uda93psRi0t5bpYDOvlM5pFugM1dLeVYyJBMYg9c9D8xA5H7wnbbc2JbcoW
KM26lKgbeEJw5RxlplBOG6WplHeU0F8xaIKrlCScgBPjsoo6yb50wT8VMKUYIZMYx7pXkBgaD2v1
4zXPjwd0+EtJE+uBDsyF69B77tzd3c4C5xtzOvY9gfaUvZH4RPtziNSOuq0RsRWO5mE+/oWXfJxZ
RxrdQS5h3aP1bb8OSr1ZWMa0J3sdT8I/iF83l8H3dQvMup349xHmSaFR7agbG2qabMYQI9l4KTKT
tjWdFpQZvgrxFJBpPOQOLFxqgi4dCw8Eq/Bty0RYWQQvGFiKtmiANrD+MFTX9maV78TF5VCRzcTP
jlhNXNGl1lNKupC3UaOdX9Q6DTAnBp6MJO5zaJo3dwO61aHGyOE5SNXc/KRQKLFThfn9yYspvfeN
o2YKB78FKSmWaEsQCWoJoOR7dxufXxUoClbfThmPDcBMJLm5G5w3Yb1Rd+KZy5/QpuJYUniXeTON
Sjsmx+n/8zc1ItNOp0myweBI8PHzlfJfpWw4FhRhhE8FRz1+7TytCvmL/BY/v88IGOLx8ZYAF/iu
egI4+wTLsroZisHQ+4HKA2gePuDGzyUHz56NSyHlPo07iXUTVcNJbaZsAUC5gfBFuJ31ceoPdPgv
reSTqXFyP8/J2qUKL/thfLafmRO5SEnAlKSiNe/4FLnDLnxpULYAR2Rt2hPFzwh3FUUdq97bPLsl
zlhlekMZtJk5FzyEuVwdGQ82vb3JSllc6E5lLRM8FANNIpyX/kx5b6ImDbweOYMJKAtXjhTTHIR1
qWVVPWT0rSlhQl+retNzEtrvDisFlNsUyQsWKZoffEmO/coo2ggTV2d9lDNZiGii5uO8sq7XHv3K
MbJ+b5zDw6iQZR3AaXs7dvfdDvYDMikiWM6C2fjGeJIl3w9bJcP0kdiZ+HEpSK2phltRlJbYRwSM
fwxGXOpZvWKjZiBUCbGhAE0IYF6CXSHiqmpoyasmpgrHdxmrtItuZKfZhlTNsjuCLJNUPHjX98CC
XE5z/ZabzR4heksAcAkwijKkvNiK3IeYO0k/iPuYJpZJX4aP4KOqfk4BBSYvDBGycCTHd/h7q6LY
yGj288+OvOW5gCZd/1VNHC77vA48G9XiMj0W88S1n3H9WPvE6ZcFlI0ETuWoEdRq8wMWW/8dehxz
wqlbmH8bLEupKCIozoWJbyGmW5Q/7azSFUhXNQDBasJBoqu1P2/gAA69E2hFB6BMMK97rk3sn2ZC
uOhaRGHU1KsqNSCCSrInRNTHYiSfPLwievwma7peWhzr5PCxhrw+6V7vDzMsY5QtAGmz3QKzZhnK
3DpI1iAtJXGnXFiU6Gn1RsOcsVi0dd/FJoatfRM4nETZZsmDc9W73HGCPu0XdhE5qFymA3mWz7gJ
GckGsMILhHImfPn5LxjOwkylVe7+IRect5fdp8mzfxiGsV4qOSrTawBtgIa/qGzVxDjWYSNDNFfw
HFFpFhtqhw37FJOrKASET43uqPvMAGLOoYyy6FYuP1GDVwlHOMLns8YAA4MNoCf3asvxSkPqp4eh
VnBcpCb0G0Yh8Ma9UnmL0qEuY1ASjXsYykbSQRnxw1hpgADZd9C+pdP9tVyMCLjc1GEPsLco5U3S
GivPxx+AisQ1pcrTI6jGUwTWJ7jdleJktU5MnFqKj8eMvMoJ4fR5dy4RI1zQoSdD/QFA69ug+Smf
lK2swTuclyJaRgHL6cyh+6/mZTWzGc+6xQJXEHRj4x35U9+2Piq+d8KQ5FvxNXL3kNTIRoDI38wK
GMgRoenXLlVCv++hfZXyn6OVvNIyMNHKz0y+phaRGMWmj0lu6WZau+OwtSKTsKouNa+C/Qx1kKVk
FQ8ECl9G7rVmOZXlqsJaFlDTp9rZ0fMijBUxt6q+StaElEal+dM8RTZJQXpsyzrxW0eIq/Q2de4e
TG9jbzg7nevwaB2Wi63K8cF+Zpx+FcSxA6xZT5e3gHBhu/QjMPs+XQprsX2Mks3U/rXZNnzjiLOi
Kh3dUu4UnHp7ShFG3pDDSQAzxx9rC9DTs+HQIxvDHwdxXK8eG3jo9EUR2D3vLn2GLAJuLcMnbXEl
4PJgf4qie+dpUUFYaOVOuLfOT27Rxz7h523MZPwb4wYBAEsZ4P/hA9bmRsXRUXm9Qs3HOUfgvlqd
i+Q/b4qA9AAXDSgh6f1oeUNdnw0SEjpnWd73O6HKlv6SxFDgskXyWxw/Tr0/idLa2dYJQ0p+KXEz
OVnMYt0o59A/HaUxmrDp9UAsQZGaQf/0OKaOubtSi5Njsv5rWpjBcfVU8l2CnbeF3SwjAXUMJ+IP
cz2NxJK6ty+EqScr02vGZKQfhzPNKQZb0TkJbOM3WCg+Z99rqkhx7QizVLySYFv6YobrBUCjpzLr
mplE028OumBe8wsCSW9+uHg5BWQZn3sFnSGXSQmwDv+wI7N4omFHEWC84wuJf/tcdloLUUIpAQhg
h8qqAetEcUKwo9JvHX7gxQdLftLetM409oYVEt4u8FfBhzQNUxksI3KIiWafBX3KTub4FY2UWDgW
dVR345yj7JrEgqZnk/jl1OFtunx2O49EZMOHrS1eU9ApLKLLIiinxRIC2k6qZ0JOOCNonU6Fs+pW
52fJC7G3Ww2gAY3yl5eq4RmCFfdPxjhtU5ohrwEprbyAfTfn0YW0y1/lpBOXSqd/sGxOy7ozUEIk
uhJCvmjBIUU5SKFDH1/h9KAl3HBCWSG3mA5VofjiwYaV66VuGHMqDs7HbbhzUs6ph2/CZRpEv+hP
63ISIvufjUoHQWKGPss5ePOTA7zYPNG23ERZgZqVkzUCD8wcDkuH4A6tuqEZsMH8XU02AAxLJv75
d0ecnipqpSSeE4TjVzUrAqvmL9OxSNJR9ZhJuvFVXfhee5I5L5ThK6Vlg+UzEkABcd3npr6zduuk
X0MvXG1MYzBfPFfeXz2U3BGgMP2r8ebcT62J17dtgEIRZf4f7jO/T1sAoWJx+B5O/ScFGOpJyhUn
P0A3N6irDQE6bkGC4+ywfUHacvOAqnM81jv/EoUKYs/D6F0uW7DZl9Yb/WUoswLbKSmnB7SaMhiz
/LGn63r8b3cVXMnUwby+6hqmbhLy4R4u61Zvy8uGamUGAKjw+y27j4LFqMeYuboIxkKWRYlwsm1P
v0LpTvarKCDmXh+rkW3KfwdhS2eJyb+UfTt/BMIPz8AuZjS0nOjYDtDMFGXh1WwhVzMsIqKKl788
oi0N4wlg3XWsEaoRMrzzcUEslTeJfhdLUCse3BygQewk8k86YB7lB2UCm9/oaaphm4rNeUu1LKjX
pOTS1/x5vIRnW4oJN9Ma1knGuPrTExzPjrZRExj3BuoB4cO0KGjvaPb3VZGgagTb5lfd2h6mrtUp
FcLDnl3+JnE/XvE15v820vugnUF+if90msKqPtwpHCMWJ3KlzhPkFjYdTSSrZWw6B1FI14IszrYI
Vx+MdQHTeg8jS4SNumjInD5lRtBqCtekYCHU/XJhUOo/yFnTnCsuuOEVQ6Jjh1koVg6aSKJp75P5
rpcp93wGsK9vG0CYGfzobhOj1BCFmp6H6Ga96pw54ip199New2jePrCfkROcj6OTR6d9wqJ/Ihgh
eNdTaq90oqheVHbOIZU06ZtIzdGPjtexUfsgW5/WqhxadqrhF4QRzObp5g/8H+n6OiIyZNQs7yeF
h51pa4ih4TP88RvELt+nSJ6pItEuxkt4Qitzfgm1kZWq4t6qEtGWpaOdCd4Z+uzsSW1cgj17g/+7
xMH519JEfdpE+V1anIi1pGcVbzaGJf3KGd2MhviK82EAt8cX+9t9XPlRfX8QcYB51fTWSJwqnK0X
k5Fq9NsTZsZYKcbbwZ7Z6r54s1+v6YJpDJ7yyYjiQdo/VXZpnoqScBKQrJ46LGgjk4IwYP2oMBNO
P+PbEItDQo31A7qVl1myF7BUAGKrsyWoj9+xXfgIyYhbCgc4r9yG3MPevtwDwo++gpY4QLRRirq6
KStATxAAYp5/cZNfZo+CjolpwKnM1r1x0K9frKB0gFjOG7xcclm9etAChdUJMobGuf3GqU5YgQu9
NPJpPOF0JjaLUNingXxxzxwy8Wgf4Uj5Zz2pQV7aH30lvEEfnATD5wB++YgFJnUnq7oNBXn5jfjH
j2Cl/2FXdAmgrVmqxlnpB0WDfds+CzzhF26nSYIBeyW/XsC0SFtKFgv5FjmNh0CymYQf1pb7ciXZ
ATc3Q6erPvmtFSx7hquf1JMgbAkOgrGaYGmPFnOpItVxX6i9caX1bKZky6t/EhuUWCMxrsg5lykl
gRzGKK9rDFoW/fxCfCBeGwwGWqoFsHCMfw9VgZ9Ze6icSY44jptGw5jspueH3yf5qQohOitU31Qb
hB4xCooCiGDhYnKajH37Yk5D8T0cX4jDZBDC8dxjB7FWAQeYoATIKLv1c3/Tpxp1pA7T1Rye8NQ5
hWj9t3o8BRYnKUDbnGtQkjoTallwivrjq2mdLWkw6WnU3ZlnpTiXUQmAbWz2y3huPiuzJyH4Ovul
K5x/kL+S+HmCqvFKBcQp6+05UJuMKJcljbaPw9anAfoWjuG5WiXTeyKoKvHaRENewiuj6jTauNb2
dvB8sCYXGqISkgd6rblG25kA6k35vKQFWELXYUkVDnipwsUo7emrTgxo5C60rQ1iOrccp40Ft3fJ
lfZKBxocr9Z8QTw+peQvKkTYwHKCreKZQEHWS7plKKmuuvF6oi8gLR6lYNh/NQclXFRI4/0J30fE
watJl17I0zoSoOkvcX59Df0wrb/Gr2J4BzklN6gZUhOZ8dSUQrSSelLtIY6rwvhccN06RzElVd5r
TJc5HuMJSJnRF4raD5nwv7mqJcizaUZ9QarFX9fgTom+NCgPqTa8zLVxk7Qx+Pl3B5zBQAlfpdgA
vRMJkTVHAWztShAjTTgzNjB7nI/QkTv9wJL0q+Azu44Apkpwg/TgVIHLcYe/Z8GGi7mnhLjJPWRg
JECrWFIzB2qVt8d+kQZvAOzQqu+QoTCEIkoGODL0/xwbFTfKJb/Sb5tsnOV0TK9rPklWiDUzqwO/
ugA1IHaHvf2wMfhx0qykb2mLF8MQ2Uqrn2Bu7FWyZ/hVpDX7Eu6zC3pPp7pqS7n8tt4I88Ky8W3z
hAbVQQurrXu07HX2fbUfFy/whFKNrnohcICEDiD+DhnArGc5j7F4pf584neqBakPqxK+tEp5drDU
8IQFT6oASWB5EhmuS3vad0IjCRFE6HXyp2HvMBn45Qm75GMaSG9G6r6ctFDebe5+OdYIHLx2nKhn
FxDpbr5jyinJXklW/Fd33QG26oVqNElCA2oOKueL/KoGbUdFCU0qCLOObZrWLuscS2jOVZAyhojr
q2GAGjSbzyWFgnAVT5vg82gPhox9DGWRrQ1OgCxZrw0wILqpr7FgfClScPjex74bkn3dq64nwsdO
A/bcxzmH9Y8Rglj8651Hq686iWb94eX52GCfe6/NsLvacG3zRSccRzMF9gSYatiD+4mYJMQ6lnAe
39PHzqy5iXBgbv3dvR0veCMVA7p3B1YxkZdCLORKTtVYCPgD+hyVt+a/0dFA2vSTH5T4HKzREo1Q
f+HSATuS4Jj138S5sH5Qd+ON3DL0H0YqSiyd61Hba0wVwlfmvtCZp9MDY2Ey3vQ+rwrB9Fpj8LTZ
8amqqEdU3cbxNXkkNQobVreJpt+yZfZaSR3L0IDofUbYmPACQ1AGUII/Pifbys89Ps3z+agNACi+
ABzu0MLe47Rk7Wmba8sZrsjvhn+g5GX+pM2oW2WkLK+uacD7vQjkKHy7wSkAxo1CTykGGuLDJZoB
xC8TeoLLgF4du0Ax2hYA6RFN4ev3gOwqZICeOJFXEVfpx/0bGrhF82vdBXG6dcdaT3yZ5pGsWUBk
5Dkaz9asPq7ELu27k3ik9BpRj+k/7NvRKT05qZMcRioadNoXgF+YmQ5X6I6OB6zdxykA2/vOz+ll
puLfE0urBctk9HPf9dIM4nGOo7aTV7q1Gfl7oTNa3O2M44SDF54cS2jMa3SykPi9+oOTeo2sFaeL
U38t185hxwcj4uahh59iNbkta/d+sfOtwH71XnBY8KsarW/4JzqLpXwWpFRhYqXQP4/XE7f4qMl9
M0yTvIL6pdKp4pMj/oDQznNeyd5GdBpRy12Po1H/UCC14SBkWSQM99vPBhdZEqe2Q2hrCoHgrabd
g0SVq+2qHaEX8pDdJzlooZVQK0wWBqYEJHS4SbxFhuxcvUuawR/E0BsL+rApOFeGiOH6b8iyk8Ut
cPkDXX9kcD80IjdlYtMtYzy+0Q0ufatDlefF0UgQrNT9VFOWxGpTSHbdXBHnVvTHATaw+M2Kdxq9
N+bEmmp9mzWOJ9MnDA7jCnFDtEou8ytlR6hMK3nDxc677/3T+N2OSy+G47RYDI/wSAJ9sIjRcQbQ
DEwpptLt232ztVVRsZcDzw6aRFREkqXFwTg9Tjyai9obRyk0raAO1SMnren+fUplCqPJKsuxS8IJ
f2ktGV5gO25N2urnVbZV+kfJVAe0FehH8e/39RR4OYbLSbDzmJ6BdUzB3iYpegG8ay2TJhKAtrjh
uanOwucQF56rbt0v+ktG+kfJ4Oc4A1JM7IXKUmxUFqvAjT0g3+tbqzf14GmNHkX1NWQxz8rWJNuU
bAjwmdfHvCfumUAWLlyGpmRYVf2qmnfH27hNz7Y3bTgYhwvSUw5DEWMZM+SvcOmc2utAFN2svLM7
NllLkeN8mkMds+wDKMHE7wEoLg/HPciScvzBjvZsl4AoQOB5NRqLN9IRIQ29zAutxgNOf+kQsxga
lsfilfLjlWmFET3O/8gP6aIsN2UXeIpx/9+u5mesMubV/JJrntvhEiJiUolHG8dDw5I7XK//2wWB
vB1Kr4HTOkZebaPO61sLcBWKQqmnNUMX9yQO3BjXMVOChjXWr5c9pRzqh6H6jZbBfiCEQGyzxTDr
a5VV1AKJF7ZctMJodnMRr1p27/sDmFLTJhYnxyDFEqAN2uhn1YYyXzJHaSCvn3gArODngOyP5a0y
raJ9/Ar6emCw1BOPdQQKFsE8AUR1ssrActDQ19mfnp4exeuz35UUZnBJNnK2+uQM4ursW+mde0xG
HzV6DwqRWy75lwTXfYTIKtg+OMQwt40QgQ3NvD0RIu6bOOe6tPL9nhbHJNB2OuUQnw9ueDYIUDIg
64CWpcmum107SQ766E+WizS9v5s81EDedr9/FJoN+M3jc2MnMGuLwNBrziC/CzDP1gxKUMG+e2h/
AOLJMpkyWjhikvEZOjtcOe4YWkAh0IDyWPpYaTt0L3GBuAYMaNFrBXGHN/uaj9R3xX8FTjTSqHhR
67G5+yXMBHMFKVusl0xeRNY+4p/bqUbELC1fygtkDJ6PFZmTE97BjFNSmVTXs916T2N5+16oqCc5
HVsiw/8o1Ayu3QWfSOdft/4cahZvZU8Vh1MkZTiJpVVq0iBwwQahV6AnIqjefRLDK9X9/9DtO6rr
58yRW9z7apTEdjVQZz9BZdVG8Ev7fL27iVJV5UbrTQwH75ZlY+kN2j56Bdz8shODnc/mPCKISB7U
Zje+ym5GI08vkp6r1ZX9e4iYOfXK9tDHN0Ti72w7Pp2QQ+H343I4Ou07uyh1MZuCOUnvMHxKBeif
V5Co1AKSfMSVXOzaM0gdoNlQ2iWtZNAPfJn9z7s+RWXWGgYZpLlbLZkV11wrrR0JUBbLuT2xYiNI
AlliDydb6EIJrm06avSG0WdpY1zlwxro+QVqUG4gR6WBzFTDBWa39ugP3DjbtRoKp30EvtdDFvmR
/F5A3VOW/9KIEMSUVHDalpHiOc/d+F2jbz4QMU5fpvN6cWKwcUWElioO7eW+wajYEHGCeorRiBvb
0F8+3CongUcTbMfe5Nt1NG69q3dUiRPKyeAMiWDgBz/zTSiCNSSrncNicj1c1FeyaHczivzblQ4h
a6IQ4DOwWIzAfobU6GGq+2Ko1z3VdrbyjJPHPCQVpmmQ1tqAh+hfuTyDYHDHRZVHzCk6VjmjjhCJ
UaVdwfBTZsLs3b6zZDHJVzCV9K4O9moZUz0HWKp+U3SvXZ5qGoTf+9LVE2tKE3qSBgrmGEAYSImp
CZNtyXzRAJtt8EgBrV3XIekGuoKpw1iIcMdI/hsrJ4nam2pzfc8yFbMSNIn76XqYv+QyW+Q5Vjp6
mZqKAXEZjOiNe1LYSfZUtEMlYyFgPA7ZqtlBAvCYUZdomp79JI/vSOZN60/WVbfK1KpGrkRd5pc/
tqYTgJ1E7YMnQqb4Aea9Bc2BBvNUq8UA64rP/tQsOiloRaTUOGtlOpsYsLXZjQaeiWL+ytcMDdE+
qUhmEGdKlHWq4e2PMn9La/9LpagwZZhaanHYcNGVd5uiNBn3epABygUOkebuoaw7nSPQ8CvZKKK7
QDaNyU6FHKPhOQHJcvKB3xiq87GwJqVp6284RV9DQUV/GIF+MdTdY6n07KqVDAPKc7BHPE85fYrh
Cpf93y7hXuhHumFgK/RpNuymsujH46iudCpfw0Cm7xn77Gup1eOtopBBCsd/30smjEd4stKp6nau
ohYyKNVAyfw38QuE/+ODTCZy4lj2XyMaYoJqRXPy1ncdu8g7UOpWFurN/riz9p5ql9TQH+DNlGQD
/ahKCaXZpRl5mlUZDHxnR9tAIQTjDeFdWvLBZH5iooenxN1IBGM0pBr7/MHapUYAojfq946lsfsQ
1qSnFcnoTjag6CjbkxWetUx+TxQbkcpcRsq8k6GcUDdpdGUfd91i8AB+Ax9SgWfXCBfvsaWyR132
TSM5HUZdCfC7V+TXKrHhDphcwNGlsdgsnglMW1uHtrfxJPAcMXiUdRa5zDieLJjKpVaV/TY9v37p
ia3XzVVEWz1E8bjjPDxRMFyH2r0KOWyyDy2XF+FCR/44Jq+JAQJc+as+VnETJJrDJ17dixLrEvOQ
elTXH/yuOsmSTh5tjOyV4iD1a1sNXbMcN2+IlUktGv1ia/qK2Tq5MtK/WrUKJxV57UXiCqs9RXH2
5pMkQWLmw8/2WugulhS+N/pJeKyyrgvmvmCDpdZbttpK9JYUqqK8Tl9V14tp5cRhFRbqnxnHJ1k7
mV6Ie/rQ4p6JxWTjVfUGEgBSFpMAqjhJTRL3d/o9PUKKlf6awhVi32kP3uPlhIkOMA8JDroT1leZ
ta7VZBlNoE5dkhC75Kk1q1QdAmZ/GXxy2IBgMJfFij1wSxlqxUG+UECqAebLe8QoGXzYsXJ0ZiEl
KX98S+zJXd9Bnd8JmsoxPaKpODhpFPRIOI8Abc9zRG90ZmgEzrgMAbl70bXioZ3mzVuFVAq9/TiH
ZBD8xyWyxLAS5DhGnQ1lc1OIRAgRwuGXKFBEsQv5EhTbw4t0ImRvWnzHeJeamhBvhgWJCGbW/FxN
vdl5Fo5I5XoLYTiyVPvEKN8LpRVo+b4PT8GR4JOJ4wRPW3DUI122s7xshOHGpbpBpkXljDWFNHJs
95pyUxaDljIfSX5Cdw+HYTWxH7E9+iwdzVth49t4e5vHtIRZaKjIRAhqY8mKj3WjDc2X3EBD50cr
uFzk+ZdhqYO74WNU+zlFR74xGA1PvIHu+Oolr1ICfMu8mhn5FYyXlmUn7dda9OHJnne/kJJC8Gtc
yYcHkVtYMewDQCVTIEto8rcYxWA3urrLGxlmhNYDjNi2B/CYPJru16/zVfN5HUPA6iN7xbt2zOes
NbviPC8hNlwlzwewK2eyD8aBfwoP6Uric2nMtvwDTSyBW4MNpvIb6qrOHST6M8hh5D2464gKo1i+
nHAumbP1ypYtQ2llKdSCyHs7QCeSt+Qw4vwEFeQsoe3mxGyi6v3sir7tMC2L9cTV5f9SKYNDEun4
Yk6qV9hzxprf0kTFXEStnSn0l5/LXKtu6yimpgo0wF3J4XeZI6Eay2bQLGOnEKu5z1kSPv58iBQL
m6G+LH863SF1P0WBgvbf+KomUvlgfJXQRXQQ3IqKqzh57eBL9OPoReSo8MUBonyWSKfjUXjIl47+
d/V7XgGL+UGlAJN4lwKiAEoQbJt4n8UvZp6tovALUWBYj0E1Fmk39M9Nvqeftckx2tNimYfnPrdx
hT8PuRtTMNaoqbfx9E5GR/R5IWNUU0oFeNRQW+Q8Iet8Ur1npJTT5HfJnf109QZAQrf56d+iE0Ta
pBxH8AZ+IfQiMl15DBjXrgJh8eq0nl3ldC5SX64RzXHI6X+5tgVY1TZZobDTzb0eR1BooEphCkhc
9f6y1t5SmK4n+8huBf/6XR8EPvXF8fVQOIfm67FlnEjhCZlkKq0WTvFSfdiaXny2i9+LnqQp/U9O
sGAjmN+Qdtxzkg7XpNWYLD9rvgntbBue4r/Ci/Utq6jlYd0fAjZuZL7qRUzJjep7LzTBI4iDQXmm
pHusc0GgwXjRUbT0Zc9Z9UWw7/pBknQ/OUhZsfgrD8ahvwT0d2O1Y7/Z0qc6M+gVfhCdgYTbccoI
5CsVOMkrwSHlcuWt2grn+NooikGlXfpPQJxRYvVltbx4Zgr7972EUmo9mTUIQ2TM2IJ3ixbIvXOF
9lOq0QdsiuhkgcFeS5VfQxduRC0zzXNA9cfTQXDpRDhGOH60tpI58Zcs9gpz6dfGBtIPa43zLaqQ
nAAEJT8T0xGz0TrCtJlYWLEmBmhDW+C/jvwWcVl+H/fLHo50EUn6lO8XHoVEbEU2mSo4LchYtiky
zGlNcM+N0Ld9fjpGNewdR+txZtydOCQ7cVW44TDMr3T+4xjSboocdqo2bq8g5p0ghkQX4gDakFns
0zHvIjxkVS2MCp+czMfWQvuhZej9FUw8zncNVow6fCbpYmETrCvc+KDkuVFEOC0TGhL5Sk5JHrhX
EqEvbJ9y3rCH0S0GKjWLZFvM2HFr+tTiSwmjyH4Bf/xfM1vkKIUSejvjE05gntm5TuehQebYFL8N
mo1LLh64WXRPyt9CejWU8jkB4xx6Wq/hiP4GwoCAPk61ulTH8JSVY7ZFTGHey/hwCY/gwjIJKHnu
ZYRdIVoOJD32XYa45QzXrFAGWNZ+AlhPMm2TikbBayBRJxtpcWrhqeY7VHLlzCN5GgUgnb45VcH+
4Euz94Q1oV1b8YtMb+Kqj5uwmGOkkQXzJfTzrcok0tXYU6Ct2bHaI7q+d2hKuPjCcs4LibUYwgxw
E8W6cPW7DbMvZ7nXBNdSSs2bNTQjJa8PYgt2xhnL7FWgQWdvDFeYMwfAobvbvDdRc75OinQrq0bt
CYZ+V484gv886vUkozTpp7Emh857O8sOtfTD2Pf78TW1H3G2W1ED3Ls2hXWuT7XOsbB4l9/ekGzT
LXObAxDZHr3I+Iq5w5FnPhq7uN8nSeieVTPZ1zsajz1B3lu1QC6AGA3JS59LJv+VqP0rJZmFQQXX
8CWhCxzdAB/2kq+2h5Mq5wNgqlAJpeeFs6/dgIq1dObx7Mbqrjx1BH2AHxDbe70lcPH0CLRXIEgl
ny05WYSRwTXU2Ec7vg/SjFDDcZzzKlNz1+O6nQgRukCZHuSWPnjKYraGwPaHvJwprQj4iyS0OtpK
KNkKMoGyfKICIyLvPQiOja+dUNKJX10FQh4l+Rv9glBC3prme5zGcIvw8qqwO2trSFJMpQ4Bp/pj
CnS82P0NpN4LzLGrmYWRGkHzZ/TeHpYAtmfLmSwwRhYsbHZCQ0xBX7332Fd5DwccI2p+UFsSlvAv
4bF0loYIstuk1vzD/mLrGCZdKFNRrbxjfK29/9RpZlIR6ux27dbEn2j/7WSJLcAis5vONJ3Zf3qK
b0BP/4VelJvKlt5iy8FKVc0MxA0cvRQ3oaY5958d2NgQt2ZNVSCofT4JRo2SDWKH6l7iyYgGCazu
6lfqIMDdIzjlz9XMTVeQO6vW7piReVr1VniDIVuWNFkcSsB0fCT2YaVBDiSwyA2EmE7slitb+51i
+gmTR5JhDvXcqw6FMW+bnA2uKrcUnbtDsPwY/dvJ1p4Y2Qkk+9bpeawmC1/y74xfDzu1XZ+Vfb/B
F8jq4rgqFITjAlclGf7wnEjeY9lbOCF1tTbvLXGU5s/ZQEyjdc+IIEVb1JDsD4OIp8FimWRw8Wti
n+fX18KxRNBMOlL0OS1TajBpq7/++aPFHMOBGTfsU1SjSdbCOY3C0uRIJqtMPopylfdRdjLSZ28a
U9qFfOWfVvQFUzCO1RvMwfGTRICQC0o5A4gbJSnUHftqodktjkiXntAC1XCmVBf3MvnfYb4dphZ3
n0F88agxHBCcJPK/wVKNcDv+O/CwjiQpFUrk7uza1l743zH+O4VV6YXiSQs/zDefUQRBQbdEqiLa
eaUjfQ5xU9EzZ1OhokJ/iTSmOtb7mxdIfxKPi/G8l3r7/v+X0F72xhJAZZnPgaaP1XheUOruqpMk
x+e0b7yCqnj3TConC2dNJR873x9W6vbsAunJ293dKoCgO7DSDpS8huA/eVSA1bNQh00rLB84wxcv
kb8nhDcxvpb/tziOmPj9uNkueAWydUwB6D1lQmN4g7AWpd3OYkwc6JwW7f2WlQARGzBPFzDyCUe0
nEdYUiB+9FjzdhCoXobhSj1/O20185NX+3qSIX3f+4lyMi2y8DKVV4HpRSzzMlDDCrWqSALr3Zoh
hulJm+QfGZ0nw+ppDG2nMXJSJZIZQyEnJrN8hIPPrZvWKuyxbwc2Wd31dJqkrE/3ek8TVG5C0NcW
XKtV3VU8c3qgfm/EMe2kHqOmJ85ujo0CVk62HMZIViSE4R8ezzCsTggF+i+/gIxPsa7TMln9JmLV
3yyH6rLDppTNuQLx6oU9melY9rd6WPqxigSznsKm+j6YMSp5hJTEsw2zFsAH3oofPq1pZos2KtjZ
TKn2Y2Z3xSRtn8ibcZo7uFWfZphOTTg9QyrSK2KCXJWgoDLWJeueuKNQhh/6majhLXbsYDek4EcG
F7eJUnucgdT0+3Fr0vjyQihYaGQ1hqX7MCwkiIEliakiF4Wu3crLf5UjvSBP6zESytvqjsgVWuUd
Y0Nq37PIkLbdKnxd/2ZJtDqDHriJBmUiWgdk/eROTiNCIssrs4E1xa2WA1d8hnF3+LSvXdSWOXIC
KRWfD4uh1q3xc5/y5ytkWajsPrAWy8wRmk7QFR3wf9yATH1KKl4KFiox0X/GUcBvag6J0SRSQxUh
iVgVEozGbrFyiPKnCNwElMU+WgMHcfMN2bfAfxEUouedkjWLPzoL6vzc9TlDLRyjnQF1TFAJRGMx
0mxHz1+LFcvjb0hGQoXHbFSk/hLWe34ZB9c1Y4MdP/PvUdXV/kjsVc2QXN4s88mVCj99wwjsLWyy
3FzVjvI3gOQKj5MECWnZ24/fVfnvt9vkmv4oFQe8n+jL0APknD3CtbsJJZncG8PEM2BWDLKuFfiL
HpyTnonOQ+YG47huscbKsB/Jt1HWp+pGRcOvpyVwSl5POgy2KTfPpKbPXUcoEqriuUd+RnlJWMLz
OZiG2kLxEYJZYFsWmDtipq+WZoMZEvWWkfOaR34XjlafKLuJjszNcaubt9wUtf+ecxN7LJ5MtvS/
yiDO1EQGnvkOOwXP23pVLD2/1yTv+ckw7+Qp9Gk2DbHbbQRyL6IqpiDjjgmROxVF+AXRUQWUorFU
X4mt5J4+23TqdMXRWg7CduivagoAz26CROZzoAJpPE3bAvmOwp0SFxAACTIWAI3tF90eGjXx0DM/
QBKCyclyyWF70fTzKS6TXFVDF2eEeWAHKU7PRpZ6fWtXwYSSM6bUU0fyf2EotY64uzMpTnmD7oZx
c3wBKJjKm91d80zZfCiDmdQTtjFL+5quCqWn3rzQGLrQAQxelWMquT9p+Kk9ex6r5kzVIlaDBz1N
lVYzsmTOBuGrRyCeaBBsPvZze5bZUnNLl/axV/fvfBSmcpcX5GwcVL0E0n2kVGOB7xZXbgVBVCyt
ISxFJVgaFgoAikCPMJP+Cx8Qw/Yrpcj6G9aYtIzR/oaRwFIXe5Dgx+KSskQrUYnkX+wxht8GBzxZ
6VDGB2OswaYKZDwEbCpDfKbFkBqTL57XkA1PJsPBiTyP2cF5zAcfkh7icNcPX8FQVnqcAMftRM60
36KEJRNMfkWtuQBG7h0rxLuPErCMv8gzmfx5XT7t8RLMt/jV3nnRlTitFdOXQg9LdUWACPyf5IER
JrMY2rbuVeU/fuMQLPux5bCg6491AfZNJdx7g43wWjiEXwJ/022xctBf3CHty+X2Z4Rvgag89F28
BJwnNqM+5NxRXBVN+dmwDjqjTmOtWHr2AtpWjxHI5BGW6QGrWn8LQ+ThesSudg9hD/KvivBp3i0U
+1B+YOdCKa3W+0Jl5hs7ydXcC8KUXYLIiOFzFgQERPnPLwQ33tc1Za/H1pTsZyafTVIQ+DPAVGiB
vTz1TmshB9CjjGS7ByeNXs6cdp+QqJ/LffzdhNwjieE7WtGRNAVEMcN5ttARaDHyNhnI7LT74290
+wckAiH6vqybWR1c/+c4FprKm82Ljogf4r4zt6oRSUBvX3aXOvlVaIlk4Apaq54FGOuTVMOrvruU
wTPYuHRVm9PrbnVK9McrMw5Q2bQEghdVAht3gmT3qlcwZQQ2Cmb2cjuPJsqCo0HKPM+hrqJdbEzj
VEwv0gu4dzbS7AhzzKFAyga4Gr0MGv1FUalFDqnn4WeY5ta+Qka31drmfbLQwPGnTLHuaeNprh5O
81PuDJMMJyCpRO3OC6e9sxQNR+gGrn/43nVzrj0RNmgnMkvuPbThkEUDcfXmX8PFevRCpP/jmu0M
aMYWEEu2o5oEXAhE/CRX5fce0pyIyv44fsBpEqp9D+HJTGgkbIMoDGk62N/cOxKRQ1mlLgmynBJn
m+AcHeOPrxOEtcPsmRpxFDQZD+6Q5cu+S98AnSD/yMoG0kRLaV3DjZ7ddgdxvMMsw+cwcHHY4GUT
nkNEc/nWKMlVoeAsjsuITeH7OzRu0yHPyulhC9M97Lg05KLEwJiZ0wqGcC8oCXns0zyxCN97Csz1
Xg3iwxAeCn4uStc4EhZwJUghbFpAUi5dofRMEmqzN3iNC89YIsS20Wg7VLa0mng62mfLrxgpKSrm
OcRLuD/8r4kfD4hmWujBzJjJiAshOJN+0mR1w5wpHsFoaCUgB6cmo9qabyDUvlp4cf2TE1R1431R
A+EBXJnqWHB7gJadeF4+HykAVxf8fVZTTRdtQQmix1UrZQpqbBVtEWGr+zT+4TvXFLzgtBLVqDiC
meyAI0XmA9qDxueJ1OJUImE8Fjz8B+PyWYwu+gOVgZpUJVyR/7WhRIdZWKXs19xi30KGnXQ13/aH
b3H3s6r6u/Tb24fygYZeATVlKn0gI5b7YeOa3CUUrGMCVDiir1rDg63bGhZvrZ0OhdSnCqzHgaGY
p+ukj2MEl8PxsUmDzgdCKVPxdGMklA4zeMfvOjQstQlvwtFgsd1+3McTkf8Aky1bBp3yuQ1ARm+X
MTWGezFe2C4rBBm4YRb0GCnnC2I4oK3QUsifzxIxhIoFHqUCC1uiTe92Ohg/EKhVBJE+OyufhPPw
pbeZYVU7B7+T5K5tdJnamrtBYwRskUKqeR/JAtoWAGwHQQVYT3iQZ4/c5vt3Tv+MuxlwWyECOlGc
ep58FW6+WsEY64i85HHOWwJupKAitLEp4/SDRZCd3cPQ5EvIccJpgpPb/0cbXYG0nHGRpjYVC+6Q
F1d3f+4cJs0QoEJxUTq4IH/j5CtafHtGpKQAk2xIOtrxthkpIiEEIt6xXHNcFAPvpSTwuBHKgaqJ
3BvGe0bNErA3pxK4oWWuSP41rfUoR/kBCTUZKdfwAXbFueGUNLlUUrvR8kVlwUsT2uCGJqce583H
LsA/GMW2MLnUxRV0FsqCjfA7WhglQYcpPUl0T88TrnILlQLVjv4pSQ4gX70jVu19qSxD0bAyVGoG
cJr4pBeIxaGDMx/qT72iOf9h8TzjN24zRx91eWxwu+Q0qdSpcOOTci/klphPh83uju8hZL6siqHA
LTkSYXQkRi/bx/gWLsjseKYInKjOg5DPX1APETWOJlw3spV0rXUJxGDL76VKekj7jXAlgbiivWb5
ito2hk0j+1y9eTNQv2gxn37vSS2iG3/bzPb2Jnln9tPSqGjq9LoeoQ0LD1GILLtR8wBzcMV5rgds
UlNzIKed/m3/apYhh4TiZ1BIIy5L39FmtECwMc17duqM4d6u/JNvOYYvx5hr+Bp3E6yzTOXPxTLT
oaq4LT5VVqBp+3jolNkX0PLXMVjPialDqWvsZbQUu6ZU1seSc2gXGFMcA61l2Jzgu/6SNhBrljuP
KKJCM7WZFebigUWwfUMc0SmZ7nlo5mkVu8GJFLNgGdEpfpipTKx/7/cw1eEd+blbEzmzL5YM+I2P
nAsds4u4ZNY6JYi+i86wrtOvbbLo+Hk8oWAvQL/hbst9Ot5mOc/IjYmPyr6df9Ebd580IrLilkBm
yieFrWyrrY/IfJAyrUogma7xxC7O1UcwuiYDUMS/rMCiR2zZzUVTqqxigJGFrcuU4YjWWfKGaHTY
R1DlhVRgo/6iPU+y9j9DSQrMyFEGvls8HLz8CB2Jpfw4+g04kTMSE88q85ETvwL9PWY/znPH3kBr
uSJZg6Z9H0hB4OZlVl5ruUcsi9RlefQ+u5ou2C7rDYP9a7LtgDLSm1VxMDH2kk2XrWRlCutYG7n1
bFVR/aI2JCSnol9KDOojnLordEAmmJ4z6qvvhZmy7wx47opRnKDGDLLXI6gY+/Bgex2aN+o8xXG0
nNYfJy0+M343mOZwXhv+stx94/VgJipsquT+gcIS+xclFKJMBjVgMubo6MqMNgf73Ht+BS7YGCxy
MLE0T/yL8tFVqxKGB9WkeLRTvPte7liHHJES7bfgPCstxM+bl1WNwxLiHiZWucAiQNFgJ66hxBnM
vZpUTeosZSjg4UWtSBpqvWfhtkLEMQSKmOZf7nfFG+SdTaxO1arVVRyyzFF7nPFT4svYpm+X2kZp
LZYnnXCnSb1hsIpBSMXMtBkDuelb3Dg0F0r4qpYnP5jpc2bPOyuf61igfow9xwBTDJymZd9b4+ik
9NoZU9kVnuBAUU9dxO4XHb4HaeG4nVuYev7xeHV9NFd1NRWJFoz67yOP6ludu2u4RSANRucKqYlA
L4cK1eJ08nlM33u7j0RZwApIfUUSBO0zwujFzSjDejiUaEGy/lH3Dx5u5YBg1XF8rxDexFO4Y0Wv
vQW3zzr+WM11hNUfCBlpSDyqy+Bk4H6N0Gl8cpUuXEI6/yVsMJZ773yuO87GXLIMfvIKT6oRptcR
GuL8CjLZUpy84bWCfvw7FbUxYhss3xW28BkWnEfJzIzcPp7/2xKksU/Xo/wxDAywHksz1Kddmc/s
URIVkRkMihn6ltsrTd1SYdUwq2DVyZx2kqaAClqkj/pBRgPert2rVCOBw8R7U5xbyCVHfsPTtFDl
awedXMo1Je72QKt1dPlVRrS9tZhcVf/2kk6W5EoBz9OAvj4RfV8LdSxS338rnOuCL14szG5SA9zv
PSVorkI+rWWX2mzyjB7HWpz3fFw8j7a/nv4kH/HIhyaEt7GC2xs4RTSR7Djur63c7UHsxuK8EvQp
pVsbna93afL42VUWDKn1uxOGsK0jAdtrgtSzWLwdwOhrUblkuj6I8D8Xn4WkoaNIXnaEqFTyqzet
RahJzFN0GW/g8ySA3n6lUco1cvjTBITBddvbsKXL5WFwnl7UraIt6Q7Ll07PaoUw/GSs4LJrA1Gm
LsxCdK/dtDJGaqXIV/vN2wI0ygx8Ts2QMo8wtvmYjlOV5VH99K2w/tAiiYsbNrI8qgrQLZ7hb3dg
POO2/uOfKepEkxdJ3U9OHfyTTPaoKhg1PyJ+q5SPx7XH9MmrDXLmN+hFqoSwLztnDqdqhp1OmQR7
CJw8vqDh6pSIvrGM6+YSk+PctSrSAmIL7c46lfGLelyGL7thUs6k18vPSv008fAhcg2MuVYre4yL
bkNYL32TNBnfvXEvRUeMLcBXVGM+Cg3akkqsRvK3IUvBFsnIOzxkSmsYEskjedSBEoitTEhgAtA7
v+IMkoS8Qvp04mTeMB2OBe5BB4IOCRsYep2VJvo6/0NB/dktMMS6lT3V/3AR7aQ31Eb33P9W+Rlp
ghKgHMGR+ruIIOyEXWigYG/6r0s+sE9wcrP8+VgznF62dc8s88RRyLJYFs+o29RxIKsDlwQewLyK
1mHEMYT3EzetrwVL/npzmWOgbLUilbRWpAXpSLu5Y75/DdvR3mxMXfFoUzeeEBxy8kIDv4KPi7rT
M9NBxrtf/MxKWCmHLPKNYyArzvY/9n7FzZfMEKiuC5mb+ZaSN6VOTFiwXL+Lm7PoHpU6y279DvN2
fgtpRlTTfL3hW8v6vTZLlvADWNR0cJchllLCVzar9PV7Q9F+bSmPcTVtRpPiiwwLgava2BnSevwl
Ly9SYSWzo/bUmVhUPsRXvC6XTSl82+otiMV7K+6DPqupOLqw8dp2sZ+nC685htqxOCaH9WrM/YZP
dc9c58icbsYpYbrpzhE12bPeuzGvLxvfFIv66bRLNwD0aSTznzDDHhghEO7K/n9hLk41aOuN+8eA
uncvy3Xk+8UySfoLspK6LD74EUf5YNL+Z2nxDAiMbVgi1LorCl5dOSAHK2hx1pooZemU0VD1n7l6
gzRyCGuXfVLBEhYNv5e5SvUBg+kfJqUdIxMdGmSiaCu7FpC7ZIW9KPnll+4HDY+/XCTbYpxFsgzm
WTsIp85Ex3ALVMIuXnKzZArRwZ0/dEvQrDVsJHa3crEfXdwFpvx4ouwfH0qs2rNEjg5nUMb+BkG6
1S6NDx7llCKDzWeV0Ft2EAS2YqUIU1MKwuNtl0VFobOsoUqp3RFcrDBSYWb+t28oAK5todCSB0+7
qc7swnWg92ywyyBXjc9aI+HUeCKmjGY22vdbJ/+OYUMuC8BpLFMnSZ9mciqLpKX+kC5YVErs0l35
IVTiXihpSDbT2D9OH/F5q84FRpZ6+AKcpx1ckjOPLwgPHFE2OOkKzxJGFjohWDBSuuuagjMd88/h
M6P5h4vK2BH7fZasSFXWOx5qcx0lYM1UNysLy4BxCypiXgYVtw70SH2UylIzMK+cufw4o00d4OSH
K61AW6bBry3Noe1QZjPkcRs/a5WZe/PuWY/3XUbl0vZOpIXe88O2WBv+/ah5fvhezJ+H8gskT/7b
KNSDuAXvgCKCcAE92e2GYPLujqIGDEiqpL3myJSxLffO5jMCsy/ZSVJJZSPjNIftL6QADjrR5N+p
8iE8b9V7BzLjQasZa8OEEuRCJeT4eKnPH8I+GK7E6NYlbo55/fX4CNBQcfdR5ylxbpNFK/nq1Lbo
Pwn+7fHJL8JD0HLHyYO6d12fbG44azPc1Dy/YCh1a6/A9RCUY6QMwWuUPUdonCN867k0jNUOriod
bsO2w/4HZtHk2byi4Qrn/DxYX5JxFdKhZ4RBkxkCLaDdq/O03v1OJzLiVy41h5Hleu7DyM7s1lJ8
6xBn8lUaApId0xRtbkFZ0ykPjIwhlK7BqdEjSEPXEB9/voUki7f4yA8seO7drsA9otqug2lYczEI
TvMg0UfA65xMzKdhC6wqL5b2UfaxJvNww8s1SW0lWZBZ25gGUOUhxWlhZYc9/iTPgMVnLDLCSv5c
EVGjk/YeFMp+K2Mb7w2TaLMHZxGpSN0q0dfTqz6zKH88/W+Kw51ADwiKJkfoUc5xzbnExZY2XQCC
cQPoG4frhFP86SF2EAmNKEHWwndinaCL9wJ0XlKyhGvfakqV8rszp/K+MmaVopdKvgdaWMt7Iggb
sXPqIzMcxa8hNaa0FkiBKKECtHYJ0zLZ9qUfV4vaycJnLpIczesSoqtRBkkNG3DOVmr62CtGzJ4W
YHfncsbZKodPneSZy7X+xBOsxdcU5GSlrSIueDZxeKcEEV3cxoFBNyqJ4yJIL46bJ3DVwRtuEWmj
16Z6VjsTejd9p/SlTcYjSly/LLzIi1fEVsFzBf195uPxj4DAqSUKYYMErFEQ1HSftq3q1HNywSlj
6PsNPDbjs8BytFnuhmmkf+aQQcS3y/ra0ggTCAYeyTcVfTpUWLuVsPI+D3wTYdoArNo09w2btJyV
UpA/KClF7EUNrMyMzB3TNm8R66AT8RvvIL9zrTtjaRYn/RwtYPkdvoEZB6f2SH46RxFHL9BM3Hfy
gZVkt6AKobCsAtPYyyH9MEWO6SLJtd4P/8bcDTC+lSm5SCvJXbqmrYBDbFBL6s+n4W3k+QSWSYqa
TMPK5juH1dow6hi1BobQytWlPC2zBp+VoLyOFHn8rtzCF/fedLKHOXUhjOl01Jjt+3nex3SOd9zQ
Qm4k8ie4ClrR0iFwlRhpR76s0wyiQk9llzLohYROmncsIdTNqqim+LKupT0f7oUtt0l9aDDf7Lqu
UL0sjbcw2MBZkdjcUhcPWGv9ssA6hFMUfiW4zxaHn27YdFzblFDcmrVX43yrqzw30C+XEvwbWHJ4
eZGViDHEUo6gUqmvZtHMPlqRrueYEOcwNAyWm3ouJQOczUK04waoTY79hwXhlRo879wQ+M3h0wjP
hK6cr3G1E6emqQV1mP/Dl9Ejkyu6XWF2KU724L7EnXl5MNb+CyvV0Ap5OPF4ovQNSCva8Vjfl+5J
/6q4RboN+ThA4T+ZBZ8l4YvaAtLcZSGCO4b9xbIigUVoGAmN0lvYSEUf6jYUskMeyKPoSvn25qH6
pMIVAq63ZXeuaIVlwK1ob1B8EF+v7tLKgPTfyC2c+G+ylie3HqCCiGQF2QnC9sh64PgLOklyWaus
xCli2ayW/qGb5MiiW7R4JslP9UidwOpV0OMwl2YXubrG/3LD/wg/+bYsC9wCid8B2t60gLls+owD
4QRDirxz5M6MWlH9v3u4iDaJFnBLmV8x1u23LxRLWZGadBoZrWtjm1A27QSgyWfECG+Y2LcyOq07
wJBexdKdPOpJsNFHyN9SBxgpRm7oe6UFkkpCxsgzcourKwICpo3JzHimAhdFIlo5xrvZIfn52+ca
wETLZ2/WjnWnxcTLUWZSLhfI5tso+bJg1/8TVSDFoV5x7OsfgDems2DxDkIig4yt33nAqnueo2uS
RTtvR2JFYtXi4KxkPGrHKbbpD6gEbZbNN+7MSl50x1FSOtNCNAObqaJIQvOspWpgb+hahfJnFdsl
QZMzz1HEp3VQSkvE6Y/NnskmI1JT7Dl25gannyuoQBiZnGTjIHVbs+dq9XhIypIbWaJb3YF9UQtb
VRoGVlLDV9fUMFpaCSm9x9IT5zd69Pha3yPVg2AdGY38/m5rLJIIlol4sMTn1aVy8bia0rp65Hfp
3pDD/p/tq5CE617TCyFULl5RO61yRN1JY/FncaAsWtlv3Oc9l3fU7im7Ch0NKwi33/FoiTIL8c9+
7Xw33FZ2cV0i4TrJkPxldYkXqux6I81o4xLleLn2Mr2VNekq2ZT+jwzZxnBVZuYqXHTTz8EAD/wq
TSxiPaAQT8ytKkXItmJIyk9kqSZo316Qq0JBd2NUEl/C2GT3+x28iX2rw+32ThbDuHW1jh7lK+6B
eBz/15nv8CmcWrAJz0OHJwPtKipQST6fS7n2CqFpvImaoUOxJ2PVPEGXgbrNaK6BYafktD0EPJLn
mlqKUvejb+m8ivgvtctqld41KSgnErQvZxRpOEiHtQP4HDg++TIRkJWz0wgDg5MboX3cuG2ibJ3a
RnRrQkWwd3DFnERj/hKEdvTqp9CK022R06zRjktMto+s/pdDGiHLlwq4cn8TUSdKo9c0Pa3qpagr
yR85RrqVnmI0RiscGT4Qanw28vLCC0tE5JQWju4tYoOk7jajl8cnXPdisNmem1JVnEk04MGqJJCB
TVkUTcWCU20Ol8j3Xe8FvVgPSfwAZnsSvpS0kAmpsRjxSR9BWpmNrOzeNWfHm+TeVzk5HZEddeHD
evwkfRz88s8G/jQsS7ZjwLBf3lZNHh3bklkksvOrpiOwmRo8JiXnQabFrLYsGNNNO1jmX/GTv/0g
QX87NqZv+p6PrZbime3orIS7SXmx+91740SecdTMJSxbKZ5xL0U/gxeH/Yf4/Uray7v81BgPMcmz
7rbyuEcSVD8Hz8z/EE3Nv5T9ktDw1Sx63FmLItE7+dq5Qp/5fX6MY8haWZ1g1QNcE8gs9aFUO7DW
NHEPZ+mkuX8Sbe/xio11oWpXPXaWOJaiJKGf7rS/e3SAMcF/LUz15MouJq07lZ0xZ1xWo/JsUOfy
PXkqPPZETxi9KWmk/Pu0VeZbt1L1ic5roPRW/Nr48iLTNboSMWmpDaEQOuzr2kkklTFMlbiNDZD2
b3lKBqgnqg1/fs/yzjb1iMz8/3h+pGAxpAIWpJuzMlwWmPHg1za3MV4x+ERjj9hd1H0Zst8xROVx
BD1r5ErP+qp8GEba0TKSbBjgVkzBQnnAQ5QIA1g+gD2qq6tDqoktjj2IkcupwihrkinFHJGeTvVF
+k+s+jUfMfXfnQBeInB2XI5MvmviH4Ku5jEs5EJFCahnASDwCt3c5Q3WiCWcUnVcVjg7+opJgTXZ
5bX8eu6O6F9+uNPOrMQnzVIg1vtQNYvcC6MRwhHLf/MmGVz/t04Vsn7FVJd99UkTPQStO9petwdZ
iLzkz6HvwQDycHPpsgEJ1EtZaMzMiJFvj15NZXSbPk9DMIkvgpAsf7lIXdrhg7+mC5ylmrZly6o1
0v7a4vVwbE/K2/LDVVgC7c1gtKk9xf4s9mFOYpC5MjEAe5fz3lvrpLUSwy8Mifs7RJ1R1lzm708L
FnbgpvLqMcQGrfZ1bKCfkgf01yUU2omZO5kOioKSsSQxoxfLLADHkny7snVj9K9DbTM/5ajAyVoQ
uqqNkxkp6gA5IXoRbtBaG34GTqBdeLPhLN+5qYQPYDsRvrOn1ASafMdSrmyLG/GFzbFPmfLsgUsF
8hkqpeh+cQL4YfPwprqcmJVrwigI7jWxS5P6Sx5wZikprI186m9dKNGQ2Hzj+Gg9kqj24SGPpF+l
tpA2zNO7msfUD/7rDUaTSfhryZOBpM5ixykPBC0EoUbc9fXGXQm73GyoZDhsaTsLyI6Ip52j1QCi
5TAPzFvUj1EBUCJ6cJc+L2rTwuxlRnigRNgxHKnqF1Scjq7pOOiv5YuTYxNOIhhuGaqP6/up0lA0
xPJYKjXFn+y5oh/Dfwa6aYkn3FKapfX4n5Mfhdisk5FFIyQjDJzAE8s319RdWbnFIFLs7eDHD2R/
VBqCcmwBY/njJADDzLd2zj8LcYITAze/98usQhJ0h29W6Dt8bCbHebSvTzaT2J0KrqkRTbXje9V5
KX+ZnMht8vGZ2T/yc5syX09B2x9zKCtL2Rf+UBDtWtuOmJ2rJf88ZoHfIZFsOYV+QuZvSykkSslc
WLb8dlTDtcIAZBGi9mkMPeckiZdrwXlqYWgOibM7FfKVQmiWCAAH6Lz8q5bnUaQqs5h1VMKleu1a
GMDnRvWyxUg5bS3yG5tygi1+788wYmxo7ZBczU5kBOAZUXuvKg4yCxAFERbWcReSfEdHqyjGPnZ6
vGJaAXe8Cc9x+n0gNKHCk544TOYzEWGhgE6vz3hhEedqxeA3inW3m+DdxvTeD/KKh5OZuuUhMNcx
5UCZi1P0XR0rbB7uIan6PdjnI/pGuTYYK3GXK8GmwuyLEWICBQycFvxShwjbcFytVFsBQLJfUewH
LPi1iQkGelB7Ynnf2piNmlSkqUuS2VcOu+ogCp3JzOyTJLHpAUDKLz58LbeOd5V+OMPi6neRPMA5
1a6xPn6Vq/c2wH1Nj9jecBT6ok0xRIK0V+63idfQhxkRCyy9HCZ7+lCjysknwRiRTAVLjQo6V4ag
DoJJngfv56OEdOGS+08RgB9p42sDJlU+bBMSh+oemnd5eEZyHqR9ptcV3CaK9rNd8xSEQHpewGFj
ll0/kNQwy+EG0dDFLPrSY6vE23If162EFAwsSLpvjVbiiaNRBU49For4CjhQb/Ne937ZAiGGp1J0
4ul4FNvVYy2z8pSAKl7IN3pRxWos7WDD6YXHK8E8mZLbaXLURqQjcBumpRcqRJ8ShI3g/mZWp+5g
fM/3i0LNvn+2ndjUicHJNDNezW6B6OIA4i/C7hv3wOtb+mT6uAX5/gO0bTXJd2xB72izeWZ7C4bX
RuIfQfgHznXBiHmG2HAULtWFHDU7kpbgdLURKs3hmRvzaiLTcdGihb4E/gG5Hy44E/KXS7cmp5+E
XADqlWJZB7sxfnEGkUGio11nCqyTHQdfZjwaB5LQzBCMzYMEnxMcrqqkVwjEGIwuivEm/vTHflcO
O9yOdYf9tEmW4FKSWTbWmiTGyjBy54sq/YTvF0Kr9+hRB3JSNEsDIYMdcswcnPXl16gXppJ5mzdK
wkPhiILFFf4r8jUcXgOibz5Viv5PBngs7SQZoNv3DAJ9BM8PvfTA1by94W4CT3MxO5cTccFX94NS
YJec7PEgt931/KQHKDBtwviXZ0MyHjFFupNU6gx9EjpD1btzx9812lnrOvySL6N7klHoQuwEqFLX
2SBN+1UzZHmagb0OQDqhMaKMA3bF08TC7TDdnCX7qZxlytOV7YFT3bywQDmB/nqGQh7t+gTlz1Gh
kjxI1yngxeQwKH/vr9TMWfx264ndjJPeRZoURaccOOTwJyTjdDBKR3QRbwizVij+06Y5tgm47VPV
OGpn1iWorGqjxmC+RNzJ3jfmhXOtLXAc/KYXI/Gk+x/YRbloy5MF+9kGCwXcM8FQLxrl1nsAl2z/
k+rX4Qr15/dpDXj6XbaFDiONPZCfTMHo73sNVdVGnBvgCwerAbxJbtt23eseV4FHghsk4vjLwc+E
LZfbnoEoPdpIprE3wzlofIEMmT/j8lOg2KWDadMwvE65dB+7X6CfdrL6QbQrS6wWnAYKjtIsW5Ri
TNUJG6PUjIy9eTWT9NFzfraVfnEK/V8xNWS6JXwtBvwvM1jiko9tT4wq+tpkXhIJO/0auuAS6Rjz
LZQXDhf9TYhW5mrEXXsff6XYH7V7F6LTOLQpUxljha8XDDqjfET0C1tKc1bAnHPp0hxldf+upHcw
k105ucHk/xdLWoqc+4b7SUTfECO2pmqa7p3H07k4+ggtVeNl6otKbH3QOLtKixAH3ubIzz8k0Izb
nc3/E+5xD1h+ZYF7GxNORURlzJs1GPTGQcNIJ+7mfz8/3xU5oYjERWtXH9H9zI6iIXQ0cHxFJVB1
T2juoVhRXuVlYZj2OQ1ZGa3L+wg+jBQSFMIRzv3wbke6c7gSncEhUUhKhSKMkn3ZxVOkfj+HSRaU
2J19/cgze/QI9JiEmpvPkMDYNE8z/cmJD23UeaoeuCeg0ybRDB5i88a8hscYoiLgr5gyyCPmVFqI
5iOpvNdWkdyX+NTyXQcdyWh9sAb8AZHqzCCHPHjwcI53++HcCV6+jdT73R4m2vsfPlVoErfYg0Mt
jbwew/IGfMkjeisSEiJvKqXph+/cg7sbAQmwhlZIPPpRD5Tgol9Sul7Y7cm2eVT55gzwirBomvK3
XfrFnzpS8MYY7gx056qHHak0fvN4GZaMk49EUPZkQfhQ5qLK/JvaxB/vYs226KGKPm+3OHvvm25v
JQjcX/xGKsOgHLEWTUdaTEBW143D8z2OWdCTYvt108WcD5q791P0PMkKomKjtQqE+0VW7VY8iwHQ
XzdQd2QNU06RanONzak5WcEB8jIo2Xrfw+Bq0cscRSvy5oOXPJVzI5aIi5Xo2GX2BvwlSfMc7Rw5
ILKp6ZRH14JRd+b+PkJA8kBOJVEKkZHv4A93UwhuF9TXeTZLf5AIAOVXMZ5LPYiqJPyCWJMRttb1
Y5sS/OZvzOe0hJWF3+TlffIXt8Pk+WVyOSAKcDHzAUw+XoegbMlHrQU/LegvRHnP08SJ5OhpWiMz
aYgIY8/DWUAcaZY4kBeIJSaMSXPp22N20vo5r/Ndsz9XsdaKKLf2WSDiqeik4Rp16T44lbKRdqAa
pqW8Pu7WW2vKCwSreCjbZitazHjiLol83R7cQc/slo5HCPqZ8adUYO6HJqVp0pZ+/xhskrekNJ4b
92LQlx8s7aYkZK3JgA4uE7T6buifeana2h1QxfSZFiJ44KUqtqF7CmwNsO7vSSNEfmFDSRa14dJn
UMbJe/4oAMNVCWgGvmk/4L6D1AnGcDvDh6P88htUlBuAnP366R1Skuz8keHAWfigJmIEjMx1OdRt
uX5W8li4Xhuf0C6S+yL4EkaMsrIwMN4IH0l7fFi8ZMvjmuEsHcmYYphigsj6sT50K6QLG4LIWk8M
2Wo59d+N9HC2R0UzhqdVf4a5tu2VRqgHyoWqJxp9yS4OkgVfC0vN6PAiTt0oC1mtgBSFhE07HACL
wGkj1WKnfWi3ziWn0Ex5Y3MfG1qX/Zjykov9XLzd8bHIWAcaaggERUOSJs+2nky7Web0+A1UDqnq
vPAFNS9g8TQZ8A54XRcbajoPpd7Df993L0siMrgk8h/YL4kP1c0ffte1+Zt3EIimgpNOwdRVTZc7
HYNObbPd10Z7A8Y0yBFrCkLd3sj7P/5v82sSLbAzX7lsEIYTfIZNKzCihQz17AU7eO8+meZ+EK7C
082ZowxeMDAU7j+yNnu5czdwR3XS8PTESM0mq/U3knws2DAiEvgBJPciX3uwOL0jxc2hFU5EBYEL
4vLEt34S65g+KO6Ri2z9Dqk2ZZ2fgZYxDyYT9hCteZpjkNr+XDTFxaLFFudIXM7uNThkGHeFXRsU
sIhaZUk29E4N9bRXdm3kiUfPf6R2BJc+HYc82ZUOI8iKHwA8DZUK0JuflIdQkZy9XqYEfNrVSP+v
X4ILumkjr+WQrDjApIjf/byIl7VlBb/xhcWVZJa5Y5F1IZfSovjkJbqEhmR/aIEt3Rlzi8rbbpRU
taihhLH0HmliEWlh+TS1NkxjxqLc328Vzka7SyO2AsgluGku5qCSgKtWFSuj5PEtITPmo2Qp+rsd
4CNn/ebH8uajhDv9kF7g8NtUCVFL/Ve0e6F4jMfLQxTvpjoTZn0DXVrrdpDBjKjMKyru227fmDCf
FqO0tmsM6VLXx5PFxwnN9IwVsxDs0EHHvKnq1CrdZlqNcAO8oNKk7uwmsu+22o1GBrdcG40BMKJv
9OSWXXPHT29oa9w+26pzKHiHJCEIlXgMfMNSc3Up4nX5owB9kMLtN4MneXcTAlFR/Z72y/jRNHIE
SYtF4BRe7ftIbOu7aPMySxQbYin+MsUGqA5s/5FNVhHKP7fwiY3SCZH/wsPA6kjccmkGq1ClGNSM
6iDKEjFUeLE4+iy6nLRt82DVBeSWpTkHuAlJAwdIFS6Y04gfbzFAe0F8Z5exZjd2sYKXML7HRQjB
/OSZUwosksY8hoiVQIUBMFB52spXuUluG4oHYDI2MHx0SAV5hJgdtTkWge5+fV/OQDvWgHU29BaG
EbgOJwIE5tvqivSCzkYSPEm+jesfgCMkHfX94ALvcis8dJ9yf4JL+HD+ZWlsxx3LcU8AuvFS4J0X
EwvN0l/8mZjRHIkxUFZvUqHDQg0TXHwHBbjgUXMTGQVgF543i7cCJMbhCvI+7CqVpvf7eG4dw1up
EssT0Ba9bWZMDPR49vI/UTOziBk0eQQse/BfH5+lZ0FzL8Bq6wtYEciIjxseSe4f0EvOscYQdV4O
O6xz67VMY/IxyLzu+LdwuZLFB0/vD+LT/KYtuPic/LYejkkQJ+fcVKgGI/Xmk2hsf6pK/GEtQJHy
RCMWcey+zJS6jWonQHEN3I8hwj43i2E1KRN78tW+rmf7PYTfa6CFS57uKjIj5VmzBShet9eZOV5P
QOIKgpGFi85AOIEQrtayhpNVuIIaGc9TPv/2XXqkYHeAaPZVGO87aA3DUvUO4SGYhzB31PRjn4IG
PNpcWC6L2aijXA0dkN7Mxs3FRn4IOBTAVLoGT+EXye/jE4t6kDOB1pEdZa/P4JkAR7z3qMgQW/Lq
cuB9zkOfYB4GyjuHmynvuoQYR0Jig+rn8gY+koigfMfSKIS5IHgKjMDaFLHvpQhMXsL8hdxyHTlT
EguQMTkH9AhbOHtJ5FlRkS+ligjbNydOeDzHhOLvxveAPVVM4745mCXhSTRBJOHgKLMKSHzWzR6W
X31oVjH5M9rTLijymSe6v5uFkSJgKM8WCsXHSDz+yCfIBbBIfMeh+atqNQMGWZ/1yVLRYeOQ7jVW
13n8Puz6U3Zwixg/7h8lEMR2Ow1pyemBPC8zwFGvMDXC3Vvxwu16FYb+cFej0aTXftNrUA/s6kJ7
HRkhyJjh9w6/qHTJ7sitmTw0GGIbdFDhpM5TL+ysan70LKT8sYQTmQfbwAA03Kbz1ZsgvqQ0n+RJ
qt/4zEYK+eNtMV6BbxcdxiTGOSQMB09DbSVmwwnR/+datcjwiB8dG7GesZN+8BYfgkAujhY2UlW5
jCW8L2hyHlXHfw9k45gx+BQjxt0ZZhxfUzMl7VYXQL9o4HbxS+e5FGEO0jaK/P6WC3VnhTnhhLDt
DNSGGU9QCk4IyuAw366HxwHdACtIeWTicNQ8qe+UthSiQ6wrB4Zvz6tOuigSj2ZqxJaaddXL2ujv
0VvIGDnfDS5wsPWvSkSJPM5OvkqyPnqpIk8/87p7Gzt1FzKoycu0d3IBns/kRPFtccCU1dBN2eKU
VwAC/ZDJyUdY1IkizK77Q8y21CLyzvB3feoT94t5BXNlw4d2tZ9n0sWomeTlGbRjZtMDGAb3d/F1
7AMQcjB+Rl3sg+F1WHnKNCKnJ9P/FJzMCW5ffFGLx9tvmhvoGTuaQ6ME58O9HTQKfMPmb4k9X4Z0
wAQPUrgsOnezCg7w/rjl7Z/NBAQbUmegUxdfLo5fI6xGLtcV4sXJmCcNkL7ZYM7qRi7zOAUBA92T
gQaeKsuMwGr8HG1l9QyMmVXAhM29t2Q1noKLJWbHymQ+6rT/AkvE7wklhQB/WHZtlhw/gROljWZG
pypwFnvkcKMeu16No/E0xdwqlAkbdK+/JQjeRVhfTg+mFMjvxrvkbQZD//NZRDUee0tkeRYfXXiz
ZD25WVuelutEJiRMzIQc0W22kOGqkXz3tR18d/0Xh6PY3Qivl9VVaX3WKrGiGDFcOqRuWjufc8Lr
0/8LYXspNosesRF5sMtg6SMuz/SA8dcUNIG3nn0XbY/9SaBjhgh0c0wy56Nr6M9+dTvizIlmXKjk
fV4mASUlY/I10doUkayJ3Vr/ORpSY2MsyaZG3/N5CnUyj/Ns1w6Flzj7qlcXOyxnfd+lhtjaCthb
5MiLeDskaZvysZt6Wa0WRo6btJshtsgSAdWOlqYseWoS3tWaNbJc1Bh++aVCLhtN//rVQ3q2EjKb
r3fLeiyqufgGufqxsr7X0iizRE0heD5qYkOCSfMYqHWbjr2eD8vrlZh9+IQeq6Fk39PnruVM++39
0HQ3vmuiyZIjMmDomfe7uuA1VAO9oKYo6axMehLxH0U2eSftqzZH/oBsK73ELHJGVlDWdpTNdEGa
cVy9VWp6kfbxtKsF9rM6fzb6OGEzDjQDieVIpVpeVOSmjTHiEaZzf/EWVnGQlgvKN8CB6gpEgFFA
xgs58fOtmIlM7cZsMI6oK51h1e7UavnSzwNCQOPjXdaB3rxoVuceR7j6yYwQ5vozsKZ8HHVwrguL
FBphj5XnoRI7ivS3tk/bJ2Jd6HpnnBAFG4Rngmxqy6pqDNrFwKPaxtwIryl0P5VzFDZW9OmyZZLd
XeIe2TQH6j8XP4KqymmL1DReDUxAiXviVK2Czn8iZ4UcoZe9u2RkaAUjlJLqG6rcCITDrIELEoAT
UXJrAXieu0SCXjEXKGgYdgpOfd9sDnoiDI2KYN80fOrYrYUQEp4DmA6jKUZkS7XrklGYahfOwMAA
w4sm0N7aSN2hk3tiM/6bjqloAgYwoB5xQ7ARNcn77GPB0slmrZjgNIqDL5CNTz3mMMrVo2NyG3Fo
0AaqL1E3V07/MunLbCe3jIL0aiA5HajDWAgODwJtWEEzqCunJC0EeRJw14FBZ+Y3uSuhdwMNjwU4
Kc/+v5+dcDCEepMBdqIPj6/u3ZxfB2HAHzGPHbUNCh0EZHAWVm5sLTqUJI+pbYepOXAcGJcCjWYb
OjOOsm2S82gVCn8SsTadBNbj6ythp5ChsZeFSbmx7kwcWoyfMcCDLe63+mrPg/4/1KEDvAiUUdfe
C2bPD6L8HQSW4cpYmbeztU+T1ZNdaJaSEPcbbqDajnL+jUHq66udgzWLjDhPeeWPNOp9K4ouWvd9
s7uU5qL21VL+Aavk34Z9CmjMyoxU9x/wVGtCcjqCof8sYfvO7AQ95+2piEfqU8kNVh5qu+nrp6TF
yxx9/PN1/2mD/sDkRCd2fj8YteRUDCFr9rTnZBPyxk+k+AqAeGjdLkaC7cpy7SVlGQeSnoxjDwnr
2H7dfgTTMmu70bf3R1f3EHPpHfaGsGiZsFPatAeGB6B36M+LFwGlcrH6gRBhnhC0tI543Rjscrei
NOFU1Qtwhh21L5JlPAruSqRr7uFb/Skv8wrxhOrusSqC4SqP1d1L7ZnjS/JP7NrEv+kgvt5iUGVi
eDogrrwD4V88EdIoIglklFPqa+Klg01ftiqAeRyS/+PFfRp83YUqZRb4oKrg3Yo54Yj6GY8xWYTo
IQU8bDvfKfU0535gw7sloJijE4wdOqKOW/dQDJVBVPQXXflNoCiQvpppsy5ke94iJT/GLap1mzC9
8LVr1tzVsjGfK5tBqPgut1+OWYdXDYkVNP9LeBK+efGHUnal1F7yhjtU+IypXz+Z7UKj1/JaRb6V
nwO/9nlYyPGskaGNHSK6I+Z32JE9ddWAntjKE603yAAt4g60z5JgiNKJNaOhTQY7vLSbre/k20F9
o1gxxPsjL6JQrlc3ZzHwVO8YZHpOUDmKK8zL65aDBsXapPXYYLShtke75QNSxaZn5gVGQWlXORzC
mjyOc0/BFSv9+VSUb4WRy7Pik7nTqOUsLuk6wMp5mNb7qhvy3mWmIJz9S83jqvnosVYz56t6tkH5
5gkDwz/kxSdA9IwkcTGG8wTQ1cr8wKbypTF14Ki554dI1fyxNXQML4zVhT1FNK8rIIk9nCL/TggC
LyKRM+U15ZGOrN7Uc8nxkpH3bRtAgNhAd7mGiguovxPsKJnBnEj0G4ejmk+aJdDC6dWizRVUx+2W
7UIgziXHmTPztbXijfskF2DaBBvzN5+/QliEDdeyOtpeIoNg4Z4lj0aeGHACtDE3M4tpc8iYwWWF
FfHzRui2iWoxqfo7Yrz/ObH7lgkdd6/Q+sW0F4glKNEe4kkIuD4IkV+ekWvGO0SXR1NDHN3U1TCq
hsqKyu5Lj0CRdnWE/SLtGXaoMDQ1Hd3fa5v+H/U0Vu6ehfbr8hXZ/DY6zuWUjiQML1WsC33P+fr/
Q6Z2jZmAZl/M3YsCPFh04+hE0xfCaKKqoIzYKX4U6gVvyd/m+s1JYMohBLex/+8QHSnoH7ShGv5z
B8JMz7/QUIfXUnxFNbrTW+NU8DE3pMUK0eEG+ghcbnGUp2qBtHulQrCeosgFCk/dya//zCnrE1Gl
PAJt2umPTBzhtOzZEril4sM6TmdJwB2NuU6w+l7D4hq+nryvDO5Ezm6I66f9XXj7rZ+Yn6o/9tre
5SGnfplmA1WItjTNJeoZxsdPCwpPjPPAZ4d8vyjZjQRF0Tz7sb1/H2G6tCXGASQswUUYh2UBtyWC
hhWxdg8vUe4mOfJvkTrGag6TeMu+SaiFMeoQrDYgN72Rx55n5XW31dolTQt5l/WQpoJibEnU5BGy
yUTVYP3OELE0yW3rSQpKH9FXY1VEJq+M7f5FwrfCbHENvhQM8OvoqG+PcP7zL9zuShfv/RzgNtCd
ZkD3TPL5X3dCodHPzcjjfWf7vYY+DYyR8OQeQGu93hdUVubkyUrVUUqvPXWzd7R//k1vv2WRE286
8/exmO9YG6xphJDC8tA475FpqgopFM4thV/A8emOUGxG4MlqDrf5J9MHjv+QR+BUhbXDC0GQzyA2
UVTJezIVAjCwbBKXiEwGiXn26qKVUBFCqtHNCETEyPNQCudcegFePnTUplWbx4pJ7abJ25hFetpX
o/+zvqWJWROlGAnzwr8QqwKyF6zzj7e+NQF4ml8Hb7qMmjXpt3CJ8kgfeXCmSK0Hl8u0zlxjOpkB
Gu/7wK5lnKE+PE0MxbA0qKXPHsmykOgrmAwC7L9URNTaCpD7p+K9dnj48wkoIYKz0x+A5CImbRRm
GKFvBqHBmtuHjhC3mez63jkdJMi6OEHqukZOVbKcR+/P2JRo6/cc+/a/GHK64lhxZAr1AfPrSwoQ
m9NhGx1mCjNeP7i8WMFDFTodYLiqJAkw6gvIBqZB/RJcTfbwfyGZUaKYs7ihGuluJhExpxSbXB/u
ONSzFSqhaEV6+ICIXeiLxSRmJIlHFkus+cXI7mQ6PrI7+6zDZWPtCv+chARBWtS0Qv1B8RytB0Is
TWTVw8DH0EGIla5IEwY69gHrfAHW+WaYEK3izhkzDhzNjwro7CKS2qrxmgJ18VA2t1Wev63vxOx+
4H8QGLMTknhLgLhllBpuT0ZbuKY9RiUOcZS/Ytnd8Q8g8xWDE2KObgu5r+XLT1qUbIkWjQbQOGkm
3N+Ig6gvSRlFeg0lcJMYbqSJfU+TYo8oK9goou9knqfBTRhV0SUmtUISrzvARnMouWJKcxMyjdgZ
ZT1gHLlHZo1bsxmXZQXHz2XGXI1n5blN0QvuuIxNsHaPGWy7+JjR+g9svhVPd1GA75O0Ik+M6r6J
EEyL/wLDzARFo0YNi7oo82IQYVE2g+UCMsY24S9y1oiCNwS/hpF/maPuuhnjhsnb6aa+ZbeNHAFA
Nlx/CpUU6hFlye5ihnQyzUkt/S3tesyBAkhwFS/38057y4GkRuIeLG7rgFG2tb6xk4Bw9l1ZWSRc
pre0xTtqAWnYQkuVduNhlUFEaiww7PslBK34tj/BMj+N97470i2s9FDcZjpf8PTesDBpl/uYxFAQ
l9HHOg6m4eWOu4B/CKe+BSOL0WSTki7skogaKaJM7OzljUDK6sq+Ofx/Uju+O5HKiLLZvRPjRvRO
/5oz2hriZk1ih24ABcEKQLkJama96IaRAm+QqMqwedc799nxEgHtEynvKrxNjJnOYppgmXFvDfeu
bYgwZSK5g5th22SeJwYv1vMEXUv3mB0FdNvKYhfXbfFLQQQp67vlkmcWk3laK+l2Nce7KgLSd2jJ
9po3yTbohYD4qc7Wa8oCvvNqGG2kEAVb0WExLe/1NLs2ZM+IidjD9QdagUHkq323PFEANi4IZFkX
zTcnjHqDsIP/viBW+MQbdM7l9gEYe4Z8dcWdYqGTf1Rr4pmSYh0+riC1I1OwcSryal7TDFveZseJ
xIoT9BRoQVh+E34fELJ0g5OXFcKbBaxy7diACWDtOXQiaZRtflCiy2lA0NATCbcN2LSfM9HeLPdm
ld35iLSvcMEzahPvDyaJSY/+PnF2kkDWXwan40/aH82c1KU+O/74sRoszpw6K1+oWmdQAXX/jVds
Qp4HdHa34BqYPFKLPLfaP2FKR7qXOYoMUs6g5696Bnre38IUDwezQmhAGBfC1l2syMkVQYTk93j2
0IIBQJKHWOKExPMkFuc0rAczBx8JA2Z3+VAeJ/wqMVBzdOdAyKEZNYBYg7sH2wHnK0ib6zLf1JYb
tvN1uCba9dSG+AKXb3ba+Sx/GTzpAoGfn4rKXz+A0VUMUwbk196Du7RfQVclVpTqY8xG94QMdMr/
64PAafrggZispjoF09qIrYp+lR8jx958jy6kv2zRZyRPGDagrKq+/plC9K7CJYD+Zd8mDWoobXQz
6wvxR+DSSoPFLmmLTqpRiRUOi4sSdhYdG4k+GTG8mdlbfGkW/BPtBeFCdpMzSopcNNHdKudChwPV
+t3+RNAfhdMQCMfzBuRgp2EhgiWjkAx0PbTAbqdgwOH36pxvouuwUmLqvmqFFhlaYZod9ONm7qIU
Kkky4k9jBucJgsejmZ9bDl5WCAXCViKZTN/bN3lpYnVyEVWzWSVFvz6WWq222CkreR9BK76/KxIi
ggXL1KfCLeRZx4amrdaemxxLDTUGuniwegPj0wTPcbDqKGRZc/NYga/V5zZULIonB9TqmY2jIH+r
62PvLfQhBR8IAFBPaDa+vgLSwln95Buuuw0S6zMVvW+DlNoxe8rFocYxcJjRMwimx7cmt+FP9zw5
3uF9LC5DFowAk1YLNbBY11/Iek1AEbbB8vU6AQMCSxTgdo5zoM/IuGjy4aYvpPTaTrPCRGvlEWTl
HPpPz59TLBAR6bedCT53CAHuVeKzd5VLSFruVSwLLwgtK2qn3KLVTHFtPZ7D6yv4DE88RqO28mo3
DTDmv6v8qTQY0jW9MWOi3nilezeKI4SO54G/km6EJw0GZgqYAB7EF3d1UqNDQk4BaI97837ST7ER
8OrB78iMq3AkdEbfKN0b0ofXMUrmQme0wByVL4WrU3mXFy5eGzyMNU8WnespKdGCsIyjOwzAQa0e
t1xhi0fSO5Os4uVb4ObdO83Usl1PTeLf6Bx1tzLxAw9PcOTldR4sxc/i+PC0CJnXoX5qKienB5kb
iAcsER4SHJGqXn7eodASpaNK8LeICAIM/e6dr4MdRbh2gYHbK5kL5LHQPvWZdrOZp3+ig1ss8EDL
ebh/br7IfuFLyCOGXlZCU9L5zNua60jU2/wnVBYJd027ggsFm7B8qRMtSe+Bd5va4Uptc0cn37FV
LUb2nbfLQFkejVJKzW/tyFER0rR3OLXg7WPvLxMdpkX+WDAUx/7MPgBwAqPzOiXRwfFxphvTKdfa
U5INZJkd57H29h0YkWFpdgl07KQ0up4CFN9xzAxrTlmp0YmukqdtGhMoxsJXcqNvyUHuOiqol6uT
33KbQEXCpM9BY6XCK4rOuXHRzZtxBhnLTCsM4E2KolS4FJgQvne0dKci8PE9cs4aibx7J+hJMH91
H5pu9mG9hTUvogPmWmK00FSbrWhWxdQODdbuh/rzBCh5BpO5aKuDCGToFcWin4XwoWU0MTHXYwpF
N+3AUMn2/JgKJVy0orw99DVNgbQihT+OExcYTNLSmtarwQH57h6xVt8MnTD7P0PgM9vVi28bWKn1
Iba3vBZkIs7J/eRRYpQmz5Fee5D9XO1IuzWmSLXg6bZ2Uj6wAj9Szl0pHhpgbyTQakcalbdn8Yo9
rPbOUsF6Cke8nJNxIj6tLM2HftJsLQpLWP7i4Q+L+8wZw3nUVu5wWiAySDVgpgp29rtECJWDHe6/
t1NfRhlloxCaFogZU4KCduisJOs9N5Zh4bzneaPJEemQ16YL1ldoMVuPhgiPoymF85ofCXl3Ssfu
1YG1AeYMxZBK2kKIraLKqNa1y7FEzn+B8wrKTUqfu7LB5l8pa8Wt6g8cC6PC4juAnQlsmJLZ77Aw
AlEcrLcnVbCq3lyGo+m/cddtbcLFAt8U4rt4GbUVLV9a8A9j1n+f8FLoxb/r7XXUFUw2YXy8ssGB
tYmW7ffs8Cfe0Yni6x9F16p6Fz2iK9dLgQY7rdHQfQg7Lu8WFQOjn8lRxK5IyehblbqcB6NqYVfQ
GyvhIZk2XHYpwKRskUsiLA2pMCowa8L4qZTaJIb/oyJWiWXdHv256d/lK2EupxHyCDDAwZLIemP/
iEnGZlprMkmzMVi9aUQdffOJPgF8Yt9THVxLHNObd6aSjyB35EQ68Lv38UJ7Ssx0bNm9ENojxo+O
4Gu7HgNSEf6UouLCcu01x3WihenJ8Eiflg7PN9yYNDX1hUWmDXKoTyNlLB8yMYPhwgRysxIPTnlt
n08qA4lwOjHVLKM5CTKbplAk67ooUdmCLhYs8LgmADYo/xWgL/t7LuDjMo+R+H6q5X+trOfhJ509
N/NnF21CVGbGUZlFp6N7jILJOnp4MTogormtHuKadKyobicQ4D//UvzQXz7HQ/gWSHu3erdOK04h
vo7VG/sA47/1uqsg44fdEDs5CgvA7uxYU+x0gS25/OTrLv5zAMiSclUPMXUEaqmjy3sAnjQ483KS
47G7NSh5o0VF/9skud4qIy61XwAoN8ns3lRfOEbOCLJpT5EYyFJPmthD9YNaitQ59H4qo3Wkl/8s
GUfLG7fCnaHJ6z1IXulx9K3sBezxS4hxnchaB0Kq4dId20Y3tTPgXMqDDaLEgHinULXR7zdVpZXl
kQ3SIeUhBXtyWqREr1Z4s3qqznmGEYfWCjxz7MUWiBaby8MXqu7HHiMiiOdUB9ej84GO5A+hg3ms
BakIy3QuwiihINgoJbdPlhniXTvgzGToFzELzaFw4fzk2iiwiiITjJlUbQF1+ht5JPY+kn4dawpx
qCMmhaKFeDr5DHGTxbZcrEA6lPOfJ7ntbl/4+1YWiqU0XSNQ9EbqwutiZI4u+Pw/XnTyOWpFnnqo
HRryBs5mGQfyFt1MO/TqJKKLyz14OYm7xgV0SMIHWhbK58zCunAd7SFBs5xZ61Hn3pMNIhVWS5kj
OnhgFtwyk6fg9lI2cSU+u+7lMxF2uEFFD3enIKh38yvTD/fKhNksUmK94Cj98RnIXznzaTa98KVp
oSEfMhW3FqYk4ptTD4SYfTSrtm2Xle5mAIey1CEkOJrUj5YhNncI1/Ji23aBU3gqu0NrFT7Pycbn
SlKtqoUNqrgxdZU1ppUGFdI1/cL6IfDrISnisR+0PHOmu1+ffI1syJO/CEayUDCHV/dr1jNO0EqS
C7QKGWLWEd/Y0psfrWu1u969rLSZ4SO1qTXYkfIFvTqLIaiQn8w8TGyHlygi6yi4xxfcNl6LrzOO
9Ke1VAmIb6Chhx8Zt6+yHPP4GZg3SEsjNvA+uubuhSbgLyFdi+X+iwfUZxPS0/as2g2+Z48v7Jfn
5PYs6ujzU8aO/8bxjazFy0wYg9bnF62XlVmjwcvXE1/+BRJVx6zg7Bc+QG7DdDeTRj/lUTy5sWN1
8L2YQ7fQ9l8FR7aaz3nd2/mxQ2+yf5eQLMgnMZ+pxsr3JoWGXgAvINU/NVyhERUudTNjqMj0g/9V
ye/uEqOAJUP8wHxsTiqbfb8sLVkZ+4lenY5jT9AzfGo5XthBh5pj/DBNJtVhsJ9Y604ZoKCmiJI9
5cIdhYUDABeeZBJnzvRytSrP1QlGwzQ53QolDNqrhp7CVODKUvle/K3FHNBWnzujI9/isrknqQ6j
9Y9Sw51TAfQWOthntQIX2yGwEp0gA4xhZKqYSZXsN2NtbcGhnXQEEmN0hlJutbh1pvIPMir/+oAJ
8W+UWPdFfbcI8GdqMUTauiq5AX/4lYoZlUJM/KpVMADhIoJgB4QBnhkztSz+e5rMYrns/WnKQpvx
owB8WdPGnfCUXtdnHdeVYdHHtourowiZ1clMVp2lTkmZ/MjcXSUOP/cYvYGwvlCXiFIdQ4ac+noJ
nTTpR8Wa1E1n5CTaSney+EbYW/Afvo1wgci6CucixJLOg53QI+uTUNhIZq3eOZOyhd6BcSqHq5v+
fPS0r6O/Kl5cLWSKdyYF1a59Xz0MV232DIi/TiAVaHw3ZrsA9bQAndW4XXtX9cksEmXouP3V91C+
x7/M8BLsI/ifkFP15hPMVjB66vUFuFW+9GVdQ9+TEiRooBY1iphSpgZPitGkGBVDZcocbEqloGeR
/ec4G6VTjqy83EGZavUy4+nnaXYoGi0szI3OHMvbVrFgzmoX7dSmznHE7a2HwmqkRE05eBqvmwRB
Ff6yBZCx7kv/V2ELY5uNN9HqNR4+AE5k5zpxEXQzcoltuLgeaoOEKJMbdqEB8o+1xYnpFrgiwlXE
QihrRoNc9tl7csCUR5w7RStLSlozd9gca4yGJfo7Sz8OmTN+l4m2uGJf3/iRYJJZQCYAfVf3xC21
OZITCQYskdN1+gS2TE9Lw8IEn6KPz3cbCmkVOUx5gqzu20LaSK44JmUmq2bLDJOC3FyqFWRoamax
BXBlylvBB2cs2SuYaS/4A54u4cwqbUioJ9DQ5BaOIgfursdEaKkG819MgJI4C1cek7f0/mX6o/sI
RoMam7QIGK8qq6Txw6OwOYagfRvkvh5/3rdlIfrQS6h8Qh885Ppo++tcFILrg1e+tI7tiKmAlwC3
kT/K6pQ3fbEwTz+jOgFQql3j7UAC2PeODElZiNb/PeotQkV6ZduEeAg9go+0B4nSSIHqs/NMvOos
ejoz0vynXRVoZYMjC4RNRHNjIPiUtqM2wo+52IFSbUl8VjooU0oP6YhSzs1UG5i8Ks3l6DKTsM11
TzK7YtiQfjrhhtAKuLqHQ8rL5A3w8h2CjfGdj7HdhTZrDYe5ka/Z7sRRQIiH2hU1cxoDMnwhZztf
dkRJC0VAPcIlYqvEQ7iyq1fy6sDu7qCybDyYW30GPxT3jGMFZVk7lp6ihqffQm+NX6NPHWwL9epZ
D6gw4NzZ1/QDe18y0rDJQK7Yz6Cl6kU8bhKdO66iZInAso1ZsyN+lczn0YaqO3Xvzh8rJVz5Dv7H
CWX02E+z3YtY9zE9oJwzrII5DL8imo4TzWr4sAfKXWdNHcge7xmDuq9zZA4m5r+X/CFLq5gEARhQ
dV2KMuXNJlgFz3JfJ7UOwQz+Elmrr7UpzYoUPRr4gso79naUScMTJXAmZYzrVk1MY/7PEjKkiHv6
GNM/DVWUxssiQZAb+pom4REO5HR3mmzvV07iytWHI81U9eZjQLfWt7ue/A84ZYj3UadLkgO36G13
sWzh5vsY0oAIPLp3Ls0zMzF1KvYZ5vKEgHV6UUMuBp1Gkv7AAMsBkKzIWjb2BSjSMvVXJM22LIRu
3zGD5od3iQ+2ff+PeicM5z6e3hP3w3g6HjRjT8m6fm0uCXrnPB7KnQAgMB5pE2yU3F3Sumdd/Ow4
vTsUpm2IwbZTW4ncxGFBtDr/e32CXn92BNozqT9O0V0h+ny738mgLSVZo7cQLc7BOmPN/pULZvQ8
UKXkcYdjEu8QOyI/qZrP3g1tyWf+JIgZ/n2Ch9zzQ0d0eoY1J1TowoijUn7eZNPbf1Er7OrYtyhC
6KS8Tl56Vp+S45QBop+pV/ee9QNVYinAbV4yt+i8HyadUN1kTIhMOw4PWaftwqGKMd+zxmUQ7bne
7KmXmE2p23GMxyqQ7ksRILfsSX16vkh4vXdJugw1GC5F/uDxQDAG53C2JfeJrfRwucEYx2d/pBhA
cRvkn9oGV0xieljQi2cB0Cl5kq37rzjdGJMN1MYii/1QTCS7v7oh2JcGlK/bktBYbqcvI10XsROI
JbQNLLT6Eh7QbO424Px9LYYYBSKyEjvuK7lpq68VCU5ssVDr8xWAD1TiDNsUbsRyY3f1YE0V2KzS
aJfQiVBzSvaSfku1J5MgIKTbeywYk+bs9XFDbQ+1OobmLOpwt0cDblm9tuJfax/+vr/dCYdp76fr
ILqcEL8xFXvPficcQjBO8CE+U25qyvTsKI3WTRq3LrxwlgyccHfP/B/320slVGW3X5LNuJI43laY
aITNWIfVMGoFa3L6bM0P8KH2EKqFNpl/GUIk3QhkwXbJUkPyMRZpmzg6Ava4EYlo2eG7KePJe8Rv
9LBN/hArVvkT6iRiWialIqrIHc3ohNyATtcb+p1z8E69HyV0erLd8YQ+pe7hGbjZj0hBRjeLFUg+
CVKoDnV2W2Wsqlr/K3ZKN2zeqeq05je28Z1LiTLUldVYrWNtN6xN6oJrS1lHKwopfElQzxx10DNb
eIAi4yoxnNcNNCZtJbwl2j9cG3jOBlZBxoHNYE7jXX73YsezjYXfMcgomUETppqxR/FLGmA8X6yj
JbrLf9OIiHg8dQZ5F5jQdfWxTYVu1OqjKmIdHA3SL5g3rjtmIrgRhHX+3GEjUL/HM7WXysGu3xSR
m9weWmw6O9XDEbmDpAw87HCr05VMrKXzsoj40GLF93wUOAgwYjIr+VIzpxsI+fYJZsVbMEt5oARZ
3NfYtFmpor16yYSaUIGAFMPHDpF9sdu4GuO20301QSYBLW0jY8T1AM2HP329Q/QvGGlM5cmZBX15
Ba2O91fStAreANZJoOoC93vYGZNZMfxKNbxIUye6h25sNq0xYuLTSfol0gg26rj/SHNddvIVaWbP
lASoNv8TXmKJzvoUSo6iEQKt7OjBL35GB8Cx+FRPKHfzPEbcjwDgtGf9BllQK10ERTMNUpFwDA1j
szEZpd9HsiXeTHQVgpxuGHoK6fcX0hTwO/7GinbOfBuF2oO/d2sg41gGiOzmnEVthOm/HIINVMe/
5+vZzh2jv6MLd4A24TVibV4+CMio1q7tpuv/pgB0Xfd03LlZme7BC/ppNQ7QzglrDIKW1FKEec6e
BvAJ4N/rRmxJ/ZLL7Z75QwIxLDyjrxBNREEXVhTbihPFOfkDRDjJ/ByatC5OY0nP1NAvXsHl9UeU
vecPXV3lzr8i+f8UI2oTpFEpr0qSyEPXs9S7Zx4AEKTXxk4oaRsnQzFMYTHu8+yyiADREkhnLgic
5XgMElHpvZRjynh5MSqQiLt7UUjJPeDYvwkFr+DzXrc0P1JG2nXveR6Pt3e5E2NbcjrT+LoSRGNr
bPqfe4zoTZcEjCzMkx2UkdXy8oEzowWkybIxrlrWBGrS9Jr9cw3DFU5rRR7j9XCwY+E8HKjasKMX
UdF+FJLAHSVNPY6o129bOoyyKaeeZaj9HyW1f2MFmk3lWTYAo/qlOh4A5l4FsdNZ5g/JLzK+pZby
pwLKI4gMfXArwpwzAMp6GP+eZKcefA/Vp5rp7K9D2uIuZ4bVPJlxqfc6NATw5wDVg3TpzBd+Isg0
hFLU1CtblOSzOSB9XktUEsYXEGuvqwpC50ZVJm6zLdnXHk0QWIIqMxnj6OdSlxsdHaY7naVQWHUe
IlnuLNdpjc/aieLwnNtoDqHXpcanG4bpn90h7vQhqa14fb0O+c1DOFBaEszxHAlpKxmKOXNhPw0M
SeH5PAUh03PDpeuPleJ2mMLcnGGZSSJPWGGW8QvyOTU87DMycpfV6ukqWivU8HNxlvar6z2EuN62
2GxEBkGSYG3nuzdn7LaQQln8eOfeKyulGqf7yqrxElFF5HI4vdG+nZ7loJBNa9lkH59KqbfTeW6G
qme402Ko47WE5Vg+t2lD/TRG6VyyjugJyHQ28CR8CFK0kaKFs7PPqIVFPsN1tf4LkucEWXZ3kbOI
ZCaygS8O7oIsTwHvZpABUj3tgRV5A+oo4y39ZX+1zHzNDHkbcgiWHa5bk7WVCY+Kv49CdTzpbrVS
vBlg5EAU7Iz3Ln1N+DST53tuY35mLPz+wxDhc0/xRkmiWRvk9Y8PzoP79IcEtIr/mgE6oD4B4iwM
weCwOu2Q8ppM4UxntFXF/oJRCHikTU69f8EvYNExCXi3zzxpsp3ZG/deq9jiKgqM3oADxwwtw3W7
opeRhq1XECfLLM/0KgAC7XR/yrkyz9vJpqf6R+ZhL6aPbsraoEdbjMTAnUGrIvt6c9FmwSFzYS6o
+OdCWbtLzoRPxcAal24a5rCGyiZSm0cMfPwQEt93oIr8b/FD0BiXf+ezh6AJKX8seYpXwZhjZB4n
jugoFLgMiE9PSmkvDBaWocYG2YYzgWOZIv5d752HsKUiIiotZaR64rAygjYDOdf8Iy+CKCFJtfUH
KZgB6ZM2kW7hyXQT5ESLxM/j/MXFgo9fNxo8ZFVQQeDC0etcFt4tI1D1329CYNlRDwfsT2BztaX2
9V62ta3C5USURXcGxOHiY2jwth0+IcOhFkX5FOZWl1LM0/p8jiVoELQ4ddftDdS/oSuUhxBjeuwG
aUvsfeSETD8Gn9LkPDgV/0Sn3U7/gImjOyizEKo6SnQKRvH1+39Flt/+3RTFb/QXuBDe2IhYbouH
MT0hjIp/8BB67zTPNfx02TLNzwcbIXz/XxpNQimbPbesvKo78+J6sTj6ZCWQgXEFi13S+KjNGpBW
YdiGmkf+J3ItiCV62ULPpiSWnrslFnyt64KMHt+gpWOhl9kKv5LuaQnM6lLZ+lrHsFGLG1UbmDK0
dvWdYYQjb9J3wMmh9edkD/YNLfg8T6BVW8ImVfcPd2oeu6F6ONC21fyhSAcJ2tzZxhOXVtxoQQLo
eZDQkoJvH3x0KT0mFwkUhdEYWF7haWvfviaIC+r1fGyf2u22VC0FLSqOtdg/6LQBwu4NZw7ZAlJL
gX4zIdvIc1T2w8Wre2R/TNTmz7sfJSw0V4tHzHI2y7GjKCwi4+RopihbxQEwEAN1WaHaYpSPrj8T
hS//V2LVidvRxQEFw11piRa5R3nmBo0ZHojF3BgroQeZFtQj5IpYxYUPCqIS0E/ufyrqRnQT7+FV
+5qXycYo5/BaRh2ZNgNv1mU0hC1DPc9mYX0XLG8ARHYOJFtlRq4zgBpjqaOYzFAxtWIu7BYx4DO1
aHPbL8mQM4YE2d/8f9RihYLMGQHmMNl92T9gDG64oee2BCm8RLQdFYQh78YzLxziD4jSaouSpQDI
gwMlSSXoipr79ReH2i/2fxetgbNABljl5Mwc17yjFzphRNIBVa2BdR2gBooZcG+0UzxZ6/x3059B
y+n1JhZY+bNg2zItcxjvH7eZ/eTB52r85cHGLsNaxoW8L5MgmLfnZtObUEFApkGbIcLZU0lrTgHu
/buS0oPXdx7NpxdigX3wsY43OQR5t+5s+COfG2IaknC9X6QiThsuVV8owTp+3Beq8FxKfUUIc3Lz
Cyec23K+8XFfTDVF8/kQ2YcUqD83uoCOzPvFxtyERlkrBN7CG8JaATGf79Pi5j9qssDgsB59CPJ0
n7d5hSjUrJkmDpaxSoEnSFYi1JLC0eJb5dL586fjniJGyE0G7NzJ3Wvyt/524u4cDS3NoqIPWx0J
pKW9Rl5b9izhVLpItDWKIrIVd5ZikHV78qsakaPMc3zykrq8HWVOPZkUYzEwulGM58gcgDvujCKN
LnLkyIisazrA3qFNAnZ7ghXV+4s4UAd6O9L3G+L5DVE2SH5ML0djavnbD8Hbxm9mfwgtnJMYo51x
+i7T6DX5DIV98J3ro9f+6V/h88e1KH+p0+cIt9yLrxTw32XXJnTNakMoNfdJfbuo1Rfsf37dTAcP
j74a8+2lbFIuIKMHdO7Cm8TSGL9HNAvhxcOyjc74ytl8FB558c7l/D+LQAbDBrZb+Go8ihX1nQY2
s/ZcE8e5iS3kW0QZPnWFfJCmRtt2NCuiNhEjSe2lKQr9uvg64RVRmlFCzs3+UDjJELSj5TUtkJil
UCP8ajtR6MpWaghsfLIEcxJfghruce1uoytffOLbshzKFxM1g9QFHoWIrWGQD5yvKQUHSbILrP15
lFMKuFu+Gj+kGvKOjU3G2UsoYaV7dW3bLo5JSOlBcUC4pKom96zPPOx0K69UiOfoxRIS6edwZxxs
NV1YeWJtO8vNR+9X1b1WB2Pil5zkS9zHmG92FzddTxdpSAlM2XozhFSZdI1hmHnwdSY4pgQTGHMY
BBSP0nL5uxshZG9XSpNDORQWC2X13MF/oDavT2XvidDIvQShvSZg6TIhHBCNJldts0VFYmoJFnBH
QxSbwtZDCDZat9jgRnA1XXh5Pe61TIO/7OZce8RMAhgs51/n7LuUdJFw2j1idMwGgID30zqKAkww
OKSABcaLKX5OjcqhCcl9t23irefxNNRKrPPnL4SJhTKvRylXxGpBovvfKQF+EqvR8HMdNJtyqx6M
rSPTZK7w9TE57YOIfHD2va5w1EA2XHLmVV0uF95tPCA9cVM6sDdDwxvx03zNqvN4v13iSE++NoVM
K13b+S94NCIKSFGbYw/GW+GlsSLG0NPL/hDRHJih4QyqnQ1Mf+fF7eRPlS7V49rdNgWFymZ7c2vo
fvPr69zazjay1QdZ0uUVcj/nthI4FKfQJYhjGAWhGOQDkkp+Mp21wvb/cq4WVvyX10dEBYmtNupk
qcPDJ66paoXM4QKM7sPl05PzZpJbSWsMtK6zLrg5olWDNhYQL0gvetl4FByNmA7AbNSDnSSUPAL6
UF/OFRDA0XUhK05hONiFmMtLGa8Ux1RN59NRFmAMkWN0SEVYFHnFo/s9fh+EM/UpJ+xrOfZmZIIp
aH4WMKOOnD5lHYEZBTkqpydlMzbJgJWUViBJyGl+N25Qqf3wLQpaCo2nUid5n566iPYuvEq6XdDg
krlDR1/eKjb4whrxdEBKVbCCnRyFNYZ8+12/XSu5TypiEhBn/aLhl6LBJ61Fz9SuELS2J5d/uglD
E2y+FWg6BSd1YMcjgv7p9hBRi23ci5IWLUlnZZWOQSDBVEk/y/jCZBzLPpO8gFk/4GaFPTjvD5ie
T7ZtNw3k2rWqsf6aXz5p0jU5hw72RGzVm0Y1UK8eFVS4toApkFbCm0UZRCnHjWvoov/dTpab23rM
f0JUrt4jhzKJ1j/bfNUwDcdJkF1KmV2b1Bq6dJlGLdOMusPJBGLBAGcyYKRCARqMC/gJaRIA89Wq
oC4qJMQ7t+7QQ8leDEa8F1Tjy9a7NAO8TTpdf26Zfu2yDPFlc+0emctsFXB1OVqK9sAI3JApIW85
hin1LmYEgZ2xdIYsREECTMik2QXUXNALclCkDd418I3kbz4/ko5KnTI0k6aEP68jxbyadesFWSDy
f/o54KsSQ/5T25ORsyoGArYLoM04szOLkW7cOOmaxiTMF13wz3LwWitJJOMCxc5+Z2WdFb4PU44q
QkpfLstchXLurCcrcLnosCpwNQ3N7wfLthV2QA1IinChAPygNsLnfIRUxrKidkd4PpChChg98kWE
cHoU8gU8p+ypTraT7AFQxIeCL+lcq04vn1C/UbOlnML01aPaSX8ldAPwJbunTnhsm5ZNuiwR/Z97
2LRLdH8lAqGEK+/zSoYt5SdOS435H6isrQc8050mn+b34tcyf2iWedbVSE88vr7OrUKDBw4WUiiw
BARa4T3sqaOz0MyqPaXu3gGCeOM6w3TmbxsSRRGDjy1aK45Pfd0Z016Wd9mdqWeIdy+dZQrY8NPz
tN6UFS6EFpj5EAq3fMs9ha7V8Zbn4E7rqVhDLMmgUZfm4RybapR5G7raaj2+5RJzcIQOlEzbETMv
ZX92IKr3Rpixjn4GfH4OXbi7gwBSUTvr6uzUpVE0XHA/H8KmcBnw5woM8B3vlavregjj3fCNcVht
+co5hmLVfupT3JRmykIgJODmuD3CAFgR+sC8SRHuRRSvlgop/N07ozaa9L1gATdXJEGIvDlQpy/z
Prq9tEZtcGg31zhaS5FuDj2fHe0oo2U9tqden4hIQfxVjFTsy5uRWedOEg80mPFReicp53QqVPnG
1TufEwdQ9+noNm4NgK4mpSvbnd4xT6dZ8/Un/ahMHw1FhzZGr8H4ifROkPRft2UeWK7HkcxS/LP7
2y1kSPaHWWpksAffzyqbr5Bzs4kYwwQ09FwrK0622I2V6Gf3rIgTf/s666hCRp66pa5XachH/jsI
WwvGVC7XWiuDJDy5pnFbespSgQeCYpHAlyYfJkA2sNAsY4gx6lOQAyOrjC2JrMN0qFtYhbRouDEm
ZJGLW+e/SqcbCg6PGQqRgyB+knOmxIqufJHc8s0tzsetGF9Fcf+C0AxrExr3jdVadBRpbDknDfTc
KoaEmNrbeZW83qIOpSCKZi5RxIjMV4IK4vOqD8fEhXe0pCko8ELkL1biNEfz3M5qshrfLEB5OTBc
2lsy6diOWJm7Q/iPOK7gFfCQl3+SaS554cBbumqTSi0QzlKeGehA2trJEl/0W+mp6XFzTvG6ih7e
X9HArEMeedbkL3wr/ppMpsVhdStxUyTVZ4stS0CSggbYzzXX/anLkbJmLqdfw5KdIm80o/dZlO56
dvTTOMEQkYPgvXeGhfI67TH9pSqZL0ooGvtPkWHrjot3fdziU+Cl7r8CyEXP3AU1zznotXdhJ0nB
EjGBmy9Ma50cWQkAno5+qT/UW5vnGtuEPukkvMm6IC0dOZP5hRwiAUHAkVg9ntPF5hi7ZiWEnswz
XHyetR0bD7Wip3dOuR4JDDIal03L6vNe5rZH9fLot2JH2IJ0n9nftG5QjIrCelfi0zRhBF0DjpnU
HY7P/jWQN6cg4EVLWOTduFEtsuPlzJGAcQYHD+RhZW852FV/tRbRsYE6LRKACtSarGeSKwIfS3hG
owbTDt+Au6O2bB5kYuDPOA1fIzN5R/hWUksttiwFUrusxkYzLmtz9VVEiWqHJs6BXliTAVA2B3G9
lkJYEsXyaDnGsO2lwRSslbhW7D8SwQxQMFvHXN1tzINHDbCVeQb+CKWsMcnolfK6prpFa03lfevh
soWpKFQ332ECriO3/XIgcMlFfdqhHh/p5pnLzP86YozFWgMk+/Qwkh/Me2NeTveUK6xhge5VTqok
oy3t1R6oudTzjBhZp00dMi5OtumZBFHBFOpHq32JYdWW/e9TPfc+N26nLcRbd4wvTMtm5H9w7q2W
u1t0MglHOx1iV7kWq0Gy5kEOjK345diLNxfKSEB8X4dKp2YSz+nOpmrOLucRCsOidoBtSs+6dHnZ
klVNdLwWwDfFbFL8IhokvDowho5zPG2UbhFOxgD9sG554Qd2Drb9Mk7q2GmwmD+56zQ8YRbSUMH3
UYEv3euQwAG5pLLW5EKAagyIbBNZPPqFT0vVc1EkF4ohlp+JMDfZGAhtT2ws+wERgEDzdaMhk/fN
c3wziCiKw4ZzO48gcsRx88rPvrU+K7kRCmLBv4thdDP+i+SYZJ2RVANhgOLhvbmdifWcpoHsROQQ
DIvyPKri2xY6imi/tLJBoi8SjZ24NxNfJ2+5u/XlHLLkrsqRCn2P+RuIQkPf6U7UAWa796tmkhB0
zT16MhhgB3y0svegmBc7JP79Cy4ySTP0LL/YleFJK4hYBUEqEQhRnqkE0By36DAa5o6gWJ74JnEh
7onf4ez+/JZvj3tv3/FOzjoaf3Y2MGo7GcsrO+TAMWoJ4CiDFUMZqGFw9M58XQsja+qneOGfxrqF
c8eCwO9CvioVmNC0xjfKDT2FDZepQia+Ki7byRCT8V56y7/G5PBk9BaGQP6JtM85cZqfl9EUYC9X
M9NmZPwjtq0D5JSUHGLI59xi2znxSVtFrl7dMqm06EIK9dtJmOCxrUhBFjrXeINlzqeAzyH4Nf6q
lLGtbIrLH8MLpDdwdFUFqT/hZxCORDko/NkD8XrmzpsntxoU+a6No2fGoYFxtsE4188m1sQoUa4W
Wr7wnsC6oTFJuhpIlcmR55L8HDAGFRn5XBMWhf0vqYEU0jCgoX0oLyV6HKDptRktvXu+fCerTCIm
YX3S0kmewhiMD7LSBpj7CRJ2rU8ltOLFOTCaoXQFFz63wiK0kRYXD5xNCPAWodc0Tx8LPnqiQC82
GXZJiPh4RhOaooMncLnVqdmm4hYkcJrInbgjPVhJoVB8R5xZWnsiMFSXgfZWOMdtvDjDd2O0o3g3
tBH5po+95Z1RorrbGjKvEpGma/dUf6uCMtCZrEOsJcQATA3NgrW0VsiQpMLbs8JUwp+rlA0PkGd1
uZq3nE4/ES1Na7gc+LyJMapyb5J61dD11s5looRKY2MfkynZ+ODyhjrYHrOvnF+YcLKBit08Fg29
0zJIYtp8WgtKOxBa0hhk+jGnRwKu7upFbcqyuJxz3zpFrSMDBdGlFds95naUVD9iYLsZEmizMV/e
9JLXch/U5S7+lv4wgIOhBNHp27+0hTsQczz9s0Cf+wczEO1eGe0Ut+850XLZe9sWR6unoWuAHILB
Lbfon39hujLuuWdCv28orvvpe3oPPDmjxINjXpLWwEnAtNnuHUZnS3MT3kQfnYRO5dKe35a0jYoa
T65fcilLGRUNcHeObvMU14Q0p7Bn7e1Pqsvk5ayPIRQvy2gyD49lfIg/W+PZDyIwEy2wpMB7hy37
Pdvl4gcxwU25/+eJWMDkI0ypVZev/mSqh1+f9HuBVptERe/gzApOwysgIf9IhvCXxuLgUqqwoubw
8haQfGUHlUsylqhMFiaXwT2N51pRJLUOJTJweDocSKhXE8ebLa+nv0HCh8fRv4uiEfl9bXqf+F1Z
vGEr6TAV3EEU/7jtBYOoUOZDUK31pUz4zhbeA8lpEXnXylUqQUMD4L33JlOqWbc0X3SK+4yuzlXX
wcxXR+J7Ct3KRfo5yPO7IpNIIHMrmtePEkR6Hcrzo0/dgaxhYgjceWK4PoSxYFsAwScp76+FbDqN
mUqi6dm7Cwd8pLbK/BRXC9kIqlpZzRD34bKfiNxGH1zKYuzEB5iil8PpPVH1Qmhpdiv1Tfv270M/
zpjKEwOrqbGe2wQXbnGqrTMQMFkixc9R8S2lFzgb//O+IBpfLWBppJr/gkRv2SteM37EKVcIgqKc
Kv+AxsfHDUzgW1D9RTEm1Tv0/Wbka5O7UtGNp2O4riTwbOF+VOSF3s3OADzmvBzpPIbUD4ZNxwAX
RMwJ408ISkCJczPmGs+f8lI/y8N/AZQRm/ei32Ehg4GRAM1rX78iQPLl1G0AZ/CZiXV9AW4JtWGz
QJpRmMl1kSnl+TxecUS4N+m9qQXX/08Fcj1Q0LACMMzSNnMoowGZ5xSeCIEzuFVLOCbNI6KjlvvV
iuaahcaMo1Y6zRhBImDokzmEUlNxvAFLn3rbG4uuqgCwjZHYI1FHx9lWalx6p/YYB3BP5ladSEyr
NVj+NKY+ED4sLK8G/EUU6siBWckKUXY1hr85K6ydtWvm3lcyR0QOifJwsVkqSujZLbujQqYOYYlw
1IAtCtCNI4gNW/4+LFKYVF+SK+PPNVTESDSc+cjG82HvrLt7cX6Tzg5xzurEs8s5Jj5cN6GAyBZS
REaX6MBqAdU5pa4Z73ce0nsMmSwvF53ZAexsQJ2MvN1SrnW3mmcY92RRQ91Q0JAFDxd9aV5d+zKR
/jKmu/veTORIQJVqKsFuYsDq3bsmCnjTlyhspuEKgcb7UVdqFbFiTwIuSQLjbcLHn3/B761hemJO
SF/9gVXEgrvonoiqyva+aCxneQ/rGJTrDLQV381X69jAjKgb3WGPcej78dlK5YHT61jYq05y1S0/
eDxssy4+NYNgDgtQYWFBlIMTJMGc2URK3peoxjUP66B9yDiGIuYs9PQQ5pcGCmEJ5PjGRhCTF2mN
gw4v10gBvCWSfPO5yrn01+x2SWx0f57g3TdhYDsUZue9RJ2ySY3zWKPvTlmlwWaCzFQAwHmjPJTD
aRHU+AsGwK/nnr9avQMH0Dq/uKCQn01GH0ivqzVerZQQEDWNW4Ec0B0vAHCppmOhd8cUE7+KncbL
A2h5O+i9ILEf63aI8Ulxe1s532vcUHIVllZeMZjROFGx50Wdq6bNNatpfenMPzPO2yovtKqFPLsz
xqgr7SGGCz4rT2qeMpmbM5tXBu0sN6G9AGdt9PqUleFzsucscV7PKWp4CGjqvgppfTzCSLJT+Epp
rt4P1lhJj00bC9R7p/8oYmVLOEuMoFQsxt/lNFUrpNKPDFWRjGmLnIVxasW8O2NOBbakzk6RsIZF
0DMso0Yh0/0Wcf6mD0hsjYBZjXH7ZaGUWdY626AgKvb5Oud9ViphVG9L8CvMst1ya1mzgN/3czc/
NB059Oi83WhydFC7w9XXYLbS+TOo31W4ZSWmB8nF1hcytjFmKufRc140HUKE/n6oLutGtV6sQ1iS
tc9wL8Eb2jPabmtU4UHM/6B8xUd9R9pQBhLCRlPS3Xnz94uQheBN1WsyfM66AVIy4ankisjOEmZv
ObhcDN6WeDridPEvYAYm6mfzPwlTmnf1nReWbCUI1rAkzs1Z23mp2NFRi3l18uEPIOIrcUJIS5Lp
W9XTwqJZ1mo3O5Ehi9INvXpAFS6oHyE1Kq1/hd+jdh5rT8qA/oAXArftW2AQYTvPlcLgbK1nDc/J
p9r7mT20XGe0skYBQYCrbT0RGIV35bkCYfg/eVjE+ImtqRcZNOfJUfpN+/Ml4lcxdbuMc4SFgFGJ
0rYj1vzol6WEGaZtLQR1uQ4uefnz7lK6MVV4LrwAzXmxSbxteTgnlfjZrk+dOISgE6Qnsi0srgEw
pjLXmlXE+E/oOwcgUxhYRYBUrlIBAimlszoTimLEMYFHJBGQKa9cSm3brQCiTBKM0w4Fi9QeK4q1
3PeMSqK5Tob18XiA+ge0dy/m6iwQ9aovX8azpBBPlXnfBt67ToSlONuaN9RULFp5nix7m1HhYLwG
nnfQ/yi60rbAgOpC1Z/MX7ZIUGQnl4X2reHUyWdrgBjpb9oeK+9q564bVjsNS9vgjVuTUK9K3W0V
sgu7T39MYgPLFnSyUPf8huPdti+Un5S7rdPBJ97DTCH9wuW+RFsK/q017uK2VfmCBp8iC/mNh7Rl
f8DSoaL8R9yzuIIOWSypra95ARnPRdvy9/jl2CD/T7Ftj4bVTbASpNCv7PZ9tMZeqAfWNAQVjY1O
oOrrE7tBROVSN7FqDiuRtcoXqhKflRY2hazEfpvQC/6IiDD1Wcfjx1CiYpfCSMX9FpDSfH09gbfj
biZ58cqrm/d7rzgOIvMWeNsKPHYkHGKX5rMmb32jyMgNdqC6H/D4t+UErOjtyf2KE1VWAng5Xw6o
Wtv3GJ4tKHOL/CI1N+k4lkJnRPv2qWHQhzFRUx0prxWEn9Kti8dLyddhLlfyc4uwNR1wv5W+IYSu
GrM/embVLHIIaN1C5HQb2G+d3QVTyA7i5H5NrLu0o8emakmw4ThOhKD0uQcIxa7c9IaBZs2x39nI
Ezq/Nw7WRi5co7x1HZs9fYVjBvIU5NPOIn045rLt/4ZFyD/XWkPrIQtbSNT/47oo+cnCST26UcRa
Vz2gX5S9fvOF6p9clBCIwp5iKFLErp8hKJ3zQc06ecyoPG4E5eVuRmjXL+3N9EhbEkwi2FPkBauH
Xqg26Pef/L11SaS9EmAcvOM9PS7D2i77Q/MTRt1ak7PWH1cgCiINAnA49gXD870qfIo9PwWlCblh
Ou3k8Ob+tFjDD/ZTUrqjpbOg6rhhE8EEW+WuMa0PFQ2O7x50lXCHHfBKmBU6dBw+s+TTKV/odGxr
raEUms1/3SuIq8hmGf0qmPwWuAeU5OKPIQsADGsJvQLLmh9tzM72ZfnE3UW1oxFe91DB5C17QHW3
kN34TV+83bwTPer8eLv9z/xz3ThKCdivdeO3fL0GVzjzKlt4b9XwGWk4dUzV71Hp6xsK7xyYqOj5
61IDdUC8PGcfOU8EFzmupEY2YHVhToA9GSWs3LXhaWDgybdHXMO8E+076guVVqM6N7E51xNlWAwX
LRIeF+tYmwwKB9t9L1BUf3RaMyEKUBSYkbk5tdc67ZLTj/Sr3aABUJ8+3EVDb/fgJKdIxO+WVykp
w0G4PBCCFyvI3uEGm1GhtRKtcLpQewGeA5rYJ/gqvzkZoNI6K8/+Xx6aNWREOJFAjGXdohwbF//n
DmAConlY8qFj+a+K9y13mlf1zdnagHp2ZKN6GwVfBcYvzQL1iwn4kprL+D3uY5+KxGbDWovsa2f7
d9QhnJt2LgkDyIODyu6AVJn+se/0X7UOyD+AKuEk1Zh7uXhwMkfUB9WykBWpTWx7na72QTrJGJMX
Cd6j+cFykV3GnttwAMPqinY7njrSge+vsIc/WMPILJ9nTenHsrp6s8JT/DUJujFLsQT8Dzz9ZCQU
6DNuxDj3WBewMIZl7s2BM/d+iQR8j+umLMUiUWlVGJVqeaBHjVGCbhiiO7cCA0BFHk1juHfKtKd9
2xOhGqAjNsiA/RG5Ybanph80lhlBY/riUx6jqHrxgdAGAqMJ8O3t7qIPwto+ID8tJnZFWT/5B8xF
LT7+uh9Lhzn8nuX6lQi/hs0dHgWeoGIYRHbLxEcb6ZZoyVTrn0aFI/9FaF8U+J0AIZAxoJfYKsnA
n13Ls5zo5CO5WB6IqFWUzZXtRZcck7pGFsJKMWZnzsP2xgyLJCCxcqkW03/RAIpkhl/IQPVqyfON
x6Can1nlmw04UQW7BnmDY5b0VOP34NYwPf1eEp10yjE1jTd6XGkE9pnDTLmzhS45x5xSbSoVkKqB
9GzosEIg/zU5IManRnN7FITig+fToz4Uf08N7g2JC61I0UyFT8WUtQd/fYehom5oqtYrce5hLvqu
Y2GPl3xcAVE6oYCywlhNNhOVyKCMNe6EEd2DVr6uFRXkQUSIIZu88OXgj9g7P7lYee3J2nmqeRCK
tbE10rRMNGmhPFQJo5n8tZidUTEhHfCm2saEwLF1ugL9JxdnDBqdYy1zlneNPYqRgAXeZweOJP1S
QerQnS0tU4ZwNn8lSZIvyiuTUuD4xZ6/WpY4koJSakO7Rzdo8Qa+sWMLxmTmskz/gjqXM1z/V5RY
jWuUd0fl0YG8tHeIS1mbt0lbZbRHjfDRGZ2l9i9cOLKGUkh3U3FsPapmGytAf0sKVYXin7Yq3Wsx
5LuQCa+2Uhs7j+6Reg7aWZSoei7PXG3KQSezKgs4GZ3zUJSL0roYAXlRlDNz1lIGjlhRHV1lKsF/
dxLfzWO9N+rGSSFPcATPMAIFS5rFbw7Be8G7Wg0OCzMSpiqC7T0cyCAPdlmqFslFCa2ccjrW2G2o
5njYLmKy9nBOhyLGvEEf0TpXidnWIj1qL9STaGXzsUcLPaIYrB7uUzcwEu4JkNQruy9ZIDnRUGA/
rTzGuXQ4XE/FpEHDfX48LcmASANiQHZxNlI8jppivAeyFdWtUmZV0sKuJmnC2aAdTE+SHminkeGM
9Ku0aC7EgM08sGgdREfNz5pflpeLCJTY4xxx9Ct9Y6DDIG4XOFZbJfbHAHyiQFTR2wm6jdKrONyu
ui3rbQmCC8QqFLzdduhAmFEARtUl9XxaO75LcfwzZnN7XKLiOHctp26e7dvzANm/+XL0AzvU+PZS
P66nuy5n04HAvoDT3NIeAWNTSL3CkaLf+0j1fay51LBHHL5R/kM6KtXNlXe4UJVGfgLz2VTrD/L6
pve7oATXUfO4J1POeUzLbivd3iXgyc6qGCZUIrazhuKG/le88yvHV6gFcCWj7qGFHEI8HzvSIK3Z
9EosNxM5OajMKHm9nj7dAlUXbmqoAsOQHVdqLXPI8THrbsOdzV85L0xtTiaRWGmgCR5G5Nn15G+k
G9EX4SHytd/hMxPObklcYTu9nZ+X+KZAwqaANGyS7BS75maLSL6aiBP7jVL+qQFrgb/D/O1gkpnv
nX1Pu0jrwE2YpbH9+HAP8w/seOSX1hWGxonxK2rxwant1HSVTuM+nvTqxf0g3X1SDaD5tvD8Oy5B
M/htQHD7lCVm2FrAbSnmr6vQyFN1i5NAZs+XkufzHDoBXKBIslojbObMOiv894Pw7XBNWhkaVSD1
9rhtWRGZNhxUADLG8DipNBroVIu4ILJ5jRdwQ4YsF2uvJ4WTA2tHrR3+ONe0N1EswDF6Zod08MYv
IuuBrw14oiyoGtxmoQzAPkzAEVOO1h6LWjFFkAtIZf9xjULq2n6USHxdJaYy6Nv6Yv2PP/Ri+zm1
k+SCHHnc6BV+u85MZn6vcja9NGHR7thnlxPsaKYI2I46d34xXNwgpzk4kVOyWLugjxjWNul6nnKO
3taVD0m5l2az/c8GjK9GNSiDNCNz2TWYfHnJEw4h7lvjuSXkC2cv2T/J9RxQlg0aAI1pNwkEZn47
s1bW7DwEzCjMI4UPlrpdGWwE6aYwoJPdJmFwkgvjkX0G5+3yiiVJ7Ru1eOdEi8v6G5mygqScfvM3
StGMii5I4pEyikDNE+pTYbOIYQKRxhBvw72up4Hriky/CIUy3jANRJ+oE++RgYB45pJfz4cNbkTD
SoJnLWZ4iDb89w7KGpvbJATKyrjwuic95u23ub7fw4iIMsABqAlYDFYgKpGqIOcwwPCli5S/dA4W
IYMDyhWRLO5Tjc7fe+3J6r/Fnb9mEa7Hnf3LDaosyadLYSNIWNOU3IVAVoXyrCYBLpVH025TTWUd
ePmJxZvYsAk6NFnvuXmOqFn3A98oP/jlTRQISFBKqLz3RUAP6qg9vSgv+0Wk6QHAYX70vYtk5wGX
9ojvWj9VTkKO1F/2dnX3k6IIEg55CUZVkqUvs3V7XnnBvO2KcaAQ5BOl0il5c+jiB0ePHGvciAff
yDRIUCxtNSEQPkGYr9u7W89LoruM8fAnAXMsV5zCoCHjaSXaKwngLC9eMc2BI0f8WB79wj9e/ftb
Gw/+714lDVhnZuMDtiXgSHZohHH7gbpcxUPAJ9cbiOF1QRKAjjsJVqas0/1wT1OERRQ7/RorslvO
pwCkP9sBOlcGi6y7/4TrJelSnxNp+Oj2ZwtwzYcYZFUSsRFu5djiMLujLyrm5P2Ic9+/zgsNtOcg
975IRQPX8llsv5+G5XR9Brgqk+p8+bDwdgVhTsElNdQDk0lBCOyeDCq0YKDPuEnKsRUHh4QdeM5e
KqIMj+oZlISfAt9LADXhJ0GCQGOMiyJAfjqObihPBnpCxmpYRrTHP2vTAU9A3kL6mdO4BKaq1u2b
+GIykAB0/BT4uhA9H1LbRFhj/SJhcvDsFXHQTkFv0e3UbQlXToXVSy5F2iOAqyAqlAa8RLGBGq/O
RHawWWYf/D3spYEIfPc0OcNAxZoQVjjYyMgM4QKZ9FRrhenvccKGDL4+Cy/9SAE7Q0TEFHrbB/Qn
grLEvEp3h4G4Eg46GtQTeBKxUPA3ln+ovQbfg+mMTHkkdScY9UALzPKzjevlPtlbLQbDq57q4fMD
aSa8cJGuvOTCR8hurhOIhdM0LQfa1xX9xEQqWQY9SNlcrozPOJxi51hhhQhX5RKt8LlA7QlMyDF7
Fdg5JGlmkZopadWuWZRbS/Z5UK7/oduOEcgfTdZUGt4yk4WlrnqODiQqo8MwdWXtz+vQWECr02xX
q6kKalmsWVk4S7v/i6z9xFakMzzfVUW9UjEj7SYI07/aU9TNBy4Z9ug6OR2mXWDgeDc4QZXX+jB9
ZHtUssYz1EvC2ukIAclqdOFS8weS6K03W6TN5z14LAbZmEMYJ08GRcNV9sTwW2a+ypspGkkO34qA
dC76ypxOJZ6ZxQKlCmtuoi08ALUW0srYqZ9nshMyaJgi6sJ6LLaiGZSUAZmmR9YYJ42YCXYJwrBl
CW2fbeDFFNDOxaFjyqUbB9LhOHBEVVDCCQrDn4K334G/vDSnR6Yf0KWn2oPr8tW8+4gwN1MIxHys
yBrwZoJ/tmRVfx0tkDV9jBHNSrm1vgV1wIvErZxVRmigult0mToYlznxqG3+cbpCBpoaR7r2B4ut
WuL0adafMav8B2/ue5y4/LoxbIHrqV678ZcdEfMm3iKwlWc4/7bX6WowVdSWhWCcfVT6C+jnBf4J
itf8hoM8b91UjZoIW74FRuvjCUVAfQrhNxpPCiKUioShUB+sBrMPhwKKvamcowa6RnjLEQRgJ5l3
2/ETOpSG9Asp9NvvS4F9rjf5sH3IPpDI0aVxEKUVN5gobhntCYNcXqozcdwOU7fFyn15wkofZkv7
QeYjMLog3uqaaYsPyO29XJf2sWM/XG//xZUNiLI68zMEG4aRK6ZQNilZeSLrJpxVkNiF7V6B6BLN
RuvYklrpvta+sH6fqOiN95x/6P8eNcS7rQ6DhY47oEXObbPbSJxduXdMcDphqSyWBdtNLZOn8f51
PLL9UvvH8gkEvZxPHwfBG+gzY3GrJuEbdrle0Hgb8PpqfYLCBQI77JklyDCKF/PYP6PC2AWyuDUr
4+ee68IoiJBu0PIt204nMXxOfO0nDawrbf4ZPWL1yLQ71oJGOSzn3VaDejt0alXKHPDojsHQyGfL
HMwcgPBmZ+bp1vUQIcTn17x2wtnhU2YjPW0nL55I2xUiDvX8RtMhrxA4h+Y4EAxUo5/uoODwgbZq
3zzlr7FPi6cLr7Md8Ld8NoPT8ue6hGCrgLO6w6K3mV+fzl6BEuyVxGDsjOzYEoC1+ToKILQK8CYA
A6UWJH0GTiPs/muiwAAXMBiFLQigsbhqy3QyJPgDUoR31hcTHRxBcc0S1c9r9J9E+BDJaMhgVQVO
Gv/3oQtVYg5NJ3KmtX7qSx4F3fjDZdI/9qVRCSlXnnPKxmOaY7lIMSnXF5ooTDILvt9MkoYTZ3Jg
9L//uULgdQOLOoOaPunpPl6eV25ext0bnZdoiKQM1SZlKyUu/JjctCZ1t7dX/f7+SW/TdHEaKYnX
atAg6BeomqafGQq08QmOu6mgNab9lyFsRYk5osLHkJLwa9DBZEFTtho1sCmTqAe620t42bpr6jGj
s9+r7m6L5LITeaLtVmg7kvmrNUiEbp0/xzEjQNKqNSweZG6cWv4iQI/Uunp0qgrWdwxdmXmvsDno
WxdTYIWHWlSBlRJ1bhmDq7vCaVd6JoJNxkWP7z8cmXhhC5DH2r7GtUX88QGaYzFiq4wdrn0WBk9j
fJpZmP1e/AKY9eYX1RRUFH2qHmOMCIyefyjRA0KFQscCFqmzr2ewS31e9kAhLxF28itB3jCkQiEr
Ptz26M+nwfL8nKw1MnjKSS2WPwDg/g1/HFwhup4+dK41OyaBdFMQs6sIHYfrfTXchLbIO77Y4s5w
YZbP3dHen28/XbfpM+Ah2yOsraf4z6vfxzrY3NUVkz4HSrkD7N5cEZwBgV+ycEKiBhfW0wJc2bKS
xVwPSVEG7ePRD2VdswVMXIVjWFOoTgh/yh+7zvkS70k5iuHfqd2YynLryUaar204m27usSuL7B9R
hVD3pymgWb+6Bf5VKsLGmLF36wdLOPxDLzsEkP0EHJfIJ+6CCD/tWTw+5SAE1izPInzNal5epUGf
otJtQnjNZududp3mI8dAAxN5x4cCI6GLGUKq3FqGKM6AWoL63zj6StOa0uGKxNu4YPhrqH5jHWCN
cUuP4b+2oHyuUqIjkGhKuj7FYPWAGAa6qzAWWBSzy7LyirUExAtjrUnRsLCHpyz98350mwtPhD2a
49dtJF6WpLOVnoUSP8WnMLvzSG2hEvCsRlJwpjXSm+2ip/4MVCsrf3SrrhulJhUjJKrG5p+cNgt+
idJhXAM8mNEzn4BiBK0gtfWlTOR28D1/lwesTBUjwB2hsevje4EIW+5WUrHphkFdQxbisPeQn9NE
MkIv6O7odOR1EAqWIAxow5DGmSq5g9cyOtSefqFSy5RkcCqgZ+a1fb9qG07MzLWOn6lacuzrPuG5
puwD5quZ+/m0C+42wxePpkAMnC660zetubwU2jb40Q/jvUpQX76EE/XbDtcET5DgIZ8XMVkA35qt
VrE4EbJlxG+5zG1XfOvGD4rS21g/NgZEnKgtEUpIldNkgFpH6LfND2huOu6BFYDaBjAbQVdAkgq9
Wo7n4H6ShlWB/FxyfVHeJxs36gF1AfpNM/4tPtUTe+paNto0/srVmoyy7vsNvmO566LzMcc3rWzr
11vGt9043ynZhjixKJCHbUzm5lD5Wfe/ax/O5VR9H74vVJwrtykLZxYNt+AK3hnRji9LByjmIDAl
mczwbhuYkIX93HuNR7ixXNx637VohS75M1sqOMQdNpe08M+7jIzQphHbm9kb539wSX4IVPG5BOJZ
pVHxDC2RCOL/VfErk/ajmZCXKBoPs9QbZXF6QI+82tC6kY/xbghEI7HVEAgC+x/SZDqezqDnkrDW
zsAflLT87Yqn/0kLSbodUU6nvVhNvzDm/Lg9uxojzNg65CP1ZDe3xhay3Jj8ncEPysHfkKhl4NrG
wQGRs7qxxCigy+2sv4t6gQSs4qX74rjTnDmUvr7N5IahxDRu65yrYJ2ZcuHJw4gMtYi8CATG5qSa
pA/EAjyLb3mJo/GXgNbbHozI6D0I7kL3L5HPU3lvhXsUzDriGr3Cv3hgH1yQq33XvrPgXAlv0XGZ
76I+tIAPqDCyEPth+sWGwYF4jd8fPuCZA82of16MvFMn/Ryu4eQvHGh/Brokh+3WO2bGFca48Ll6
YmQxt69jQZhzv26nKpUAqjOkuq0EOyXL//AglaCDJBVKvlUGL5vPgwJzi+Ii0of5pFNh6UOtIyvG
oPtETl53s51B9ptWt/7plnnncvKvoyGNSyoz7YUOZn2K4eog1hpWLG78x0euDD4GOFnfmX84jVU9
w6rp+MIVvkkr1EMPQn09M3NHwOME6j0293oK0GwrLvI8BLX9WYsKuIT+xh0AFKVsaJsrxq9LcoxK
rUEexnMQtfnVDVWVrHKRQLVA9/p6SmR3URUO8P9OdEi/B2AdzAIpzy0A9KpiJ2XjuTDRKJGHPQ2H
6wmUK4iQoDCMgNdNw1UvcSrJKcQBUEV1wHLg1bAZrjce+w7Enao2I/WlTap6zS6Q2o5R/I/9QrOg
eOwL1qVu4Ln7jVfhKwOwfObsTYNHruNtjpSTuJ+HLa/N2w3UR2PWLNc8lFKNBlTlzjPwYFUtgzBC
y3FonvZbl3cOav9NNJ4uTTtRwFpTm2uUXax3vHyYhZ8euVMaTwsv3tSNr6n072449zJkb8ov3bgC
v6w4GZvBHRSsgWNG0mPpHnbkV8Y0DMWhaeRIjI7KT6ourwyoo3D32AQ6nGuV7VXqTXKM5ghTCg+u
AbJiHD0oa7tMgK0YKTdwc7854IVJ9n35qfNd4yGTKfqqgXx0woEQnWrYrgCaxtbL/+ww/WyGV5rX
xC6po1Z7LPAvHZ8ianCq9HFSpwjP4SpRViLh3F5haT8I8zzrhjrvloUrSezekgv2LMe61eojEj+S
eMZ7ukVWAju1qL6XPKqCPc+ip6O89ROWAF0kSa/V0DsCFaOWPZUla//uJHb7fDKvUDr3lCgnwmA/
p47r2TbSjh/yA9ej6YIC2Kvh3FjRZZu8Jm554Pktvq/DkzW7v9O5d7zUMD/+vj8ZkzHtVFyCDKCp
DDzyi/Zghw7108GzbuEXJmEO3J6fQlYUaljY1o19bdUvK9F/oR60Q3x7wNYs1lJ7gtkeoVvx6DDP
wqYDTRJpLHeQPljsfryFxJ/RPT3DnYssofp+gisWI1ShWWh53S4f0OkdVP6ZswDbsyjdupAgnzGh
faS7v72nLitG2kKbItMmUFK8lPiHxTT+Teizsdgq1WUFYLgmoX7kk/7SPQD9tZbjXlepLJqQj7mu
Qe9utWmk6I8GyvYqKnma7+EbUumA9EzV4VCnxx6jkXpO9UntFEP0bVVQzgEOzSoagmkz9gDGV9L9
tEh2MeRQBpDwe9TP7CX/Vb2oR5olhBvAKKL+FqyEg5Y9hOdbSWDXm23frF4ZZqjYfRFv2n9UzNRF
IncVTcGDnlTc2/pmleJXDRReW+a3Ncfx3qzrDGZevEpimo8fLkrlRyDuC1qy7wZ0gdPMjoN+oaEU
8hKxLYayy+t8DOBOKQVbS7eMaLW9AzknptBGNT5frQDgH6bmt6+Atsgfo0TbI+cHggUvwvVI0pPJ
pH1vA6FCwAayyP6D6ue6t+SgO3EapKSeS8kw9Sdgpjco1Ptn3IoyA4gSFpGxV0GCmAGxcSm7s+77
+/YQ4mWm8wINVbT+YOFf3QVgelbnK5FtCFoZFRd+bz1+myXF7FgiVC1XULHJyzivu39oIGPhFzyf
bGx8w5xLN7IM6Zuh0PPtPKy6CgUMb8RLPCmUC7p7ywadBAvKxo0EfhyyKykxC7OHgkBXJcexKFjj
2DbRxTVbvtWFYNJwjRxs4aXozITlN67QF/0xnA+QSj3IIYGCWbN04xw4ZtsPlRMX9yAFIx4Nmbbj
nZUjn/9cJ30Sl8IO1CLU2wZ1A8A+a3HHuvxRmwN2zDWfvkyoWnWMwSu+Y8qIZsvWXafmA5zc9GWN
NjJLHM2noPpNu6QomJT1VqR2a8Qa5VKysIqpxXOsKBvdszUezYsEAsILCCPs1I0sql9wyzdGY1H7
SpTCFvhY4rvYMSvb8zS+ApOG5VygAPkjw5m4Wa3aMv2lbRQqQyTBn64zPlBBXS6Sd3rYJt9kXpaG
UVqlu/qcPz6VYeqsUYFzT0vMv6UaiJz6Kl2m7WVtGRMqr2/gtbQ92UTgwTDrSRE2zfpW+Pwlrs3E
ireAVMeTk60pIOE7TIK5w4VRLgyriuwqWV0caGlt2d+k3WskPwYO9QwaaX+2jwX0fnEc3HMjv66G
8vGj+DdPjd2ZOJ3T4uis/Zk7vMlXhqo366QIh+C9zhxR5GNigpcBrdnksY8Rr11+p+S9YRjP3yf6
DyZ+Hs5o2mlmmvVUlRbHzb9QqAri9dceDfUyvRq8nSm/EnE1jaZeQcaY8qkgceIpGsgoN3bNTGtU
wEbQKAYYcYeEVp2z/W9gKUJsfoekU1alg0m3naK5frSOT7vmvSc/7bDs2hxRVAU9z2jtd+KVT8bt
5FbWb33MUvbZDI7ZvyPP9UmCakCbcK+pvEGvi/szBebfvah8j9DA+ttNgrlgxEkHXWPxIG4oFKxp
QiDxN0NplMWpqZl+I6JwwdiZZoDg8/a1i7FHki9YR0Qcs9P0vm7nby7Zh6rTLlXEwZlQkaXR/dAU
Ja7XqLgo3pwpUZnEl1EMV/Fjb2jUflXCfutwtk6i4CYQFqtotrwZ5uiikqiDn1kl7IRHXpjyz1zf
3/DdwEkbAOfG26Gg4Bvkrypd2BiskXegzPa7tVHmVhhEBYrhM3aLKygLoIfJSxl3NIwuE8sUzzcG
FEBVxZdGN/Q3JmhCrLbmGPW5xFgFfCF58HyvT+V3K6Vv5xvnp+s2zWnkDgfBAG7w1sPNlr9fYprD
+70SUhTfQp4tj9WtaCOmDea6ZObKMqqckEeuN25J+FcUKPFDpk5Og56PjIPd0cmB7q7+OC5Qdfed
uqTQhx3wrZiLhoZDY+u2UAgsAIZMdhxNNMIGqnLu0driu74oYoB93fQiJeoCGNmFpqVbDPFWi9iv
85dGhI81E1+itsRKsiDbx+zAyqrFLD5jGRIDwK0dlBxkbv5+bIC9siPDLa+ItETduze7pIu789lU
VUq/sI98GGE+pcg6O1ZzWSggZLA/qf3Ylb73lTShMjxdVQq7vUjjYWpdDRIT+sAqowd5jEap1BKp
lLkeN4kp4Ih48h6FSeB2ip9UTNtge7hYz9G4KzsYPH0qXPj9OUBa4vjRmV5cWDHdsT6nK2OFxpsJ
84fdxc1vjkHF5p+UBf53mAYo9z5Veus4PcxfgnLBwj8h/hGebY5G9XBRL49b72CJDMaJR+07dnCC
IlAdHb1FV9/XOh43vTiAl0BcSb9+Bd7c4Rsci1StBK3ewMPyjHTrEM9lNn/90slfU+EOKHO08wkE
77sw2oQ044hZHE5NdQez7pcIJNDvSqpE5u/N+VT9S5Zh6iE5J+NA1yVGHUABHNWUxcwm840xl/Mj
dyr3tTxiEoinsFOvIwnkHb6AE+khKLPfujGyMqnt+DQTkfuKv+BhGT5vIpB3zdgNPzrDi4cS9owK
gq2MLzkm7wscLILoGH1D8SV7qn057RbMh/wqQRavsp450dM0JqEApyVNwn0U589bfIksS6aaJpvH
oNHwf8iXgzL5Wi6oa6fQdANl1BDbg2wYlPNpKMp/Gr6O9FOVqXLDfvQtZEG72H9REqADNPZtwKBY
hpvSRQkrsaOE6fT2iyfvZCSDlLDUvufdWnzi3jI3NucwAEwE41cdXM/xTNSMlVIx8MCYC4B9qgJT
UBrtjLBSKhV46oaPZ1oGIrHATuALtvAkx8huYaUTo8IVSWqEptBuGAycHrY2mHF/nVZn73ZHUdFB
FngCQjL7PPqnmIQYPOqM9vg0Uco3Q7WG/5+/ABlcQlfxFp+CZG20M5Wt2yhmcg25fJMw02/KqNYm
Vx+2t9EMpdlrF6EC2b8nUvEQEZ6QfIU+/FIfAeruThN58Oz+DBdAFU2nDoUKtA0PEqIXcxNkViwf
tdHmVFLhFNiX1voabTRKk45zvVxnsiLeNfkBPLcTA7qjGklNT9C8sle/hIhImRu0n3IMwU826JM1
sj0E/GmBuE+nwwPQcSC0CnsFTliLGesyRa6FXA925TYNrCXgTerBF/SugOaUge9u3DsHpE3pp2JP
NLsHdI18osWYNZZZVHvtRZfn/a2x4lfMdKM4+57drUbAGQXYZYqPYNNF8NMsL1gAFsO5thrfiJw/
r0S8YEQirA+9v4QnxiMx0BSHzNe7JKqs7ttSSujIVFvBiMnylMAgmkv9RDghmTTtGQHBwdelM0uA
+P6BKrYeM2t+qqNMEkzBia60PCAR4hSLuIumWeategOn3SaFjuYbPlMix7rM9sMYqCxNRCDyLJyK
nL8jekJDpMaXQxU7KUPT/marNQvUTfAdOBYInUKfFdCt2j09kHcqnAg1dIrathLzHdofk28AvND8
YCDQaiq251SlnJgz563ow/ml7XM0mCuUVACxdZ32d4MrjJEol2hEFZzY9FPFPGrQeScDgMn+gXO9
b2s4PAnUKC75pdXJNNsbXLRVVVSV3W4qTBwbpWXheaERA9Qx7T1jF6huIw14qrnNp0+OF6zeZdi5
eCSigrkfwr19jCyy4sttt+D8GNtaSgnQ+LDIblLwXoi36fqg/B4pl9+xU3QrB/na+r6gQDa0RBZi
sZe88x8ZONu7skdJUz+ICtLf5dDT66uLLRDTO9aHuiskGkO+fYCL457INKsTPuR85vZdlAxTat+j
coWIUsGdnrsLtf9ajwmHtOvOzRVkbssmMevHQiri8hrSl3wkbaXaRRq3z/rE9jZGBZR5Pw05iFPk
kHVXw+Q02m9Lr3dB0OkIZ5mKZG8lFYmuQWgCkCTHaMV3TpcZSrV8LfXn5xB4CeZ/Og4dogT4d0ls
bndCKlYCGTkfZM5YhAq9bGA0loPsu1i2R/Ij1nwl87scg0JUmRGXq49KAP92ktLqHSC/inLVIdFB
nnM46ye3loCejb+84wFG8Ddj6GPFCEIforrsqBM9fj2dFOrGgpw1J0XyirThGuhoCCXAdDB025FI
8w45P29FfUFAQgkJiq0hvQf1cXNLSvR1u5uvYVGwo1NyG7fOy+A0BFt8sAJSk1ViyVwZunl6HLld
tdqfHem44BwqO7MFOmUojGw+6HdtYJ0kz0G+74AWfUyEidQPaZEmRMa/d6Kla/zJDMSYC7JjJQC7
/IqJJr0Tkw/QYd+0w9KKOp5cZgn2Nx5pB2xXo3NXoe5KZbPC4UqVMv4O9cfeX10oxhk6MfcBXhW2
0mUj/z58r1LEcUZW2aa+0to9WvICEB7hAvqf4vPnr9+UgCRTBH6OuQF0oijUbiXK8HBWX3XpZdPz
2+NKdKNyuwoS+zNa124Xo1dXTtcFyA0JjX3MDmo8lkrZojAGjtq3mVtFlAkycH9HDtOMPGHaJznS
9IbiPgRcia4KEY6EZFLuEgD/eYZWu42lbDrDY5+bfED8PHFvpDygcbIlvevKMGFIkLuh9afkiy0S
ZUxB6xaW0k0uioARxmBWRW85rPaefliMviWqLMFrVVy/6zSLLIortyhrMcQzmraNBgnNr2duWVPF
QYGEwig6Za0Vrd2taWGKQp33Ml0agF92f+sBKWOIBDZbBms1onOzRs6LvPNM0op8R6WVmJ4E3rKI
N81MrqQFqUI39THfH92xgIfAKslhHG4bXjkmp824L2aHPL7zbW/gwiMfoTT9MHazwuk2pll9QMm+
apEibDf2S+IBNKnBZFKslxrj0IOevZAjIlQdmaaxHhRa1wTABcPqnPhve2TkMJFadx/rTHrwUMfv
fJ0mt5usTIecTNq4FJhVFlma2jo0bSdla75+Pc+bfG5tOXOtHd8j58S41pDQDHvhOr1JJGXhNr3e
tOhZH03lUFCWi86ZFBf5NwE4FmdhoMBFz4Z30DHWJ8tkL5n+0BbEbt8xv+YdpuTekjMW0n32KMyp
0GdnDTplLI7zXGwAf/sof73Nz0s4lRxFzJEvMJqgahdPn3eoLID7aybeBkrWDnvE02xvz5uG715d
a+K2dnYe7YEL7avpnSl5EDJOW7BvFZ1uWCrD7AbRy8+uZpjrNklBQ00kH3ALNqSgj0GQFx8ospNI
fKZcbDuiS3JKvgdJayS/vKsbfRV7iElfJ4xhPDW5rIsSx6cqtCpX+sKN7n8eUAeDsw8Un943xQFQ
Es0t8UkiJQad60oBtVt4LAUUxGrcDZbpdtiImomC07BgQNlOjQJrdlJqxq25cHyS2DdCegOaCraO
RHXxuse2mohyi2vwJP7V2QgofUtf0dJpU6Bl7dUFQfngRmU1Un6WtgyuVEIEQmBFYV8aD2WPDLa6
hNnleGpnLP6gx6TwZsuRuazsudy+qfnDsYuhzF9P+umK1ALEX1fAzcD9ITMXI7kXjnmdKLLuNf3C
XpbARSbQjMuyVJkYoY4tq4QFc+1xiQtKkCe9nMM0pA0/Z2FFjMnf4TdpY+ROb6dWOef/6loEzW6j
RJ2TI/pA/GisWtLjWrCYOsCAn1tlVXia45dFcPzIqS3j6XncQ1m0qpG/NWMIafr99TLZmjkUJBPy
YLI+Z3T9h9eVgHII1VvMdguEGCmJK+1d1vLpvY9E9AOo/ZHyZSxBk/lCMm021e4RQqzXq4I/k38b
41glXe4oUKpdkhlTDgsWegmQUl5Q8mdmsNDYiA2eXe/nlY6YCKxx0fopPXuMx8+35WKxvRMOqrBI
BWwHriX9PjHvvCXntoAKgzysfzqorXT4hpYFvtY05P4l6l8DwgBs2QBFEfWzKaBLvzVqC2QNnLBE
33NQI1Cne0nmyMYRim0PtZeK6OIX5EggXxG7xu3/aX6GXd9+8HaGdg+uK5zAXERxTZ1gSK3vpvBa
610z5O8wVOaTa2RHE58ah0Pz4V68gUvoPK7uRaJYgcy6VOSHY1+pC6aml52cMJnyaxfSL5iEAXuu
IttgzwnP//UcBF9qn3Cls1ytu/EfU381DOY5Xp3FIF9Vtukdz3PC4WdsETGq1vDxlV82JRz6PlXZ
ML6z9XyuC4GHmoK4skqmP5bsl8f9IwoIH2erFLr/tisJcSQZYTTAEosURviB3OlFysPrQnOGnUG/
ZEEk764e/si743a7mnJAt4JS4t+HISFHicZ9Cs8l2qJUevD3j+dIyy5t4cw47zwtwQsuwZO3JNvf
baJAsDpaF3XfK+I3gEsC5rFu9Y1zbXzotMbDGrU8xUZDGvFAyX/2RfD6qaXaE6UEosc3qNYVxKAR
ZgD0pU8ewPNbnYvj2+N7rbeQjjQG6zTsth9F4l/1JsvMBuARaWO2hNxB79sdtZM4v8YUF2Ysx7gv
+MdFkmSP5v5qeAnb/8giTst8+kdv5MsU8qFeqORnq9VpS+kMZJyXjNVsytiDv+VIjp6MqJIcULnh
RRrN/XVt3bcmvZAr1PLwMcJP0X8NGaa/QHng6pKogOcGYWh2p13Q0pip9QABliIoP0Z+Nvxehhzc
17IiQkZPAb+t3oYOifBLEa/Y3ztl8Wl9O+vp/s2AvH34TdVEwhdxHdGGwghdyYPYLEJDp1q4lgXS
MRnN1ZCbHWi2Qwp2zLd+sCysfOYU+TCUryz6Ny7NarRRlsab0SlPpvY1fZyhi5RQcUTCHWLfw8Ft
xNdpQJGyKC5RL1f9q69era8bAfhSkvK0whYUhJ8WKMewq72r2ylmBII7uhST4o6P0tnqYNVNRGlF
2dmwRXHjjrihzTyGsULqSR7DjYFtXgLJuweWWlInDG2JbQWYBhhPkKtspSkOy8KEvOPFdn4t4LuO
1PqlcNR3vKWLFHenJ7zG7rJdxHzMDxSWgtcuUCkbHnjkDEiArudkwtlP+LJ1MbVsAaiHbKEXkP8y
TftDeiiGnOCypKVyCW0L8wlRzSRKa6Z/1u15jzXnGnY+CKpL+oKJ5J6Qg7dafPfaBnKoeBRaIVx+
tq/6LhgCidNdRlXRakcR5vOVoiBr7vPAzhMsNyss24tCC2VW3SMA3GRYZKV5SABLkVEvajL8NNT3
Wu+HMf/bmYPbWFdOYJdCEoIRGKPYu+5LhfTLWixJ6mzHZh6JDY/GBRbjwOJpT+TXVc3x2dUmpUJz
7TIRdG/YPUfWgjDDWkS1w5jeoC+8f6YfMAS6UHLZVqBeJNxqPuqI1wFxAigVnN/kj22c/WdIc6HN
kVkYVWohwSU+J9z0TpUWqUspRPnoNuT2hgYP+xH0koi9I2mJ/hWRba/9oQtLstViygTD6h1gKff2
T0fewqHfwp1DSxXlbYTog6I/hz2sr6pHmpPJFALdiB2634Z8AyZ9ZtkQbLr0A2OnopzxH0XyTE9Y
tD+JUqjEC8DqHAf5OYPKQdx6X5GY2a441V0pPW9ayZOeU6enRDvTgsN1hknbAv59AZJVeCGEn3p9
57kdaIInHfMZONHmQHDO74pyi4NBZLJmLNTmc9ajC8enJA5M6LPfCzR1Ry3eDSCn7fyG6sYWzKx+
Wy68AWLYDzT8eo7AHdfOBGlADfFZDiwLFgsjGxWHirIVngbcl/P5S3ZKTglJUePk/mrOZ5xfipha
wocWSqe2iNhvFDoEds/x32sBZyKnNHO3MFaxUJR0HgYb6VsHWa8uiOuVFF67ohkvqywOY9ERF6z+
38l+XBJXss5eF9PNRNrP5muAe2LO/WLjrb//331X9gx0YOOF6U/jAXhcT22BGsr9BNxkkBvjUGgJ
j7KlNtq7e3kPWBZiE4kpfjkm+YoOuGh6rpYrVbNQlbf1oMIHNHukqBsZBTM9YxMmdy/61B8q69Ju
D/+zpkFzFIz2h97n0mWvSAQTDf1LrcWxg5UscRQ7wiMjthldQu9dMhJY0hOAJJCVYhp66j0SxPpg
QY2OUvFa+lJZRLaV0tFI/XYAmrW5zKJKXuisSmhtKphYHPh5aCdDjt3DN17XadEZaVKEhX1H9zCb
5u+LGCPJWR8uJ/rpWNjtp0PO6EqMnbwjniEYTFZkj8ZvvslvhxuPoWzWQ+j7eOXr8VD5TUbSAp+a
RB+/tuakBWPLN8gzfcSSoprEydB9bBCUMt2RckJvTFx5onEDpRkRR0KA/U9FRBxk88hpRiQbOJ7G
7WdtZBWkLCul1467YbIGSuLd7xynYiwK8r01+mKfqH2jjbpDNIPGzKEsrzGjr4LvHKOX/QZGZLnO
akhezIMbaegHFAOQexZx/tvFWsOnXS+tBYbsPeODmBSPDb0sXdpJBlDhv0540URdePizwypNgb0L
jq3ERWlJ1Sh7m6VqQDH2yYsUrI0kdEIpDA/zBjFkAwKhgYJZ1g0u1j9oIjwKBKs34s1Fp1VvzGeh
Vs/70tmHvw7tUdPT8yAu+hBCPkltzoB3sfWZKfJCUHUPvF839AXpXuxV3keu6a4x7GI6T0i91hm+
64XCvkfJp/Nislkg5RxnNcdCLn6gRDNA09od5hZSF3a9HKEH706ftq809ZZQx1MUZhVnFP/UdSye
vs5DDl1fqDtD1J1jZhDQ4E1SZMh0oL+UWc9U+TGik0gJw3P1w4oXmESksOgMoVmKWxYgdre9TwO+
9FxAleRGl+8tk8O604VxQobLbmuw8jwhFLWt/M7P72lGrPeMT3cvI1O7Ps6koanbvhAV8ZXjjC2i
MsTiyqb029s9nBRRmR5aq42vTIonOh/WdaWrhgj/jdRA/asusCy0nNTu3dIOY/jHja5T3ZZnnbs7
lyDjlNUP0dulIZpIKJhy8mE46I8H3M+GfPsUtacWscbeTT2CiwNE9X8VlDZrPTCILmp35QPlD6tB
Ziau9EkLAuE8DeWs/lb+S5USOjpPQ2KbA93vVfqeCGd/mSNsXaZMCgw2HKikFqxE9YuaTx3BWa3D
pCTbQqIU2xv9K8Sdi6/CLB+PqRsh2P32FFNK3HLsIDAwJOgkDJqp4Sf6UQgo9S1N9B8SSxqRnyFh
Z2Eyd5jRF97yV+6ew11W/5OIc7tlhkbJ8Foto4d6Bxmy5y6UStADvy/8nKJ8/4D4Gpcrr0va9NXb
8Wvtp1krBm6xpQR/fAVfn1/RtkGviiWmcKUPyYh9aD9VjCDlIJdmgy0OQxLd4Z0F80qakTg1ABjt
Qw6XbaHLmtuqTLsGFrz3RJe3rgb96gfbRQskQpP8aKjYDUAe9GaKqLqFxwP+m+/0qqff/Ur0wCKO
9cGzg8YipY14sx4m/+roqg5zxzeTs2wlDuRMjxt49VRNKXwgH18gA0qgwP0NSqasa8MbzWYFGOUw
aTEMWgbzIbUdwI9OpzlOsNSW9YrKoG9jwwPChsbnjlpH22N5/b4dEodYBObAtISGEy1mNZY6OkE5
HDKjOzZU7IdvUxGJiO86UQHNj7Nl3dcuMOdmz89CNIQOib7f8DQTqnXOKv7+k7juUQIs2AOdeTYY
UNYz/lxJca2t2Gw9HDrnLnQ2KBKVyRBnH9JqpyXFw0n2Yk86taKtdwn3sc7vMmOjhO3N5Rkn4HJ5
XR32hQsoxOWO5CyL3T7ncZAeTPm70diYEYXJWA3vAHvH1Ituy3CgPdGQqNSvCS8dPRNXU8ityhg6
YU3P9dXof44OOaYl+p+wTi4GQa9YJd9lGebKkYUhy1IelWc+r3Q0qF1W0MahTeNX096QWtO+f5Mv
7MsuBCcAnW/6gwUDaaYNWFtWh2lmPVnML/kUBLbZANJ+4f0ctHMkjBA62jpPiDwxyUKKexSfBt/K
5RVCMU6sIA/6wNXQBs81LG0ZG8osLyPVAolL6oGX6ONR8az6Y6htPuqR50hg4cN4y0xy4ZxODqeM
m3cwwUDTowz9IfL84XfgBrBLRoS81yYixppr1VGeucliKlBgtzhmGaG67V3xaYS46mTyXvMPrlT1
RoYJ88rHpf9vHyJ7/WhuGfxkcTEefmTJKjgl3nbHBZoY4EMJxDnob/bBxgAsqZOHSPfnEpFICDbn
vb+IEEqGwtEAclj7ALWXcRAxbqfG70lGmanKVRigLIPJojhO9W46xV7fkRZY3bih0io6sw+UX+48
FyXfIxNUV0pTE1IuFAZ31kL+GVnYdIo1QBHLlg/HDGjb4uK7KnXSsrQrYv7iIyDEeyRB7/2+MxGt
mVRjtUvO+K8KQRRtOIqdh3nPNBV3gxbfk1vPg7xp1VAa+fq/8mrmSbaeblqSnDnGRZEzq/+h6PLC
CjjY1RQCAVnooht8T+xUqu4LG8dmV7GSbM4yzrJiuAo6erxCrCr/FGamtiISgGjEYE+X9jBn2sto
wpuPyBkFFrNW+VQ0OJNccBRIuElYwb9bqCpyt74QakPwSSC0nIEwLzJpkbDlDwErR3Z/lrXK4v1d
uGVTOjZB+8rON/csw/f4/v20xPGan9hr/ulEw5IGTxBm0GtRIJ4hPX3eCl32P9N/JQ4vDrdzLQ52
JpRii9GDACMmlETe8hk1F4o8JTEpuveudGO+ihZn+vi7p363C8Wb2w78gg0p9wtp14wGLzcDlyr4
jZkpLQBdlKgDDmaRXWVD8pIB+/V0Klvh8nS84a7j4iAIlS7HFvIsgnynM4DR/RQD3QNMWhLIbSq0
/6jt3EUjaJw6GpOCoubVgGFwfXS44QSV3lc6eLBnk2TkKya8A2HsiaBNwx4e9TZmuhSwR75XN2RA
xPNO3brIMkbuJS5qLcmNJXtpjdl7wTDKrpKUlPXZVUxfJa6pNV6dHAWC23ETKVD/duKVR9kaVSsr
JPILSdfBRmryhHBmtN6kwvs4EsEI017Cx4wzBb5kPqsVOgSB3fOCOBWuTsqc0bCZd1/w//tWarPi
jYRTYRbZrhSuMVOb7E78ruDpYOnCaCuCqZ/NfFSQtpneasGYLAWfBWXpE82lHMTn4dmSyC7Amcfn
/WbDyYot9TkZ8yy0/fv42H9tkrLbnBc3QeOhV7kk99HYL2tbWgVPPpMIfpDfZSQ18oxvfO3q5SwA
+H/LcGLc6aVWFBMYYThrE7bIHfLy8GtQwV4yrfpqJXxPcwiAMzCV+3GbgRreRl5/KcF9SkbiWbNN
soti63PKpuQDFpTKgr38y+zDfSUqdhch6B/SlluMZ02TIzpWUqOg7sNUh/IlgA5zRKygEhlNxVtq
qV/sNZCo5N/uL082E59pP982esm/s3CMCzI7k+t6n8UJc4GK/AjxPjUuRv74SV2OZs+svGHJoYq5
rIpyROtNfl9OL7bGjpCt9o7M6xNESWw6H/+551FcC1rQH08cmfNQcGhLw8g6sqm56XZoKx3kqdfq
ae6azYo5takdqw6QjYlLKW/oI/8fp8A8eTWtFD1P56BRcev6DBB35LvIfMO6yuVOsE7DMNj7OI/S
rlepThhoL86/3rFzQt4z+crbtPopPoYCsoW7bnK58kea/XbiYz3ej8fco5gAcRxjPi8N3qwxtpyh
sNAbLADgzMUruLR6H3m2/aKxbmfAW0xy271RalXSj/x15ud3hPjPyPNEZxqHL52VpRSjQifgEGKR
wM1pFlAt/Cpe/wzgcVD9W1gmkIVPHcdrT465PZqpOe24/GfS6SGkAkOe8nyqF7vKcCZnptjGfY+A
sheVHE3LVDSAkgJM5MMru2rzV3QLeXFZiyJcuVn1FReXnoZYjEjdnDKsGhlHaWUEnZ3vkdn9TZf5
Bk8xeW7lu72R2AaLiYMwhLA2bzzKFjjIAYo2VkTQG119/NxiuDQLJKvGiIchHA8LgvV2F7+/pu+q
/kxDnSmO8xdV1nZata59j3U/gibwxTcwbdlLzZbY3LPszmHS3Gg5I447Yh2nL9T53PHBis1ukOSD
jz9Imi/0fixzQ/mJjPV2nsRVfUtxKfezg0Pg7zKxaINfVfUeQT+strNlAFyS5xDtb/16N+QrOkE/
MmOovq+iCSbpkmCHlvO11WFTmReGeOixldoSPYyyCyDPimWf+RFD+t/1Kk9dDXVIwjGFYFnvHhnZ
47jLr7eWcwnpWyMVRUhs8Uw/BbLeLtadT6R+mEJmZPsaMjM0oxleEh3KTRbUWN0kdtpKOh23zP1E
RpKpo/MMA9yisDlGrcMHYrY++S+pS87KbTMMtFOHPZFb+vObTNqWvfhDbvO5wsnnIEUuojNWRAG0
77SW8GwQm/yq+LZ/2buICL6cE3w3ZpQTUPSBy2G6U5wVH6eoMccJr00UkkQ1ASIkEC89o00rDy7H
epOCl2lEGslPUfIAaUWFW2TcG7ZYAEOJQHhTMKHylz5LzuCoUlLZz0MTUxjm5hT2yTCLlMsmEZou
NIq2ZB5++/E2HlHzts2/PCw0NWgrEvBOPgbqfp+Lq3zYQH7eI3s/Kh0fPeC50Dqqdi+H3VG33k+g
st6AMy0o6tuj2Or4VSOTYw9PK/sFXMEFSHs0sxzU2iMQtu3af8M9Z+qmxOhERPLRGaBe8R12ZO+m
nGuuVq/3p2qu779nhOQ4l9zBFdIgUP9tfUqrKJe0x2LdG0FGxY5t8Jt0kNbDxIwyvekYvcZEz/xt
PVgJrGpSJ/7yL0EQ0HeMZp0xSSwDY1ByueOJv8A0+BkooELiBQe+cdGiBycaIlI2w3HLYiZA36rn
rINm/o1U8ntMfY6TWms0XlRU3MnPP/S7hpPBS34Z2fMM10pXxFJnM4pNet9HQwOgcm9kiWq8MW19
h8qZ6PBazgNJUGs+Nac0wL3FTji82gWbASjeSaRmzUPuF7LKHhJyMsoDJ2TNGwsVqewFOOz/tuxn
WiI0WkrM2WSxkWaboVNKF4e2o6wKijgRJ0mpmquBz9ya9wp7cVzxV+aFRQDQ1pP5Fb3orqElp2ba
E5nAfeEWUOSTGHNDTWqKIRwfdPZ1a0KWDJ4jm064UasFz2ca3S6ZSqWy6fdaP/mpKsnWGEZsCCan
02iwm0wf08lCCFoN+f7n7ozWBqQ+UOyzqodDrGe8jLEyqiSd4HHhtGAxaTrhtS/sBBHhPi7ViSFa
zOx0g3GGsul/Pz/l4duI+qSpBVfJNtaKgJwCEKZgX4lqIu/43aatCaPhveUSxk5fQgj286q/3PqD
kSGNXggVfHx10YHsZU0KhirWojMRfgglHh6BKGbPIMflpdLANCd/GIvGwl/zu0aemC9KKl8VOz/z
cYK6nAl/hcZua9B+cn5zGvgqH6PIRFcSReagOy1W/0i2vg9jqWbPz1eMLBgQ92Iwnln7dNfZuTMM
Nw84kPqUCvKFxPlarVrYyYRVuB5YxT6MWxOLXyUkF3xxA5o1dRRmVAI6Ml1E4mDGBflDTTxkA73d
CVeAjSqUa7Ep1O8k+FBxATT4ul90BNKVUqoMB6L1bQ2BK0feqvFjiiOO5HSBQ7c6tPj+bFoSHpet
1GO4QeiWJYVt/WnCTscKrpW1EL49x6yi4C+yEe2Eyb/DjQ9BSxHzw82UPKVLx7SRfNU0I9+VYH/u
TdAofho5Q3IfOZzawt4mBphaEIIZ4PsEPyxet/oe/95eHMnDiq7m7fomD/LFOlXkUKevgRAzi65+
wpw8r5YOG94BMp/9SalLQ0FYMy6W64cGdMOls/6Y5twmNdP3+CtWc2TZMnu80Dx11ZB3nT9au/VL
b0clGj58Cp/5rEiqrMd5P54aEA4IFBDXDYaxK0jEm+MHg6HytRXnACJUZk73SEp7oVBdpMP2b4d/
5j+A8V7GqfMiUHfvGW4qN0XagCUQDO/rpGCt2qtHJ9UydqcxNaxzPlrkFMHT6ME085ftbmR3A48D
v7kXAXqJJ/iJ0IiNT86v57zAxwDQQM1Rk220QDS7bK99bjmRDHODCz57aCKQ2+ZfAMNmzUxJ6wwc
/KBb3b5FrBMyTBk9gx7Hli6p9+LuV7/Z8RKpzAGmFtFxhEqkjDKclvhx1wFACDufnAKncIZ0UES7
Fy6hflulPx1cvu+7janskwhBdugbNsxFShFbP/H7tbhmIrE1ZpTYkUnDzm8fNQNXULaPxS4nyHdK
9ZCqNTCGRlajhDxb0zldUrmks763LZywaoR4L3i0lUujV37FdWLWnux4hXAJUTovjYdqvlju9Ir4
K/u8od3EkKzMrHj/5qdOVQLm4qKgrgdjPRFVjDh/APcGRSMW0TiTcfaueOqH/IjI27hlkvv2Ww62
18SqJvboTk+Ig4O4gC7wvLp7BLvQ6BMK8DD8cP5E3LU+Yi79MbVRFKAFlCyNE1iqHI8/vBb/LH8T
hUw+7o7RoU/T6jffWak0PBqothiIdR6g3oyLcMUBK5mc0lhj32ALxYnDkOMXBN4j8s2LMOBp8utL
5nvuIrUxBgkOKqWI8iNdGBNqpTAFla7fpdB7WUVfkVXBgTw/k8M3/zSORjdfS2pkv4YVwFAxOj7c
+IMgw/qFrnAGsMpBQDP7TuA2cbV8uoVGqFl1sWw2Wm4GAkT4SFFfSsPBv9CfmiN6QUVQfLCZfi+Q
ZkGXNIBxcpLF8q7lp2hmVuG3KgkICLAFI/O3k07pnZbCdlagVpLrwm6iolYk4z/11dB4OVvW7hzv
XOnSpW7E/MT8G512rS72lx16cYNcJHI89Z1TMMcnwK5HtnjaQYin04s8a8lShE9OQTRVO6b6S/Kl
znABypH+GIEF3wmK5XvpOeG2V4fCKN7W/Jp53500DvShLre3guJaLAQN+Pd5EbZP7e6xxtV2qSxG
ZBBTydK0ZTff/pkvC/5Yc0UYk9GiDeQ0NlostYH3XIpxbX8RL27zMcxdzwL++vUuaAp+hmNQ8lJ5
hXbhQlD5otfObEK8Km1ZbNYvEGCSK4psTK7Ioiqrjb11GTgPwrOUFKM7oiN+A2DoYyaBlg2y0wTF
urdIAEsb19Zt9RL4DmTbEnMSslVo+TSMEK46mr7GzgAFkHua4IRlCuu5UZ0nofRtll2vQL176S6w
WLTLvA3Yp4HZnzAnwvYYwKRTIiiSCnP+BcplqDZJqjeTTVXoGYLXZrrat2Mu42dVAvRFxtN1y2Wj
xPK8tk3Pts/mcoD8yOh2ei9e0ro/XpJhHPeA54hEgibh887wzUJwTOwA8RWmBaRl2xw8X8gwAp8+
i2+kud2rbFARQb+cVrKm7+uESx8NLl/N4jNNcxeYkFpvIpx1RRsyHRVXMS8t/u78CD4MWxY5QoDZ
Oq0MTjIUJ1KPX/yHfNqHqBNWxp5lmfdEwmqQD/JzNxcn3+1kmhm9ucTtsuDkxn8xKFeMxT0wRkWn
diwCIz559i28lSgmk9044ihmKq5K4paHCbx2diwmIi0Ug06O6viBeuvD5zqfqNfD4PwhiLFtJK0D
1S+y1XOD1QzoCCBJO+TEeZO1PihzUFLuEJSav3trz9K8LpXaRGSh/pt5LU1l2Z9/fLJKHPf5mxsr
L5XiX4aKwQN9y9BOc/UeTXmx8xok3onmUCCLCWAhnjSlwUoEg6SXORH2c8AKBltY9hZv1vCwrBlX
uNvRM63mfCT9ixo+JeMZ+nYKZJOzI/cRr0ysC2bn4CYPG8O6PN4XZqifFF52yxU1mivo+qBa5V5f
xOGvLD8YmqTU1NgeWNqPWIWPSrESfW5uQ3OOAPODsMaFWYlB8MuYykikBsOPnkYASSEp/7YxIoXt
OdUnQw50sroFdKcrBo6LVZjkVLh2ud1FzS8AwpYGVsMGZGIK/kMzNFT97Ceg/OOA8h9N0qmsEBnT
B6+istFDUzAEzZdM6HUZB8rR4/v+R+sesIqsDihI8IPlL5YAOlnyIHMjak0d1xDqLTwzFqN+R1tu
U/fOswMK71qzUfwU3tlo7drFG5C/9C8LYzjZIF45kLC5AmjHIMwGmlLiHmAf5uyA2fF4dE06QCZA
YwyFfF4AXtDQDR+V8l59lJ2Z1U0K7ItUhKNJphjU+BuYAvx8MLpF5TBFrqnjQ1t/GPQ+MVk1VfD8
wPFO4xHtYAsWG4Hp0MmnbIscpUaPbDfop66UhI/Ym6zknnSrYqV7vM+/pxuPMVb7lm8Z9HXQGt/u
e40nK5mMj+NmMbviJynxkxw9/A+Ab2dF64kESue9D2yzmMFu9yjOY9Vv6cZxiex7EF8JJUZCH8tG
m1sgc4blCPnMblSoLWZR8rCioS9GIdIU8oZ0v8L1rvzdZZH9R4IVYMQIy/XpHs2hG4/m6AymPXRS
dzs8mVxc/cQDKcBFQPvQClbz01bZz6j36BIQQLb7d2NEOwg3VoDC6k7Mdh262d94QSsuCZmpcazS
H7NRFmcCuT0C7Pv9B0+7vyV6K4p3zIy2WfJMOw9n058Mo3eDUrAmDxDI/y0hmfHeSycVoaA68lJK
NR8D4croszmNhhJ8/rBEUWCpmwaudHsqbEB8nu3kQuI34fVpRDPQnAo9+zLWHyCKpfiYrOQMGKZV
2E2qf61hX8hXndAgCki7Xd2zN/04sBm414CGekkp9QwoM7zWayh9aFAVppVcDWw82Uzu7BmLG01f
ZpSiE0KB4tb/m+3InNhN4gc2b2Cq3oMVx9a6OzpxFZNZbWY7PBH02oKkn3/lAZEHoWwPIqWBcE/Q
fc7Q5Em0589QuMEmXt8yJDbLr5browWmA/J7kZ0JARCTTTQx6DYstm3APaA7B0L9cutjGZ3BuIh4
0xPs8RbakS9lj5WGO8Z5sL5twiwdpxFKHK/55zTlPiu1FI0yJX9qxGuy45pN8ubppvzCI+1SoQgU
0luv8yM5HMLcmRG6CuSF1jzHP2kjmeQ9zQ+Uk46fgxdeLypld6PjSVL9MtilJIIoM/plJNKXzwGj
R4EksBet51ARkDump5qfllb7zY2rnGlV2TC2UgAbrkvRns6eBBCGedSf2YNZEhCUIhNoEoLZ/eRX
lY4zw3dXdcmUfWsQa06pKBiZQkVzCXfi507OpsfcNNoj19zSDLMWVmWG2zsVl1aas3KAiay/2IUO
bHwFczk2nxhZeTMcotiIIxm0n8Kye9MR4a24WbN6CKgXHFRiXOV72YlnLfPpi43KzJi6dLyUTFKq
WXwy60tdZ0yAfgtXjxGc5p6vhpzcEjHEsc7pzwsGkwhb8Bfo45IZ+pp8KDhrZPBj/ZIcyyPA7KoP
BxNZDLdUuhqPjJ05yut3XARH9ublctmB2TtULYAspFUCgO+D0gcCUZp0h4neJuL3YZK9SzzEbJzW
Q/h3wie502tN9FtubqsMxN4NVUKrVK/+dhCeDEOVxNJgG1DoXMcLpMgTZHxgxEE4emrjAiorTzUA
ac/OU5bJbZvmRWPRJntSfAwhdHCRwrNtBPjJzcz76df/FUbfScWD8cvcjojuR6STginUVJbh1tdv
b053RVHGhyU1AacSGCYmwpv8jiZWL6av5Hi4Dfoqvq65KLAes0Uc936cEL5wkSd9gN6afb0T9cRz
oplbCgYCtuQNRyBVLRalTPoZTkBA28tv73idXnwc5Y+A0RNJqjvgu3uXk18HMLX4aPtHki7hVqDj
c+fBdoOz6BPE3rm0a2t+dro28EKsYvULmpDNAELwWdcJ60vK6En/iiXLRSL6Mboz5C7Qnx6qQ4Ot
uugkeU1hq+zVoj+gwOrSuks39VI4ubyh87PyRDoGrZYZgOctQlwc15D3JXWlR2JLcEThh/hx/gHZ
EsYy3xwEKQMQRLYcMkRMMRR7Qr8EHd9KY973JDf1Yzh4MVdDyALcdLAIfZEaWAGQI4gSp/LrXWCV
OQrQakbGtLOnVAhdVaFSPl3DS9bKaStyd2ehEc/4j/CRJJTdFxuDJEZ39vfbOYlN8kWea9FmVsSB
ZDvERB4QWtRfQ6ij0hE7u9wkLOb2AacNRW1hQ2/4amGqMzLi/+/wUjmIFFDYb+BeJgAdaTX3XmP3
G2t1TQM7TNM0aSguL1VW/1ED1dP/l7m+z6CG4t4rLHho4FVs/UORhBtGtTtZw1cO9ti/G6AwtyDE
8woVvG5r4iOKsKihFaFwtxMKdU6xFDqOdjeskvz+R5QpIZujWTZcD0mMYG5qKkkZfhuaUCVIZH3W
NbEKKhVWOp0mNE+ahzOYntI2g4uBxUjqTKXUgpobx1cCuREGX71bMPHNFwQjJCtVXoHB6Ct7WtMv
rinyFF7+OFkJ0FeUTywtmb0fWidT1uXIPacJe2vBjLnfQwh1f+7cUtN3BIxQs9EPq8Bzyyea8FBm
9L2+DFxpSQ4BVa51jQ7KQQ5DfZPCY2yQmBZ/xqJymEMK0c/DdA/xpEToOLvLygM5VbevQfHil3Da
zcF2SufqjSngEIvUOmFiAfANXLWcXFthr3JepABQ462F/aYhFU0mRmQ6GGZIF4ssI5baAFjV7RAP
+aB3fMmy9p5C78HseUQ87t2jPHhVJ53Mjfbl7Y0dJbs9Ym5mUpB2yb4CyR2ccLQMl+SKY2yPEaSR
oy5Lk07/ENXXCvpEAASMZttSgs7EqgECpJ4crehdMf20k5MwmQG+FbnCaMo51Qs6EH9J692v7G4w
V55eFcrgYyp8D9LhtygSUBN+/aXufz5gin/yJdG9qQvb9Nzt6NjxcyNilWxdliLgo+uszlH1UnUq
AcwBvCtbDXxmS1F2QMt/m2MQlXKVjzfEbDCk8vxZGc6ku8G9Lma+T0ZibG7oSF65OYiaEJjI0kV0
AfL/nwSCBGFmKF/3lnigO8rYQLgMnaGX1WoJ9suBWWUCOy4JHB73+Vi+6geyTXgcQa8vsq042sfP
FSAdfwjfDKggYmhgyJueMaKixAMZuri2jdmwZ2wm/fl2wa2lhEd2kyNGwMJ6BXKBN2ffq1WsJW/n
XdC10YUbujJaMH2/b4dBb2A9ChqrhQGRobrgSGf/Kk8R8GXbS7RynrCZmn6Yq+KwDlg4Y5jc2xhU
IL8itYZ6JHag+214rxXuTww9GrrYn/9Gq7esUN3Tb1eQdDw+uPrkGNRWHME7izrVDnIpKb+h3ymf
oaSAe2RAfF7zWUhpZ+jyDaefD/mqvaBknCYJ3CY4IGXNh6TR0m5gNykPg/zQLz+MyOmhF8rlHb6j
hz4Sby4kaiuC+1bfY2IlrCC7LHKCZ1V/T25KGFoxGDEGH/v17sfmfjDgpWbb4FAM4kO1RNh87HD+
stmbVGaxfk2R4ZOIjKMa3w2XAEggky8zrs7IdaTVkH/YxzMGsUzO4hBZEH4Rq3wjd+jmBbj1Ouug
TmIdAbxglnVc9XLG5PxvGW0R5TKwo0cXoHwnYoD2aGGocjerqDAljva5OlFZ6CSVfWMN4jKFXKk5
vjieCFTKQcf56PWNINMEb1jdj95zI9uReWyTUsoDo7TytGy3pl7sp/iWhnqv+vz7Q35ktG+eiQTf
PgsNbrCTTcuBSBtrXnFcDIqWmni1z43e/O8h+tKH+YknimWoH3n5Ic66Dowt/teGw3LphuBq4m2K
ibIpgjdrkf+HPbesCfsQSJ46xABLysLiseejqOFSBYr6Awth+XuJbMjDpepeTJoQnycat6FL0ZeV
AdLUO89+v0npooMkCP4maHbctXcWinxCCjdGqPtMJn8C4wwMyBj9hxF2GZg/FrwrqAN2rR6BBEGX
k5/j3vZXxpXbekB3OKp4Yrwyk4RRzTmYNqfmJEzXvwbkrwDZSaSbEHKh7saA0XuCuZpFAh27lZgo
V7ky4Xs7P6zlxro5yDB4NPhfDkKuManGOM3TJcyn7x3JIBG0b+ZSjxPrJgYfvNSRa3zbnVPdWTOO
mlv5EJXxbSOusgVATDSn1JZkRHqSDG1gM9ZzTFfDy0soeZwLkbJ49bPLk+JEE8Vrp1dbIdu18Lro
w2Oc+d6BtBrUr8r0Z/KGadPBGJMKGorp51JHv+aRIePV97v1Qo9X/6I8vCr/9kx5Gt75OnoQnkdi
FM8dbPHdqZauH5ttBXjpNxTsOMyr2lMck4e5ugHuCOopp5KPAyIxTnJ0CQ4YEVvUjBRrKkJNAAh8
FENqJQTPU9v4gbva57WHI6ae+6onXo3Mf830rgazhqAq0N8i4s3R37H1AtK7VMlJrGNWEGC4TE+6
MRMpvPDagcufA1v8MYDAkz5AdVpBY0lKqteXyqCMh3Xrud+yJlDj4EYDDN9Kt0ZpnLXlYHJZhQ/L
+0AnOPfOSpvLGUS/0j0i83CErwpSvbQMfBDi5UAfS0u7kk6olzvyhS8Nkf99nt5PoWh24aWL2f8W
Mhzf2ONcNn0BYrXCvOT8a3HPrDx0j1ReNo/JF/TwJCeaoaH//oxZbwDcHG0SA3AGa8VbRIqQuCmT
/QYMvjYDrk82tqYiZNwMluUmLTBuMX9gkZDTPyBg5G30ZZjqRbzf9j4RSVIpSNo5QFxB7rwAhvaI
y/j4YOAGfJcNDLRAvPuXRILd9NL1kNhIDhcZRF0dqlfX75k0Fq0WqG/Cdlot5mSR3FIA4h0TsnqL
4eISebHGmmSWFUoRDw0QqDmo8iYTuGUUzMfmC4Rc9DVhKXbpigq62I91BItdlnG+ITQkpzQ5GxEk
+mA8tAtr1IJzdHclD2YghmW2MDms0j6/u8OuPpBeboErBEIEEg6dFLc9Z+p/rY9vTJJkeyXnlkJ4
5cKG+Wz9gZ8WV2QZujU1FJ61S1gBArG8mwPs///69uvdAv7RWq1wNFy+UU6xxS5xkpMQ6PXEm/Qd
LAbUFkq2r89xVrm6J8Dhsf7cULjxbqhYyHBcNnTwPcDlhZV1m9n5/SoaM4El/WJVmzdLuQHfGgO5
5+l0fEBCdrRp8PRHErGj+FpaXBIcfzpLy3D3IaOuFfav6DCcyyeK7riRz6Sv+rsHknsHxPixo9aZ
XcLnate9BXF2P2ze380UFZeiLPA71c7dkFnb/Q1Bz6Z8vsfCTT2G5pBg8ydtpcLVAKsceJM8Pv9p
R5KQOG3Mr1Sv7KnbhBDfpBeHQZMHYYNzBpvjpZWDBimdMWnlgS6KhSMnoGV+emM6lUS2oQVCGoeg
qherGT/IlClNYBnUvMUTzdrOdSNyozGXBxSDTzLH5gZtO4GC0nUlW5/5h0qEgS5r9FJf96qG+9ax
uP4juqxprDCFJ+Jizr3+gxvbQhomE4yVif/jmQjKOjYfhCc2EDkjUO8sOxM/yp2gg/d3Ve/U+jrS
Pi5TfKwRFiERrI5LLuUFFoKPQH5VXVUiJArfKCYgkzd8zuSPN+8V4f/p+7xodCxUY5ZZm1GtM84y
CjMXGeLl32KpZI5dx1Qe6BFP74GtQ11AMy+lvaWQttXVQ0uTLrO0O0i3wDoVX8eSkFlY/bZRFORc
8/ur6J7Gm+E4AqQMz8vqBEFuRYKbHtMUxiugndTJIqx/mkcfbrYp4o+7Lt9vO83NMP/ZSttENkW1
c2zFg2em71tXkVHQep3ucKOKAmL4yay/mfizNmjFYkBEC5JFSR6927/hmC2x7P1nUeE285IMnXLk
O721l1T2YYUzYZxrC/V58gwwppP58w1kPFYEPITZZZg76da+0My6G66x4L1/eycFTZGcfCoeQGu2
o1rf2prFwrH04Oc8wtyPqLb8oPSy8fMr0r3J4YA+reF7HYElRxpJrerV5lJeDsUZX4a089RyKlWi
1c3VGHX/OskO1q/JHaareErYXJDD033nWd0rlLdel/y/5sPZfhaCzpw4UcnG2qWoOxN0bE9Vo5vL
OFbUvZGaUI96T5Il4BRI1Hs2NP2q6I4TFGNwiYKcuNnBfKMnpU+TjQt0sd3+i71mL5QNEgG2Pf14
/zMt+tQWPw56AtnoQBqxA170E/dIiVqyY7PAxMoeaGxuS3UP1ETexiOAf6Maq8z9xuh3b3ySqBhk
qHqtmwWO0b9YjXUUFIEpTHXDiZktUXiXTl9cj4WhTw3QfoWt9uzTraqYVATB0kBcJjeGrv/ESAfh
bzPSfIFQZmyGB2dhJbkptmNNijagQeiuRtQzrlnpEfRKTfwooEa3qz/SrhmOd5WuAQYgXAerADBD
088qIbY+LP1+Jm5XsFsUkLTUu0zp9lkjWKGMpeMVLEP+8/wZG0jWN4xPW4z8uRkyH5bohrNScB51
XhKrXLrUhCZdEpJ1VAaBpbKibG7kumGtcloQsggwx4xDZPruVDAKuYT54Jw3luflyTXQyxNYMuBs
GR13pSfr82G8JAmRq6c1Fn8Ehg7X6Dr7xfFr08BSpNeE+BmMj4EFudyHGgT4MgUAoUJgRqHeaBM4
9c0g3852eOGpxzfNBm0clztZm90AIkPYHeUnr7mucAWV6JyIlM4xTpzL22UQbidy88qkeel50o49
L+Ko0llBcM4cR3qafOprYwmAdPeLkpje1LfRfNTL2GwAh3gwcl2T6BOjmU/HaN7KUGB++DAHUWpo
yqCMlA4vEbO8B5m/pw7vCoxO2vfvbITpjlRBltkUHfSDliajIuhmH+XhCBqC29gyt8oEtrpLjGI8
C8XqdVnhllYJ3N+qFtO6KFmhQ+yfm2VqEniF6o21LY6KKV8ad9f77ar0tiCOE8REZG4jSPN+RIzB
Wpt/3DXlFISdZd+m0k+XFlBxfJ07iGlMPJXVbpAhVYzZA0/XWDihXAz0rFE1EmpfBea1ckjPEEgn
cuBn4fnBYRHikfSXj3EPLQ6jn55wHgVrt8XXRcMQn2Ogwo0HfIHFE/Imkwgc5qTojixuGBLO2n0/
PNeufHuTQlQoErkwDsonBhobILORQ1PCBo7PETLgDnU6KIqn7hxKNwG1zXroV/C7Yd5YxsdpKzPh
uJp3Uu5tg72cbiGTWDWlkY+7mePnsj5JzsiDWoqhfPi/xDD/E43yZZcPJOWi3Qb+IdnTfo6dzju+
jxlK5GHm8HnT3K4s4PFMfi+ycWVgSIBZYD600tSJLP9/dsmozMxXV+D7fiiRtA9fP71s9Ko0TXu2
0KS1nGrPctEDSwYHGxo9Gnnwg5L2MDvaRW463pZZqSpAH1eyxLrxP/+t+HnPKNXRw3LkUAA8+J8G
Hd/8wEep0p5l8XcckdRaYWqmU9KBasgzulFfrNAVFODAZ1rx5KaVmxyTWgTsLT6pi8tBaxstlZg5
5rpZLLTliyKUWW56r8SZr8AILms+Lo/GSUlzc4z6sMWIhvLAym7tqaFoIZmFZqNNAgL9NBAYMog/
bST0KzW8o/OUsJ61+PsAbRa+QBjbQ2I1xIM7DySkQQ6BozTOuKhrg8W9yXPrebSEoLI0ZmRIylAq
hFbOilKHv2HK9lUAYSE25aJEoXIlmxlJqt4rzOVwLJmTBKHQRDOMn37qNbOrP+NGik89M5HevELB
3PfjQfZcZuvFbcZQhMsRS3wSO3NgoYJZD1J4YKmZT7ID70nKMj4hVP3xQ/cpfJexwYHcLRkpnh7Z
w4PsTTt1/HZZDMI7xP563BQnmeCGOZqqltI1Z3oY8eBtOLIA6ncRJJ6TRLETsjeqBSDME3xy2oCd
JtbyRvTBHd3fa4T03lJH1J8RHA4os87UG238ALoxlVOyya6GS1ZKuaMpxOBlnd8Qxu+BD1Ie+pCN
BK3VFuZovK1Na4HsJzJW7RU4NLxFn1a7sKsiIM8F6+gwfqKqwTxVGwDK47/V+8jmXq55X3NSx/b1
4OiR4JkLkNkFywwKh1Pyc9Tw3j2LBCcXDvoKONCPr154UMigD0zBBh3XtoUPJasPPUPiKzF3Ga4B
OQQ1jIFGRLpIWkPkxfJEeUnTj64EiDDj5AlIogmHyzobxPCddF2/Z8PDUwtHQ6BqxOABqfuaddKM
Zx+D9LVaiAQblIN8Z5CGz4cfTIMa5YbELz/uUOfiV3s/U7l2GQ1isHDfUdOLL33/RNCjwQ7idbYf
KTPkKvcG56tzqFjCmnANYWN3qg0bS+RyMQUtfYNNYOn/2yACET9wTQ9P+dPKE+mRXqyuDmUWlj17
jrU8fB4cQU8ANMS9No63BRxyVAegVaLovWHJZom/0S3eaQEQzzbDhgnbM6KTtZcjZ2ZABeZuquYM
CMiHVB8Sxe6FqOkw11aSWNud8KUFmOBKEnFY6rKaDw5SSBI51KmZyJLtO6gu83uuElS0NeuKKs6I
/5Fsu/zVS0n1X03f/9p2ObobYKpJ7aemIr/IVbhiGPceuJXBXRSw1nbd0RcXJNDnyAtKQj/cLTW3
TlFZc4m1kp6EUQ7vZhCq+zxkv6hiLdsg9Okv5UApQqwRE1cbA9D/vFBZyqYnXdVMWMZgI6L9Vs9R
k3yipTxEylBz+qhDFlcKMpVY7VWZPZt7oT4fKs6QQ3bGk6GNkPbCbSkuSuFBrjSAY3FyU4n0MTL+
nmNhbzjd99XbBKG/B9I88iEO2YNtIcJfuHK1bszRtEQOL8JCiN5r+2iZLxa3HaCNqOgYqYxo2wiJ
liEfOGfwFaE5Wt1LDhSwqNgnt6niyoasnW9EMdvg7/EBgoJIgEwPYbEETyUiEBfcvlAabolMKlaj
FMVjHv+xtIQma/rCZ7q2Bke9fD2Xw/t2q/Se117JgLS0Alf5zkq9CmpLoCttuA93LzekovbkVghG
vQRZQPMCe4vwcM9HSXVXONiuy/c/FicvgWi6Ij+FmKp85Ro9AeRXqr8tGtVR08lPVwgtVUzJu4qp
9m251mWS9p8rq9mb1vmLnqwDbd5tJOE2errdoye1dGozqezsn222dgJ4HHsMCovga3G2K5G0Rg8j
PMqgIvZz8sJP0O6/AC70cqQT5aDe22ja7PlLooE4AcW5H/Qobd/eH36HD1OTVhkxNfEZebgV1w6E
bWwAsiqMncITKpP5/Hq3ICKVeihmEJopBs7bDaS9vrM1KE0pIi2jisXsIJmYJZdjNeIpXnGsGgWY
+xj2RhFdHyINV5oNyb4gKfTa08UknjhjKBfdo63Ory4kd/s804O7Nd9hd0oAH6VknP4lAxEOBNBq
A6un7+u4yDZpzZVfNIxSP6C5Fur5ROz1sMg/fWa8cQDdYM+8kmFpQgQ3cvrCpu3DDvs6cSdgjn1u
hIars+31oH6DqMvHDKA7uxQFqwWU8/dSpU9jXg+Q2zMCqQZTviTTAOqTyNeyn1EDAmoz6gTRhHR/
t2Vugwc2y1bHO2lftG7+a+r/cHcU5J7vfh9e8buNrIHDly2z8VWDXXA/pg+oryAvJYsIKR9qv+4h
G+hp/0kkzcwccdf9Z4wXsbOFl4r5qOIszeQlbggIgtwbiX0nAsQZ2ZpKj8wBEKNGP/1sv7eUWvjh
KGyTGznRS7EJWXgEsxNtMbFaAh7GY2NnM1ukTAv0RLElt9EbazpfY4tGRIlKlr05gk9hTafCLxcJ
d/yXfzh0DwM7FMBAS/ibbbNFH6myeAZrTnfDKqIy1fDDB4mK1suATQWsqAMq9iGcVG91yIFtUdHy
EomycWNY1yJnvU2f+HsrutfvXJjztXEev7PGBZT4yvH5y/13KSsp9smEhL8dhMtHL26AN9co9iJ1
BKsRB+nEKEm0rExFnlhDIGvuckn7MvD8ZzkOIaSsd2l58zP8iA7wk7d94JFesIvyfbsT58fgLFdM
e8zNFlx0IxeH1yV8BzpniGlA8YhcM/Vcs7NxS5v6btUX+R6ZDmIGa9YnVomWTnFkZ4oRPtgZfNEO
UlbHkSz5n3NILf92FXgztWuW7I30VtUmAAH4o2mjyA91l2ZPVOCrjeIeMR29mzxs2WHDXs8hx2Iv
67c8uluSNW92u/CBul+pITLpzHTbFmx6Z2q7VhFGwNFH0AUrGrCwXGtgZR0QNST8RizKN7impbH1
+D3yVq85Oqzclip7e/NN3X9GX4Nu67qQFOFZDYt0JZjz2sYRlA4dGLm8mJgYtZX9DLXEf04D8wAB
mPTbCdujFGrnxLIg6/e5kRUfQ4PC1qslri+OURLLRWyHfy0b29UoGwwS7KWBgF7f/2CHRIGlCN6b
VI6SxqdxsJ1Cmr+21bib9XddidJ3Xj1150Ed6G7sGdvFmRjwgLUtIu4wmuEuNSibV+dQQkoARUQv
PX1s/pvuhmsCIg60ywtcJuIVYvVKLSOhnkOOmgmfSF03n/wcXexh7qTX6cuXJZv9XztGR4ikkIJd
dL6CEao4KDrUfBSaK+MLZJCRRLnhckRx32Mc0NEFlZtAga+SLrCAqQnwAccsTXzey2jhGhbQe9Se
x9PJslH8CEgpcuOJquOUDiNw9OUwap64zczWyDZitmdHdDvFoqeA1xzbA9Ha4JoZBqQ5orv2CW+Q
/6h+IIDMf6tHMYc6+DAt1ba+IfI6YR8cmV9bjiuQ7+yHQW6ND48b9kUA4rurJYeaWl4KORjkdyrc
lUf+mPf/VCqhmvB1aAnxo2snK5vGNH1YohwdIOnkCTCb21x/77dbsTVgvCN0rtecefn/a0tj3yi2
DtNYXO4szIsB4+HndvTEKbD7SXm8Xos5qlRstO3bpMCFfFINHO4Tvwxif7ibeEASCTRI8cJ9rocC
SIfpzbsVOwzy6mJUca97mQcC4b4GIzq4v/+23GcBO37kCukOOMWDtcUmR5a4P4drUUlf96bwGBc/
PAj6YlUWdujLUtZMderRJTrP8nAwCcy0pnp6kiOkbKLbRcYVh8tWpVxYinGqvFuQyiZOuh6mcI1F
JJoZXpLqHRVsmiS1X0Z69sQI1UYC2zS4Hyfy6w6KUz/uRIp8jGoBIqXscbO7jxzwpKw/m9/ZdEuR
W5Yh/hyIVGn61qoFd0uBmdvV7+wPkqdfanKDA6AR4n3mEar/3aXzcK8MzvGOE97rctaqEa1wNkF2
rPoSe3IeciFrX5zNKeea4hC2LgWn8cw6hwjbe8jocqFaPda3TR4x486AB53GTffKExAYBNNqYHKd
QGTaB31tVUIwBBoYrt/jQOOs6a20GY6COBGL3TJrjIsAH3PkjdjMi/kedyJskve1PBSwG734Fb3r
dMusiNIs3YAE+/HP3+5CVuVysvCce/qrPWkhD4hirldOoHB6RXtIFGvD/uROFwA3LlqXfzbppJLC
0+/gbz+cGddZcr9n1moRr7BnILmBy9ruzsNGJSkPm48CH484wXcV8YNTPTtOCeoESiXlTeNdcglR
xDk9HCJqtq95Xkt93fbPwlHyE7XMv2bHypPp9CR60IzB2tKBJvr5vn1DCYtwMJoy7u/kB/B11bHK
wn/UqlELTPr7jD+G1oNAOWSLE3MRhvqCefh3StthqhMMDiSYvFAlCKY4ZzpgCBwVWjfyk3EQGNgk
MhggZ+FrUMI75QnYanFKBzDbwjaLMNt6j98tD+OcDEiydIZ8yMmQpiBkj9trHx1/KM55mOGjxDj+
xfqmmFdoGHfeMwkBn/hPtJZjYUXewEVT73j8m+qtzNWcsx8PcRW3aLNw1Iacc0hXFUgSwr7nIsYg
r1uO+2pv818yuUz7VLalkTdFSHnpXfxFL5GmiLU4bHK6bY2j637XzY89ebKMw/jn/NEJNNiI2egh
e8r1ozI6q9LBR8efXadgBcXlkOfHNwe/uI/Z+mLr9/Ut3EnYJcITlehUv7XKoXVqd5wZdjrw0B1G
NqNNHKLLMELQXtGpZH2s/+kRKNCrTlTz+WEYw3G0X3FhCOUXBJzGWPNswldyaHH87G2BMDmuduKc
P8cxtyUNItXp0MdQbpGZ9Ih7+5I6Ku29sLAT7blZEh+kzs0fKivv/RQy9OVeJezISv+2TdTOeLYw
DmQhbXi6TnMMXB7X4qr1OBM3BJnnGjDGOHoyhZPg3kHLNbanKSK8b/+UM6qSQdKR+WNPOqjqzH8a
MhUOy70LHN4/ym9CoX7eStpJ3glFZwncAZURw4ApI8zIv6xTj7GTZVjJqC8QR9ObZdLRoGpHnrs5
YSEKLms8uolGVVqnud44tktdRycbn1ThXL7jGwhHiIax6EgP7HewxaJcPoMTIUE2BGa+X2OvjTR0
Y7J5ZUThRHTCZcdW8lD5kyVn2RF9MSZy9+VyPaGxWFRSXNLyHl1vyrFZW1ErxsXDfiUMCRHVR8j8
//dy5choe2wfx1RgHWwmaJmFrndNzX3W43RWjHBL/lBcSLIy584CqXUr1nbIzcgYzuJB/6l2oYoe
Gpi/rlFN77lpXEt+zgZ1nuvOdmJYdJYPjUMF0fu4SaodjvmtPi5QqQi7og23u1tI7iiKVES1EwA0
OnE248wocAjp6mzi1XL5PMwq0ozztHKtWZQyTYSVafdBYCuQsC5sZb/2AYdkeMCVc4bSb8bgO36N
JKkraG6hO4MRoUTOcaDoL5WAUturnxvzSYgyWIx/DZtjs7mSPK24saFMmzeWnXJ+S/ORW0DpvuQW
LEXXp1unbLHkY2/AgZSxkcGDHKZNBavo77vy9LZWcJO7VUjiNsyh4KBtdOVG7CGWWJyDbXva2Cai
dyUVjxgC3wr522q2Ec6bNdozZh6xlBM2Vv0aAntZcRuyuiOVg3FdkAmPDxPTdDnXMCu3dMbTprNp
Y1oxkB1BErBUiVlk8zJPUpXwtOu58h2kV/Y+WFSJJwtJ+mDw/ghvA3DXScGEbiTuus7jbv6qi/d+
0ibB8ghaHgpOOOeoJ0hMR4gu70NKI8+9iBMRBERfpUqI+hZJCtBPUpaxyFpSjZG1tsMeSTD29ON5
gsi5wTXe4evElMGiQ4qZWhxCdVJ1aMFFO0DrwdIWiXEyEq8dWctRMqS6da7WFaAgmbTz+80lEtpj
XSxoqDe+8Edrw0cS7oQSyM4IaDh/tAJH6UIY3PK2eCjgFzL69oU29aObG7k4/SzgiVWtbKxZoYCQ
vVZYvOykcJIStY9d1MqJrlGisV0HQ4Ra29LHAVgV84T8pn28tgoMCJsZorB+UPW3lvx5QIW7axy+
BoDo25eC8HUyjysMKh/jodStBLFzVYMAWpXxiWgeQkykb8JE4w2mdzP/+1D5GTFqNK1RESz1ro2I
cqpg3BIl7uqm8PkJ2JqpMx/BmjGJoz2E+K6uKOGKeG2sqr/3eQDwenJG6Ot7XoR6cL/MCPEaHp+W
HEd2GhyJOxcpaLaWGQcKLEoaD2aprEVc/38nhfv2w+TBdd27YeIUgIiL/kbsq7q04RNhBMSi7sQ4
Rofe1N62pMZC7gR1X7uuXtkQ3a2W3tfRnUcTzyqXQPJG/YFBt/g96DzX9yVecqvkRsqdwiSPm4Yz
5+/H/o7h9vBdauNZB3uQciw9Eu2EmRS3jJRcc86cA9hfpQIPp1WAgJJEh1TrSXMv5j/xtzjEtyge
kEblqvjlMitqBFF/P/aefCE1BkupNud5fOPMuWUbH27PTfckDnNu1lHuAxpejkvIUz2o0SJgBq/7
+T761BSSqcLiJ3xd4L7tWTjLDWDl04s9WwQh2nnTaIq5zrR2SzeB6Qhz5JpbPtSs8mA5YQyG6J28
JqABQZTqpgKs7EyHqfzagBzdDHESHmoDtHZ7X5pLc3peP42XXdCXMOIJkgynCu66diXyqUmZN9hw
44fnRM9n/IliOSryfqLJZ7xTTNwIwMUIBYXwNk+UeIPVE0i0Re3DSGvNrvRgFbJ6z+iUUiMvvROq
J3cr/yKtcYZvTDwcdrV0Y8NATkQrgcTsuJ7fb4sJI4cKQw9S6lrpakFGVBqyxJ4Hro2q0hJEjTrA
6QqMC4YJuj4myzaqjGo6ZZjA9lUxgVK/m630Ul/GxLVMOjSyn5p+koQZs7kON6Y+E0CSxYTw8b2W
HOlrYPPGSWq1Xwr0OKRIfMAwlVN/g928M6A8mfS6Hzs8+h+LLC5llB8my9hAnLwajxUhkHpLI/6s
DdLQHBCRkGHA+2dOJcGZDU07gPKgRXyCKbLZcU/xQdexEBxIJ+PX9V6NzQ2CegwyCLJBjJyU+YHy
9o3g6t7MbRCrZaveRZbU95gr/LRMnGccL/BhSjRE9UoPoMGTapYBLXyKfbAaBZZUK0G7Fe/FAxic
YzHziPDxdPBfcy/kkGKabQaQJgnK2lbPKYhliQZDkvqn5lDoCI+eT31sO4bq1clTuBHIFbOYUZ7C
zx3QR5g2eKTta+4W1oaO6d7KyPYZh8Phr2CdtDzsIUar2Ey9gzmCSl5rRW/Fu2Q4ZuJ/an1Wd0lW
Do76+p/R94wGfzKPDlLuWQFoJn5Y+SYGQ2n3ujgkT/cHUoGXbntkiDEUZV5u+MGYYGVrMNt/jLsz
ERwEyZLGheL6fcU3yaRc8t22gQjQUkh9J/d9AS6gUKYxMPvCon4CEKqIjsecFksFI/dDJgNQHSe8
vw6Pcuz2leYcsGrCiiq6k+YKhhUS+WRfow7cnjenUumSPQ2awdD9Nyc1kgh6nDNI5cMCn3eIeeX+
jYqIQGZKNjf9DEXA1YqBTZjQPQYC2EEoGvrho3cX9im/YU/UFTu09t/AnbQCi1PC1SrAeFrmJ4mt
8CliUu5KjXm2tcGnYl04FS2U2ImNOPRyyHOLTYXy4c8ZMKuP1MgWg4YwGaOKeCC4fPr9XocU7xdR
VvjKBH6F66JsGosm1Wepyrf4Psc41wqXeiTLt/SzqT3F5WZpMD2RNfGnbv77KA0jnceWfRpmRLTa
71T99RC6A9Q/QCKOk2o7VW8/2yxUEvHPeBxxUUPXiYhiHMgqe+n3nsAsrPZbRv0AroAel06sKnvm
UaizwkhIM8tcMEAdlLOC71LgtGhMYSdP80kbNXuBicLLtHiMq4ML22hqZKzRPHCkxZLEck0wkPUG
ZvwHGsmA6yr3LIsOmRv/QDQf72BTzV/NA3xQKhGasQIAW+vCFxxCdr3xtXYrmRdY0rkOIhRIRuWW
0xEqiUojk8qxLD3ecqJ7kcsGj4ZNVt82gIMMtSOLM3BOhMDGR2e5U31BJ8l6ZU6OQzaHkDD2fGPc
Tamp/gSfze22SgiycFazsQn5HKpIKScfb20bb4H/k60NFsDEPn/KoSmWsRtBXuFIFf8YadRlNvQI
z+QcTcsBZxfO4qx5hwYIWY9zUg5cwHktLFPde/bdLLKt/FL9cBNbVNcUvUHpoGRmQEo4oxKQD/ea
q5v0vIK4ikQCyasxcEfQCZ5zop49WnaChb2D+tH5M3Ct2obyIdRE7YrHwR5K7nRY4TWDGI5wcwdh
3+jG8tTcthlXWsMbRUxLoYg6dDxl/xE3Up1H2mpPCzkWlvEuhwNJV8KF41zDBMKPYIOP9tflpwf8
PoOHBhQwVxEY1ZqHjbZNVcl4EqB7EF3Fed8bseJcPLt8YO3XNZnc/Oh9y+VGYHDnokgNiqHu6Ety
Xk3X2Iz+58HSnGROpa1jT66QaEt+keBG3/o/D9wzvtelkkiN2IVlsAG0d0kesfw2gqr1ohxuMDEC
AK9+lYXcgbz1sZtsIfs0A4g96ieKAOWTW22o2qXDcFZh66B0Kk+WutFBXCgr/ZTaUpUYcJfOSkvE
SJtF7myH0Nx6sbLB/a6DLseY3oqJJyyXuEj1xABpdjWCYUYaGplFC63GrLi3GEL58jqJ4gj3S5lA
XW7dXF8sc5X00apry7fiZXe2IfHKN/emuyZlxa3QwIE+5UadazH4qpgACHHXdSx0jhGIXkIWgAaR
G4Xsq/ECFhrDvIQ9Ya+hQDVjLVRGYbGVfKdhfWWzma3fhfN3/ryw6txrTgzUq8LJm8NZm5KZZBHb
cQm8Rf+sesRDSKj0zauzVEvupp4aT6VE344cGSxzGGT6sgy3OdtTcGrbvKISlnrKFZB9oDqkGGAi
7Z5u0D6sXgyhpmCcOTouWVmSpBPRjyTIHfrXSXrZKfRJvukgMV7apjXraarpThdAIsO1O2R5oeh8
OIdcSxyEXIfiommO6KFRGC8dpss3/jKz8AaQiRvoDd9HJyxjPbPtHEaKTsPVcofiYBMuZNUM7/+E
kRvGHX5LgvILxOraDlnNtPyJicROASuZdRNdXVpJKuLD43iUI8rg3n3lkP+bSJU07/CsFhN3llDs
7859x6DkqHGv2JByOTgBlz/PlpoVhF+KINlDsX64fiF3P60dAJojNpiqw5Xy9B5T+SNx1b2pHLcT
sq1lXABWMDuLqyOEvfEvqGpFKVuNF1jts3+XJvAD7cbznQPATYZFDVDi06Z7+U5p6ViTEIoBlenQ
ytQ5ME3hFu8Qe4GkharNSxWcWaOG20+6Lnpyw6FBYw1NXh/BDhyAoOQXcr+iXY+5/r+KibHqMmxP
s0bxlUgkzHyxpi87WOkUsU299bXzjFUF9dyG48ZK3D7bj42lNT3CRNUrr60QxBj9YHszXlRNMWS5
8RoZc+lKdLgD2Jlc2RtsxSHDr3Cubci6GxiQCQWrLucB4UfTFBb1kjKEVt8XA+6DExfNEtGMgT/0
gjHR1EN8wG/Odtqg9uJyPiOA+IQx0kUJl5BGufU2xfDQC+mPF9awCIctLuCnXVS8bD6jSI7+GXpq
aJure9FboEZk+id+bHoygms57vj96zxaLRX5xLl0c6iXBrcWxJqJXgw6vothYnpYZSyhCvQDF0Gc
YskRLI+Q6hZgqI0pMzuHUpDttrr1s8/rKgpQf/uCl73apCRU84OETdbG19kt47GvYgqIwhx+phsV
xK9cqf8q8B6cFFy2zMNxXkiC/sQ2hHGrJcYgexFBBdB0LZWxShu6LWxRHEif5FW1YSpw82vKR8Oi
4Hecwx/1UtDyogy6TmWHDZ3cSj1GC1d6WwY1Xu6dDlUUApu9+b/XLHXTIuEPOOhJyusCjVH3afLJ
rEl/Uk2BABcedVSI4OqALIp70EFzGeiTDJUcjPCg+yk94k95TitX1OFM5Utb1qrZgDv8h2E1i5v9
Hh+D1ApYE9ew17zQhw3T+FikFOlmTNqqppkKQMO03cKBkNLFDf/qrd1PS0OJFId+w9lnxc5RymrB
c//dn42jyPLB+cQME/DhTTkoHyPrazqF4TVCUi34sFxe7iVgk9Y7qSjS4pTsHD6jcsX2pZ5cEVvb
yWF/ogQGU7X05MrGUFqjTom18lLaal40HwjUdB27g3npZ2sToPTaQkcx6r92qZ5mYuxSlY4GYQoD
4LJQNiMw4vUkueQnbQmIuRarY5G9ozmcSP3aa0E6FjeC32Ekdmrj72JYtJJDvVuWOGZgqS/MTqvI
c4S8A83qy66ebIS0A8QfdsPMraZY2Z5KZnQR1J/zTUOMw9LbkwwfgjYTmyyq0pCdNWvYu3feQhBk
Dnn0QESSZa8SH5tD/IWFM/d4h+2ELb0psxWsc6HfPvUb9wLGI8AEP6fe7ddX+ZhTs9QhFZyCy7GZ
rc/QJqB66jkqxwsUImG+NcPaQ2R7ZiXRhEIwGBwZ3m1+YFnMk1czDAzQOir3nI/iI7AAJ6MA1cTK
kBx0hlpxLSrqf9h781xzC2Xr7xU4hGF87h5ABNdRG1DSKAwaIst+BpBk/wvYE3cgWcjhXLk4eGhk
FRQ1Iz6WEp8cc8JBAIQrDFozcF9QrZBiCqcp84GFH2FtrE00rbt5mJFUsLg1gdXrY8PTVm8/jVKj
MfegJlKL5NG3FnQ+FMxz74IYJTaxp/Fpo+unMhxRVnUk3vK/zDE3kinMinRduDkvQK0EKqDG1C/0
eyZmRSsf+eUoDfCQaezCK8l/dHdsOtJ53Ze2qg2Nt84dujBDh8OZPf4kjNKWSyGWRBDOUGFJtxok
d5JLAYgkghKNKRweQRTV+IhXmZqiCVDvSkk2hv4hMrQKi+L/+gO5eYHg99LIGYpxQtrKUxm6YlT3
sh+B0LK76rnbTLqC0JboPdw1Hzem3DXWtYMgNi14M8ojIN8iWpzv/8SKLu23zjs/3c5PfEPk8LBL
ObuTuomKsS4JZ3Jl1KKm17oM17tak3LeKdfTKcP75xSKGAOO5/amu3nQhfy5AuHkZS03fvb5RrM9
Efv6voyCo1nbDYsmL13oL9MnEspFIYEtcUyNjC0xW0A7o/0DO88zM9EU/K2zGKUEOfoW6RbUbuVZ
Cv/FTMQe8qdeLmNGi2+1lJ3U6pK1n0Q+sh0tqk2VqbVGRyfwK9p+4A5bENmGlP9+M3dNs6efVfue
FY2wiWlDlW8UFJIUAk0oEhVLtwRH3kda5lcktrbEOMwA/yGULUmeVmA58MTg7iGPZImrk1mV4GQS
d2nwMbo1suFkUF6cZIUYPvDzAHg9J10TjYQlHny4b6F76f89hBTppJ3sINUOBg1uHtp6fnFN2c+9
sIdXEacSMRymixlW15aqxc6m5Z8MuNCDBOPID2IAPb7WTX2ugghgcv5DjDBp2dAn3TWHVL5JPdRf
w4CazOwF5kroJJlCN4zCEAj7kMIZqldZb8DwvKH5hYbkvTKd5lV18pLSI8R7vlBBX/DfT0cQ1kZB
G2ginVhkHbopvyBwZotsGPq4gXwAvU02fZcaYcGozhvKav+wEIR0+Xq5t3Mk/nOHbzdN0Yo3SR2G
07xnM8oB8z9dWM5tNRUiHwbw+uXhTzL2kB8y1lYTgXDwveOYJXCjsLI8DAzswjAmc3DkYpAM6QUf
RBWarxlMjCKTci1THfQV69/cGzWPLgmN5V/DEz1frG4ZM0pRUyZXkYaCwv3oFpEY21w+bjN7QR0b
Tlf1vj29roW/4qjTOZ6Lv2TK1I9d57/jESXAuC7lKbst/JbMpeb8GY9dDNMSbI/a5dkbuHifHQrM
obgnyZxKeQImDt6joiIDOt+A3eX+OaKqBSBcYO4L0/vwrNh9ohR21sXKZWLus5YLlEcDYry7ilx7
WSO6qYfoxVuR1mG2tmPn4V4ndq+tXAUmQ1Xt+NiZdYSlDfWb2pQwAUYwb3TOFkoEV2aMg+VC97Qa
/f9Rj1YeQsaGP/tYSo6wFvsYTjLgJ3Xkfyodzs2rEKnGAjmJ+1bV1hvV6S285izHfhSVtaOVS9uV
OpQX7js92GxKeMfG3yHG12u14LOBs7UXALBTD/i2ksLU5QG9PlOr4wP3l6tkJvwoFahkjW91NIg8
hgwxyJzJl9dkLICVO5tMVZYjofKlp6+pLGDAEqJbCmhtPpzmeMBmuzrbDEqiDOYOUjZcYjhMACx7
cqPoNSRbmhOASFS0TksiI2AGSJL7qTczob2n5Tiw9+Z8JfnSrQFNKCPS21Rg1M+kYweKTsLYycXZ
hrYwc43xe0hhXv/AgGfWLQjV5d/j3upklKEdiu0ce/A1ilz9CNNFOyoLSjPokuhBLwNbo85i5GL6
JorrVOnyHMlyQ9P+b46ep6b0sM9C3sD1Ie+EuQJH5mJRZhdu0vNjZcy9sUSDFbUkiVnrFgqrk4lO
Vvl4pJWbAjD99hgGpKxFdAxyuFcBmayL9V2FM/Qqbj/CMkFCb6/B6sBjI/98/gYjNTUDDPcFeaKh
crxoY8bDt7CAWr9G2bhl+x/VhOq3LTXFquBTXe7i1yWzt5ss9EFvahqaR98S4SaNDyIUYEuPvaax
g2sdU4sw2erJqtRKwpURboZiP/9TUinoZsQmCBYyBs0vqYuOjmld07lsxuuHvlEQLZPK5ItIuFFy
egs0KKmr1EVOj+gaXGewl3JoPpCrkFq+NPaLgyzSC3FztxkECtEbMSSU7h9vkqMTwgu8jTuWmsx5
MEJvBDlxpXvR+v3X5xv+9yGLX8cvDtCjdsXRRXoN61A8GjO5XqR8Qn2Pto47vjfQrQqLw8BhKdap
cCASfCihwtko4Gu+4xXNJNnbWM9l52zYD4nf/xbrK3j7p8n051jR+pqXBs0D6A8/2wmfDYTand3c
5OEgjOTSf46E9cH3Uo/RpwJcMkftML/pOMbv12kfDkB6WOJCQk8/we5eChl89bkrc3MLqTB2KpdE
xGbLK2LK4Akms1Z7/EWummblAhZLot83XIVIUaVtv/QA0NYVdCCRmMTgHkv8LVH5gbjQ294p+XPh
SxLq2KwBopSqhnKC8awgHBtNWV8RgovFhHc3hDuXGUQ6dyiibNFIblvZM+h7yvBVLKjmRMIhIi6B
1Gn2OVB5rH9Tcj7c9Xos+gzpOxx3+u1dCqnUXFBCG7a7Wa4kWclkYivw6X6vLZj8XzFRIEY79dZC
2LQmGlFzlRGUjSkodlc+IFrazpbT4YrmRuCUp3EI+d7Yj7FNCzqVhcFNgIe4ww67m0tU5iOlXo3l
QY3l9NHxRbzdVqsmvBHJZ8gJXgqbgkz//0yQjqs+Kk9iaQbd77AaYSfZkD09nJSCJmPSuQKb03O+
Yt6hKOfIRp7kzfPSq2q71tF8XSPHjH+VmlG8mnZ6BcjsNDjy4NT21DorMhLqIiO9nZorvzU4jZtj
S/gWFipAy0xQmEmFobJoa994onF1v0Sz3tvNV5nZn3kf9ECrbQVQC24GYmG2YGcZw0OHl6v78yRL
eP2halmDqATdGcG1wdLggXVN85DV5pFmkR3g4gcFxFRQDs24YLSs4bdEJDPAsaOy55tFePad7XwC
1URiTd9FMS0OdgdOO9Wp08YqSYECzZP3tOJrhW9v2K1oSyMpbWz1V0WEuEHS3rU1iTz6UXUgcvDp
nJz0yJj+HsGKckXaajNbWLpO/jxWddIg6DHFva4CeFKFGzLtGoUPXjHmVkBDi7xFgr3eUXSNUkbR
Gtg9x3a8Sq5r2QBv3epdP6/ltJJ1gkUa2hEeO4uaptTDulv4U8KKZsAzh5g8H7ZR0HFD6vlyr8c+
AOzniJ6H1Ex2ZlqCsjZti3bajVy/tlpG0TtXJpKgMBAQikJ/S5M2Op+XrLKA7ninz5gbp6iOQtTR
8q8vtV4VLxP220NbNXkSDWnMAyIFL6zn8U9W1o3gj8JE8D1BiQShKoM6TDj14HhVLWT8NtHizERL
+RrqWtenBoWmNcP3AAfcDVZhuNGHLBFx58cgiplnFCVTKpXJeqUWvfW40QIGq1M8I0wzm/fhRrvr
7xhLy2rutZIKDaKDceAySILp+h7cP37CKDDyO+dpkayozI1XQOBVzaCR6euEfVSJsPsWLBsYTofp
u+jqup4+pajX2weOFkSxjL5O7AglfBj7kQcuieKivQTRqdt7i4Qwo4vNqXOyIr4ZDD4CB+ez4l+E
x3o0GH45gsZ1t7Vee8jiu9dmCdsVcM85/cTAcUyuw1+UvF69ON5bp0nIE1h5hoXOTl9S0Ra2AtGa
QYbkOPhcttyrgUaC3SsCuvgffC0d+88ufkE6r1gvBoTCNXeFNMs4DvC2AowpFnPLhNAzCDG2LGxn
MJyTtq+8pOENmrEqiWBQfX8spXzy0r+ocDeOxpgUDxIP0VZ6Cbvj40J03Yq+t/GIz7KOuEroDHuR
7/gMH/We1zLnQH2aZoU/l7nGFsD3y5zRqqWcRC9G8/6V6VToUnR+xwd7XsOrqX3JnnrYUDSWkue4
23s3gjMAd7b2wzeviiK1nINDDNyumftUu4zL5MPCvLxIvKMc4W0I3B2eJUe+GeExj6zcwRLWxyMp
jx16AT8lYz+GWo6z9oG+mdlpLKkr8CnVOIBo3PARZpJX5cMiUXsWYfgAK3fRWdjMjA3Xk3o0RJlA
2tiJ9zf54QSTeOfaCRxKj7E8C4l4K7IHQeYa45ZTl2FHJ2DXSJMJrgIbTLpoGGX9zu1wWvXXFV1y
tzPRfAU9t8m5Y3zLv+idn6eA0CRAhLjVLcUMI//gpkqvkxyZTa2At/til0a2WkwlezlaqfbUbgmY
juKfMHEAm8UyWN76qHzE8Vl++sWVUGPDipZ3TuYcvDipXPTTbjmdpO/qWbTmKmKl4CPWPLnnyeuK
n1PUTO5ZC9uqPQ3D200RJim9R4EaVAk1QleatyPRY74uj3gPVtv/GAF8GaRS9xzMo4suHspDemvL
pAO4snHUjMi4gel6UIxI/WsK8B9WhjNYkGmOA5X2KZBf7y5b9aF3BXdZKIrQlPd0i12TkO7V0uyU
B60fwPgqh74tgTid5oVdu5k3xaCoZQ60/TDh4v3M1ZSnsv3hnAKT2FKeX6vpHt3w5iU1/OXfCrJ0
fhLWUV1rv92NgXuAJiukG0bHjERF/P0vFq++vZ9z6rsiT5vmvtO3w317p4/I5BZlhUf5ATyoUx0w
3W+WfmrE0Dw84i+C1SabEZ2NV+Gm5/tb82S4rO+BmZsbtzsh6/rgKh2udPZWm8zs5II5t+vMZw2N
A+Be+QXnHfIDJt4TR4tGNoJFFJmnCU82yoe+BNJu2Kl6bfzHSyFoChaD0i5JLD8n+pZusEEiPhs6
7jCBqdMTPvApjgp01MbjUgFVg9SkphgzYlmaRE02+7OcW9elkWBBxuopylPcaldAAoPmuJMhosBO
O7297IJYy6FJbh2o1Ho5r/iCqQ/aSgOwoGAl5cMcaBRs8GNrW3krAOR5dlx+cgTjva8AsKjfdoxC
KQLIOu7hQvnLkkNaKIKUovk0WnRKwHwS9uObMygMrFypK2FI4Y6QDhxf0XQOeTNA5S9ELA/09gez
Pa8l7k0bD72CzFdkO1ZIFv/4VxZxReTiTHfu0HQd99j8DuEh1H116zUkocaN2zr8abX4ao+pa78n
9GwOhhjIaX3+zsfLseaOX2pNBtBQQ5oTTdG1akK04fGMLRXOmsAxfa/pmAiOJjl7Gg2HnMwuNgFY
VYzBuKsr5AXDRkakCDs4f4GwZeLkp/5abns+to0W5V++yYfiKSiwTfdrUbher1OQOp+GqufYaWn5
PZBdtwmJSwwshMu8IAlg7mwGcEAHl3hqPQM+sLusaSISQnDBIf3xuoFTqBIbWOA1S2R4VTWsuSBe
hHWzTDmta13PN6Am8tYiNcD1YGds0MARzWIpVZFo5FtvqWBu7euZhWFnsn4pBxct9JleNDcKQUcr
YSf0pcLe0cOJFkGDeLExVQdxbBTKAtb3waPNR69zEvs1nRKcFYD68kV9hH3ZPqzD29Gk/csHUzED
UShOeVnxL38kYMYWfrN936P0N0bwCCxHwEukGfNL/G/W/ZBeQ64TDXstoDUoofLZ0DNJ1dlmJbbn
3PBE4fa+2XFoQf2YECHr6ZpRo9umxNXPRQbgBDFNLz+PYIuke1GKbwwit90ckD9DSuwIV0AsW5p1
W5CNm1gj9L3voIg7vJ/WVNgAVJ3EubXtlM8dWMuPo5LU5R07K/RaCEJGIWbnwoVscoxa/YlC4SVd
aAXzvA+L1KZFqz1oMa22cEktCCalAYCOEImuvffxKajp+z3WHzrxwZcCOIEHtzjioPKNRHMHY5CO
31ln/W48GhlsAEX8Yah+R7zS4I6vlZaRxI+J5ULHAh0Allja6EcjQOlwtgRpyInCNap85tvgVKnH
vuhRfSnFwmLVh61WrF1TgQHnIv17+yGGKXLfvTI97kYDOg9d4tTMJCBytLalCVUttG9V63rAqwqJ
X97lfuCsXxtFRkjmJ7I96AQ0NqbhTiddVYz1h80PEHn3HOAsWbVetULAYzCMiG7DFY0ZFF5aNNog
yA17WQh5un3O7IrcQqHpDVNQbbfmLWW/AjVnq3c6AylWnFouIKYFd4vqHQZWo9AkVqmrkw6tLi22
HaYo6seuHQ+1DEQEHNxeJ4s8UxI6XXrLjHmEvw6YKHIAxQPaGQ8fu+hrmHYeQvNIkHd2k5AOfA3a
790rfoh2Av/+VHZ8iq0aetmLa00HZxR6bb8AHxQsG6cZDwSch5lLhzsE0ROA0N+TwEb5QPNBP7m6
nQrMqL7CcOG1ZhvA8zZ4ACzZ58WouOmLRwPbnez4hqr2kl1gEs1UT3U5b4tPZmNVSAt3CI+XD/uR
DrwhE8E8Ro6EngNQXe6DtG8LnRHmbjq1usTrURJ4FJB9AOdUkq7QMFCc5+YLdQqkyPYZb5e5HZRI
V3W6FK7plNBppNoIIIxJ2ujSHRDvnDY5Fc2GLHVipby7d8C51CcZgzX7cUPbqLiEU9chxaRu7aZb
qgWzsiw2Yib8w2ihKCgPc4U5whkj3VkGnNiTfKy8bvNUDLpgAJWI0pUAc/fifPP4zfKZw6MXJazC
SiNFh6z2W1RPHGbxQ4a5INfCT3JgzIBETkSzIbCNj8xPNcjG9THgKT1GHFDE6+0hR7/kzaHDvYsC
k+y/bitTid1eSJzpK2wXSSRseGojBxpRZWMc+n/G8RL6fudhO0eoXWtCTlR5K8CeaNWBiF7kQY2w
dIVKeV2Vof8hA3zcIMeGbszYTUJ5eE10ZT04Uvgj40dZM6kO8p+D2Zdz3cMl/VtSYzFidGdc6fAw
p2IfNNdREubOUJOq1ta8UonklLqWuFAgbs7V2/4GRoitZDk3aq+EERevIk0uKwSRJAq/vzHiXMo8
ZJ/sO+2nutujHVaLpueDECHki+XnjbBwv4CU0yzuiMzwo3jk6hio5IHqN4gfzd9e4UG8y0QHdx1Q
EHXaFlGAVpoM8X1rOVEHM7eQmwgi71uXwlnNWKE3nNuocof6hLgPxBbQ5hdTFbBf7vooX2JKoiBq
uT/7ONkP8Fu4EWCQKjb109vTfLZHSPd4Pdd/+cY3Adqbrp7C3ARrlQWW/vvdHsgf9JDcqwT8z9xK
iJK0jIG7crs8cEtsNhw1QMO0wpD6bA535roFpoQhdujTJpUQpAgqmlkPDVHdy8LaWUVsjqxjk0+r
9OyujbWmltfLTm/mToYCSld0Alw25zHsNFWmDSG3KpmLUiOiJ/xbNoFnYpahK0YlbQvEfaHmCQrJ
bmYqL7NML7R9IDrHrSlwWUqkHV0uceT5tB9APjsjT+FgMES/1C0/JreWn61u94sdaoPKrzwlVcMr
v1nC3UbCA2CZ56jBhe0kxMgt9UtedHp1GwLdE+JdnC4KmEFNx5jzXiKLxCt4dCbbXJZJ4P7cq+kx
xX8mGzz+qrcWHYTu/Xe0eGLeIRztEjRkEJJzixBD9MvZS4RKOa4YLSVJWLhAyAVI/0q33iY+tfgR
GkwGmWzF0Tx9tXTZxkEe4glDzYaznCH7Baqnf8KmPtTlDVu/XVuJwy1dzF4CoZ/CNYTkaub5oYQ1
mCvpa7dQRmmkSyT+QXXFBsSfFWwKlIag17rz16XasSmg6U4V65Y2hvj6xJgHVAGPlBlQ4MxQGbqp
W5NGtfZz+lY2lYrRkgH5w73TamMx08kRnhGQiiW6XcWcBae3gh6VKazdLhsijCfThv2uBaItbhbW
5vqd61ReHvR8pGlhuEo8FgCoBqfVPsGVkOp3We9bZfnCO5bJsrQwqdkSGkifUFG3zzaM3OuvPXg/
uFi9WJZ9PITOCs7bu4Bs7Ao5oPwc3sdF4B9jht0lFCJOstDPckJ1y+xZkceRbR2V0BHW3Tmzf48q
LK9j3ZZEnctR3a6zreTrnAAcJSNd4V93Suuj7CLINCFp+IAyjBRJvsxph9i+0jXzJxFTkxHvEirH
Gh1txZ9llJJKw2ytI/T+ZifqmKLQNApFYet3gRXPpdbwo0UxrYrLMqJOL9DDrgbMbL+0S5zH9kYB
vLRfQ7YDaAixxKh9sRcSh8e5Dd9+UA/EXSX9d4JujXYeHZ029WE4b+4XsPVDSjQFgDzd1EWkardx
FRkQ+u0TQJeT7xPxdvVd1ldRX1ZY75BCTv7a4CqyPnk9xIJ+Ist1EQN3TK1byjQmx368lIDtDn6o
zNlOCO93Gvd33GdBYJRFmyg4IuAOdxrKcR5eglxyxgLCY7WW49LOjshXlO0GWBcorykv6v44AlBn
InX6nHj7ZauhAtQD6xnxbscUnVcU4wO6irI9G41yFMSc6NQbD5NtyB9Wn5HpSyzXrLMWqw4iO96H
DdjSbyqf8oBtjlyI8jeSRM61PYxWFMnyX1Jgi+s17L5VQc/OXi7KU0KMCyEtrGFwGrFaqpOFvMnD
Ln6p+eh4ajtBVR8C1s3r9bCoTvZ32F8JeH1fDEgm/Hy7GozZP9tRLKYxuxlfdmyNMGeZcJ/Y+VD0
L1NhQ2EkcsBeNP0sBMXkWrYM16GRozT4/StkeiBpAAodoj5hWz4Rqq8CQn2ftPGyVuNS13MaVBk8
Uqe07bRD+Z46VvUUPkcvgKqY3HWswFR1PsPhetW/Kh6BFVmJFMr6+sLK96HwXXXyLGKckKqRhDYB
5gKn8J9oZuO6D4HNHJX/SxiZuwiNVkNufronl25hb0vUSkW/UC+z5fI0SS/VSvL93Y716LoruQ3B
JBBWycH9qP2pLDm507YlbjJhqjIZUQKvcwFi+hnRsYeKD65SvFHqGI6Wd4yse0L1D+pTIapwkjuZ
eFxGZF64zQ4th+5CT+nfGGAeEOLZ9XH88j4KH+7Nn91wvUncuo2GkqOQ/LgaxG4e/K8SM+8wUL6a
yMH5OKByVcENChmOomrv3fRYxhAlXdZ9S9XbLvgO3OjIDLo3mrGKFlHiyLVm9zBKlrXu1B+OAKWM
Y3gVUHIVYTyh9omhJ/ngWXudSPKlZj5v4X0Az8SUTMBafHS/YX+tcSo+ZEKIjQI6APNPaoQ0AqH5
5se8pVL0LKNrYN+sRlZOlTkj6c3lXfXM+M36eGNITWV8dqunj1/LmtK3iJURYdzktXnhz1GxQmy4
iJJmjdZJ7fUcc1nUlDMiRFOIUdWhMgPASo/yM8CRYMNs5ih+EQrRtzE7wEmFdcD+2IjoTLI0EcYB
vcgWCVyp89wUd4MKgayrkRdEhzPiB5sA9qL6pEsk3gLJ1v++dyYTaOKargYHMBzepIXxQNAZd8FL
lm9Zcw3DyLxKfPYlxzWdbIj4a3J2XY+qelQs8pyZoz4DghXBMEGfHSiO6WUt45JQVKli4a1Jzk5U
zBJgro84WbJkXqNJuHc5a7/kvBFRllFxXYAPuwSt2NJpvpTMJBYZRFNWZXDUls6vvOi2KMONVSj4
BW9YGpEJOVC+zUNzJ3u3y04hXikK5GPxfvJZlfsSbSVKciH0jgRpN/ud1j101xUsbCW5ea4/fr6S
Ki9oCI4aY+UacK7cxLXs0kmFchTCn6F2i4hTNIAATv/8AgiN0996/7sbRDF6ZCZj0lw4myYEoabO
xsabyUC/6W1ld7yekxboKFe7919nHUbPcVWT7y10/1a0I02avuwCTWlpDwOpQvkxj6YuZUBIhDSA
JCh7HjPLuZEHppCUYGkpv0K6Ogv43xXKFGOR43t+seBJeO+AWyuJ8abSIJoTgkuI4vFTzfpH5AZ4
GStqA9aYRh0FF30O8ehXWp+Zu/2XqluCAFxuR4WuX7geh+RVfk8Qn+bw2ZLKMCiiogITVjwAXJcS
K8LaNGxiYLeSgjSFSOfZybcfa6D/F3bz402ajrZHLk2YJYPnRrbNlhoTg1HEJ4hqb53OVLLDYVJM
5o7cb1gtBbVDFmbAxmrkGPAZ1kIU3fcO21T/3lpkH9igmy9d8lnLIi8MsuUXeRgjJTmDJBqeTy+7
sdtPyxSu5ZW+Ky9EkrsoyKN62qrNgeTckqOv1c6LvoUx6F6O+RaCk3jLxzU5/x1FHt2wKGecsDLC
+a+4623JUwumWfVeU5ffpvrAjX39KFYDX/UWTkmX4Q6MCwnwiLe9PN1CBo4hxPb4o35PZ+nfWWR+
+aKiOUhF1fkvFET18VhbrMQ+cwtcHfGp6fRguix9V4dGdls9YYuW8UWVYQA691X2koNFxugKykqd
cHWIgIzK7yYbWcWI5J9ZaxXDR5IdEgquPhpqeGBSlfb3iXu5+4PC0NdBvytehknbQRUmF0VuqjNF
xHZDPmONlkTJP/8Jj263CJhqeZ0Iq9dsAO4AsgOmLhLShoRGEmPWfOfaclw0AixVDQfcQh8gnH48
WB3WlWRyei9xSRh38B3L6OMCSoxrGYtVEN+xwyix2Dg+u9nY3KE+7Z0WuiE67XVFbDOPNq5BrO6J
emRV40KzOJCsm43YPbqC4/SKt59MQBhJZEzPE7KQzjB/u3Y7lnBojOCXi8n13JkDvIpiIIKI50I3
6agK1C0k/GOnYy6Ax1ssGaDmy1Xp9IAz9en2ndbFUil96j/Ov4F/f34P+QvTHzy2tkZkaMznyd6R
sltImsMdOTX+b2T1lPWYK6/BX2cPK9s/nNMJ2skSgSJvF4JZWVk9LF4JKskXKWemz9mSn8vg8QjA
rmYhdwyQexNZDlfjE0fbvvpAcP4MkVdCQZx8zQcAy6F9UDn0GbKXQBQUFKNDts1oMlh/AuQ4BATQ
MHaDgIp3Z2XrBTHuWnv1pcJ9bHSTIQFbHrFX1YTfigKcnoE4Z2r0WJvl/0RtkawF6sPwPLcZzKEL
MPrWrWjJaKR6YPQ/ZgFGezA8qDgQwYWM5miMXM3+J8ANjgbxnVWYA6j3P3O2fZZBESXoMc57M14n
0xwyTR/afZ6V4q1r+vnlO/a1OSrv088YE1Wjww2Js5B4COqDovzYP0U993h9eOjF2AI1O1SHOxAe
DRVQrshmigMwAu1KrAMYE7mzBmmqC4KvwHvt0h4cRPzYHEfh2pvCu4X140mg+Zi1Cb+9ndLQObBG
jy8dUSAuA6Wr5+u3XsezAHqd/rx0H1aqf2VxJKPDcKpZ0PcVDJnYjo9RShAU2utH9SSu7CMpNzLW
nYD3uAtmBOC0x70L6ZM4cAM9W/DGIokWiu7Kk754E9q9ERmYjLDtSl4k5qecsq3M/5K5Pike0Org
gSlCmrckc3ksSjWVKkvBpUcgII05+M9ABA5hynh8j/kvwMEJoSVaoMDbsCX+k0AuWzvZb1V9OIef
351tvszvQ6egPn8t4+vio16dVpX42jIXBrnRyvg2T5M5xXy+0yirjC61wta/foFPPt87wGleolHL
Wwhnmwd0/blGZcK7M89DkUYuQIM1J9nx2ve6vn1mND2QKivggivlfWLez0IAlGjSniW0/nbTrLSB
DdkRr+Oshq/dSbkMcKOeWwc3siVbsKF/1FyakqPCeRJKV3RvSly99RRBAUDGSWcxao/HI6a78VTi
RDoZ0uh/E84+huFhHEsbpgUqpe65WHMtZ8yvFmTA+gv52hucQVr/bNUj2J0vPraKSqZ21wB1HtD8
vircoHVFeBfz1faZ2GCaJQ9Pgc+5u69mqWKUI+oU3Ts6GIvcVi9I6+GRCAi5Z3Bj2q4B20SFm0eT
QZ21WZbMvFEWg9vh6+9+gsXYfXXM4NHXEIv1Rrh+9Gpnp1u7kK7bhWN2IFeO1Cykx4xWZ9C2EQzu
idbkSr8yitrxd/TPOFifsk+PhfhZTSFxhvxdO13CNFnIrmwLinmT7BIyTAnetO9P0kiDGVrJe3w/
keLD06Dn1/mSOLpF6ww2xZoifC7CMg8eHqDc1q+256QiQWc6GDuw7bXFcLgPEGhOlSxmsX8xQJu6
oNZsBT3ROhYBLHbH8hB6QWWOs2y01YBpl994eI391rDt3YXVKx9uh/xc0rCHdzocvu7s4YQww4kn
3bJqBZkln4a0Qs4dBN0hpkcZz5gPXpW16Vn/CjcwcUiX14pSw4+CyZd28DB1mZaUoQkxxeFlaeKj
CA1oXvDLIMINurcZ2KeSp+gJg+nhiSwExMPygYHvkHbauo1vaffy3DfX26anoJe5nAEee9V0wQfD
JiCXyRoZ2s7a7Gp8Cc7PqZKqgUcJVzObNlv0KRDYH0hOVz4fwINVpktZo+/+HzIGJHbbfl/uRiOj
4OMZWKB87nv9pt6srLpEESTZr2a5PIr707HDjw/RI8XOQPBn5CZGfeCeEKiJ03d/jrqeRhvS81CR
wymODypE3ssVCx3cpNt7kbdTAbHPAXnSA5sd9SNfG5CGngFfBMywFQmRLiFwC52AhDYmt5sbDFEJ
2tksFcsXlBoJkjrMQwr4kT68nyzfRTq4Ou3QuAPJevRVFeL+jkY+2DrBOKek/LpBduAgyOyBolOP
lo+AOhorq7ST6T1BqKSNDEdmzIF5NPB76Z/w3smPne5ybtXi4G375o2pVCH7MLlzFV/S1/HeL8xE
OsEQ6mzEKwAYk9tSWlAgHEThzbORc5E4zqm1CG1Uw9ELJ0Rs1HFc7x5pw6DMPsQ4j/7MtM67JfTl
9Dm9Z6baELWaeJxShDSmvX+El1qWe3n5kJ3S0O9UiH7fHAyFpoCKTnASJfxHQIb5n2DI5OPnGYe6
q0s9AIqJDMSbFAAIw41EfjhaoeiWlPiHxeJ7m3ofW2Mv1QUaJuJgQL1ux2zr6TkUwpTnHaA5iRow
NcsugsDbeFJe5v124t5As4+U8c7dvbXHdjljWZotsIhCGArsOLYh98YQ3vnh1RRVZGoAhU21CLNG
ISjYo83+8dsgM3bJ/DVbzjPeraaBodgchtzVrJydoqs7wn83niMBAAJzWyFe+j09Nxc10iiBC3W4
j8NY7UGD4ucamVJF3CJf3Zo0b1seVT2N1Q3igG2S0+hIA8y39a1JoIajxxBteYa8dkzFH4SyahVg
gI6ta7e5AvtjrhHtWw67mmDx07+ijJFYTQUvk02u6McrAQg8zj7NzI36NNv+NgQprRvnCCLKqAFN
680zGAa8tIjpSbhJpKrysT4U3rpX8hC5Ux+VZTpjvqNiFp0bfLHq5voeRGC2O64sR7LCTrU+oJpw
CWLBAXoD2h0tsNT9g5XRViPBk6Lqe6MxcV4znsbEkCUHCiyNatl8FumHNEYU9e7wVXgrpEM8uRtW
r+npgCbDNvKAkh0GzxvWnQf0G1HcXT74Jt77cNCJljm/Qmu16GmNIqXwo+D4QnxFzg74EDoR6F1P
SB+lf6ag1W6CjEMmdxzR3Ux9dR2wgB9iVmJ06vX29YuZ21hgUXIA2feu3Q6CNQrbiKM5hT0/4jPi
ngA+UDYFuwGHx9PN/0hCzQTt0x3yMf1coo99dMLfMLWcgBYRIF3G8vGy2N690KEHxdu2V27QoGUq
Ym4b2Cz8pZZimw0XZU+u7j7ez8PhKtjhNoQg+TCkgLPMO7ai218u+d98yxv+j/gD8AFvwDKIXTIC
Q5OByGTcwQjensBerZsOIABpoyclWAAZ5bXyIdA2th3Zxxvzv0FXk6KHawiJEm1q9JZYTKYH8EnL
jzIRgi92G1JWjxhX4MW7BY7Nfb8qBW+fRlRFv3Psg2C9uVbA7bDPVU994dd/Z+R/ZNKugndjPyjE
tRdBgyh7VuNaPfj0PUScWbnkHAWZpjwEI2REebZIO6ZwD2h4UrDTdcGOhWKL57sF2UvZSjCZ+bJY
PBq3GhoSMRRLtQimlk8N8wpiFFzeLjJprmijmnB6sQLyFnZj8ZqfPJ/FlOroa8GqYOz8n7AAgbus
+TSp6MX9yksORHTc2LStLETTO4F6jXVY2CrTnQHtMWz86E4aNjAt9WKdCiyeVEm+OIbAv38mxXAC
yW/kvEe2Tq2PbDXi36zwXWXd+05Ig/ZoGyZ0g5/X8mBH7Vmsev/5xOwEv2NrsMRTW7uBleUgtPrg
1SzmYh3LJ1XAJYu5Zkqlne3bM0FpGXn/1Byy0TD40FPy5SkSn/YACyD0zxIsiz9ZxTxPH0At8BBR
WMBZn0ID3m4ieexk+rwUegAkBF/ycV8NNTHZK7CIRZRvdHFfV3slQUHdxSeeqOrzvu6Buft0BEfS
nPCl9vuT36mT7RcLnexOm1/sFR7cl/hDLiuN0tfacERaeRNZe2PdSQsNf02fizSacCsBndKSVqZs
kgKvPtbWJnpi7UyR8QewX+LrKJjULZO5QV0VdYMXF6iAQHmccDydpYc4b1tLHm1iMGjlIsBtaXJr
gb5o/zs5jBw6nPyAx6vRZZrKRL0TfMKyU3d7ucL85NxGm8gT/UxfVJgBFWFj931aaVz0uE8WPDRx
5QFZ7f+pe1hFEdOTR5d1eHsePdBPDikQTOPOhEYcNb1DY7xxtYK+jij5Rl3og/Dm+XpYHe4noblu
N6smheaVjTfPP68QBv8Bs6Et4NwuWwILWZonjwHp97BoYLfm7o0teE/txb7IcdjqfukWJ6U1EMf6
bKfqcqdp7ta5Zs06dzceglO/DSrzTrS2vW06NcnJH+FsX/5/+NxVDr1UEi807aqxBC8Ghnd7HvrJ
5INhCQ352pMGm6NedDveFpitd1jBg2sCxlsVem4Sd74F5vF4oRTGJhf3nBlBBK/DoOkHA1OYWKS3
s4kw+aQuIHs0HKPTT1m1EuQIauM0ChH3qCkutxNdeTmBOK4jFM1cgLIAAiYZ6VY8EhENlKEnGjQT
9mqRfbK5v8Ex0KBOWn7Lv8/HPX41ezTfFaKxpaoocdRyjza9oTV0GluPIjthCqqjZhtKrQ198iYA
q+3PcRuIwXxYJxl78iK/AVP3OGSTfXEMVEAzLsl/PVQ8ykNc36bq5Ntohm8AxPRJfNucXHbrRDwn
2jsoR+Kk76zMtSnp80HIuNh7X9ARz4LKtawsO/K6bGaT4uAzo8yKWK8Q08id1FMsL6DkebBBIFoP
j5COAPZUnz+lkZi9uDX7RaXKjox7LhRAUXAsGtpYvQ4FQd+qY4IwIpWRnwvJ3h1cvpyMgVDMi58h
dlOp3yNceytAZwwAHyUx+K6+vxkXD+LHMKrSks2qmFFY1Ulx6AP/0g/HG4Bx6IXqywmOyL16U6qW
H2xJqfSOfklLm13fieUM09UWhwvVHPsILUN3mLJaFRYAiY9tVxIVPKdZPK5JyoHwqamjPIbEiNac
RmJ+xvZql2/hY0Pxd7zTKSULJcH6KpYYZ0+G9ymCSbhoHmPZoxskUDWmDPtnAxG8QMgx0SUPanbl
IH7GkdFTrR6jLhFZoBeTYXbgUUiqsKCvrGrlQr6k/SVh0UvGmHOz4vxSACAhpacoXTGqYx2r4PYo
+vslJ8/6DcO8dpEfdVY8bxk74Wr6R6dGeKk0jsUkBjSAIVywJdh3d5E65QFi7Nx3PZVOt2uo3Gd6
NgJiK0Mlf5rSZNTBitRmVeAhAELdVnGNnHy77hPLmGf4pGtOnuzB+s3XiiUSlcXzjyc8uEFroUgi
diA9entrqlRmojrazuExbu3n9s+OHZ7u0N7czn9r9MMZ/aYhufjdRpZFwR8rGFQGaMXgAIJOkDyj
ZsKOLseohgqEggn5CXFEewCMb3K8zhncvO5W1f8UZpp0sfQ0A/mekaFyOfMsccNuYdffBehYBP2G
TxCN8tbr98pnKYVSDbk9J/bDBSL/yQ2V4AzwAN495MyxHjDIWRcnQ+ojd5jmNV2D+qNwvFRTuppS
2NAFOgHLoe06djl/jrSLQuflNejbCmR4IPAHWtJswyr8h9MeJ1yNJP6c2ZOsGpkNAUV5F/pfBewb
eT86GPwb760nlyud19Ye5ogW87N1m6ckcVVgI2KBUWNzy0p54GxKuwaP0k5yBGrWC28cddMX3chb
wPYhIc34i1ruAby+nYtBmBLBT+BRphaON+UD0SFJRYGKPAOYjrGF5+wf+0Z8SedsUFXPjXyb7YSe
nahK4/ykUOGtcnaDpWZEd788fhc2PdyKAhkS+rW8wmeAw9b7AZ/eXZZDYUUUo/IHE9YMEHxX7hDf
R3tK+XL+MDF5qD3U7gmLP8XbqwnDVxEb4odJq9do0MhLIuDBmIrKuzO2/Uk1qT/RfFBfcxNviqmZ
hg0kx4oJ4eefCqqnW9L923C6z3Ui/oDy0o/V2GNAVCYnYri43Mkp5VffRHpnScntXWniIfUh7xUj
SLOClEN6bxD89hv+744rRXd1waaV7xjpBta8M4I5HXmvNMXXByyFBcrLX8cM4TtmOaEN9YFCYPE8
Y3QSyNwYnGNn14+YlZBXX0FXbsbnIiHmb/LnDF5gkYNEhFuz44oTJ30zjPJWyOVFoX6MVI1HwzVj
ydZLznkm2zCF1Ex+LiBvHBYYahSI402zo6W5Q5PRcrDT4hXo5KoLrQ8mm1+TZNboGxibdzurepHI
Mf6BpMBD54MWoN349MeAmhQ9xfP1mu0s947+sINwVpbNn2HU1ihdcN7fyJk5WRR8wuJ5XAPskQm7
HCFKJEZMtXss+LvdT64xqFmuU2pI8baStDz66TMN/+Fie+Xe9bB3x4Slg7r7VsRSmUKzefRsjGNr
wkC3yFNOIXLldxZCAhhMPh8GHgK6iVshI7rPQADNJqjddDgnEq0GrFBp9B/WbQZRiukang6sYUVZ
uQHcaIdMvcjrbUxUY/hJd+ohuj1cFnel21fF6RUNksQYxfWIzkNmTGr96YP3fduiTWc9aluUpszp
uDOtbjeJ3cuA9CIFojybXEu9pxITsFweLtS328H/F86ntxjjVL5HJkdA5SR/2b6ghpo4Kgiad52p
T7b/Ddcdw9LQls9pe53DgevY8IEi9esDMcsHifqmIflkeQ3AJp9147G3AufSHn/JpXLDTPsx9HHU
uJB5+PvYZeferqBhOmO3QAKwOrSEmmIDtkVXlio0dW761BTz3MW+M/lZUXAJZ0A1eQWGroeLwvbq
8UyfTssSfBoSmXVcTuI165MSCATFBvcTk9SCIniIntPA7HT2xaKuJz5y/krXA3Teq/hE4LaP869U
Agkal0kMVXOWON3IZDxY2ZNQaKZbNIMZanuOxEPdJN5k5IS9T++fLe5/P0uYrDyeN5U8fFVRwvvB
Aln18hF7OHjQJzOmeDyEFk84uJbNebJWeJEVY+8HZamUv4hKO/9ynDE4HdbvrKFPlIl/TZCptmHd
7OYN/ziT5Rd+mM09Z/cXcC6z1RTli3wPNPo9+vZVPloqg91dFqCigAdOlmSSax6jmCJHYXadQ5J/
F94zzg1041LnkljxAEmif2YJKe3B/AJfCKwqN0cZE2VE5qd4Ip7h+FAVRoQC5LNozUs6NfMMa/gs
6DFAxTENOB6tSnO3lavBrRMFr982AEWfTeKcrWYUDnr0/A18xmQ0mGy23TG5S9jr/2kZEnuZy9O/
qFK7Qwd3+m8aFbWo5tSGF15RjI5zdRUVs5ctLIYaI9ek4j9tYxLYqN4vLTsCBweVf6uu3dvqRUm4
s17MRCXqrbtv6pRYkru1FnNv2AZTvSplglcC1h4t3FTjdxykzWtKsZzyF/Ic7xI4BiWnXuTlYpi/
QqdHl6XdBqS4vlQEAI5I1uCnFTvCo0XR3gReGQS+aR6yLf9m9qUhz/9+HO3rGGJFj0ObZZs6ZNsd
9V1e2QStGnCS+cgTrMUx8F8aCWo2OF7/ugSS9ehy/L1E7SWCT8JD5Wc5Ssu1PIDougyb5NWx+Exy
Kt1IdvwBBkgCkG/uBJnNsQHZi18yw54krn92/rQ3js0IbVC4SXXy6OFs6y+/3THOImo4cn7bp25B
inxsX/9I0QQi9rP805DByXP64gPmWHH+wSv5Mn5DcbMZFNGHOvU6dlYyq66pAPN0DMf9g2D57/8t
56MkQ/WUvjc55ni7bp6QfFCuZmXVyMOTpq+kKNHRlHnTqCHEkHttfxJ5cqSID3F4MoaKqkUhcUzV
M9xc8W5cnFPEEfIvILD460zZSHif52pRWqjpRaOsUVT+y3PabJBcg9ExZvckXmBzbO5USvPh5RS9
qKUDIEF9cb/FD0s3qXlGbVoHLyojDtJdEzai2y6p00xUKlRW9zvYFc4HwJxvV4ptcG3fn9RwrnoR
T3vr1dqtVsyfMHF1Yj4m8ENmQvseZ7gtmGpci53IMb2iWZEJ8CN8CYQPfrArnFkTFFS3pcnB8n/j
VRrY+4MivRceB7kbDKk0OgH+8LLvJlB0mmHlZIXiV2yrxM+QnN08xHKXJz3cojehDnkkCk2PaZiO
CqUJ/hyXSZuYRX5xEzoM3e9+EbDyeUD6nnGYUcIqt6EU2tIy+N+92RKGYIEQ6awX6XcTIwm68ApY
zaYGXU+WK80a63Oj+5HkBdOeqrxmY/XXcllDaty0InPICMWuc9hsDDU1dkOKrjKIfwgzWICyMkiL
eeQt09Vkzw/0ARFG+DM8P1+ztrf/6FjjdzUzJ6BjNUUSFhI3edWcWc9mS9oVSkukVLz6lu4ZEZgQ
6aXmRYeCwnymMscpAGMwBn/fMKr9CRLB6rEvEbfI4vRCCSyzczFQaN0CZsHlsChG9uFFldtbApaz
JCwn6AlYfjDFNwitcvviREoCC8veE75yqijXpUFSpFcx2o6eOTUFQJJvBl1l2gS1w1qWfaHcT32H
xrrbf0On+fStstJ3YRmufHWSxd53vH/V91htLkKJ1IE9JvnOQsyX8ewFDz5q7IPBrjFMtBx/P4r/
AckoNro1X35AbL6w8VE+fvFAr9IXs9I1lmFHP4JHKD4ZdKjD3i3KBIn8yjCnZ9i5JsnXp6tFZJ1u
8Hg53oLlVYD64bRjwreEX3sVk2RBsbOF+3EQim8Hc0b5/HW+FjC0QBqx3E+6mhVVyHxWVHsKbrWw
4pg4gFgn/nHIfwCsG6HnFe68RImSxpf6zV2zoZIof7JAMm//RhgX8O+m7Fcugrmprpk7vxziaxT9
4P7xWqiQLEWoyIB5sjfTdHs0kGwv9s5gzBaSXdwlXcENLY3jUQSgU8vQz92B31bBkUJfA97jXkfB
xQKuoK8kwUMyWEHMYPGcwikev2kNT7IZndmj5cj/j/iBpiMDnXdROvdg/u30ZK6woShcleHN9dM3
52kN1874pu0Rw+dV9Loil7IYeMbjWYgkiATsmMgfLjsADWEzzlgwY96RhT5u1qo6vgYmWV5bI26m
54LT2HXo/5erbWXnx6Ou4KGpzBxwUn3AGjR+A65Ig1pf6PwlRCgKgEtUEMxMWbqWWaF9dNilEUnl
cs+Snst/BDFe7BhOOQdwmsS6Gr1zgiDZVfk8vVtQFumXJuv7St07NXDIR5ZVAB9+bfySHJSAmvAd
HfeOZteuhUpVJeQI5Qt0ulZPFcv/XqdHPJsFNazeZY8CjkH6Ow/+C8YwF2ouAIEhDll0aqEAI7YE
N5FvidMSUIFEw+xDpSwQel8A7oDceHcMDebeeZUKbkXRjkJ0Jvva2QtkyXlPkSnmz78D9QNvaZ2+
drWyIHV/ibqNBhZH2lnXgtfDGjnIximEuNloC3wSiWmiw6R5EjGyDTF1XKYobB5WaPrewSQwDSZI
6/eiPPMwu6GfMTtxc7Ll6YvNdkCKnSIvi3JGRtRHxvS5VEpazi9RDkx7iza9HQK+1SBEkkk0F1aW
TnO21lkJoThCWOPpSGbP4fO23U68Yn9YsXl/EGDSY7eXkbUULCvxGfTj/cWOrqVZKfbDbm3e+LjO
SrQ7D6cHjWn+ZJkoI1pjaRONdLGUShbIru4O+pgfI2y5+zGgBdllTMVP18wWZZZFyGwcqbPT4eKD
GsTjoWJ9AULVjwaMPR3JMxfNFiSaAFMsBZdyz73ua1gdmeBIiKiAFM4PvP0o21DJGQN9ELdvmpUM
HN8u2PXMLfY17f0CROZrjAAkUkYf9K3pBTySF+FFMbua0XWe0rmtVVgDdk0gr0EwYHvUkmHgMjSz
KSq1GRrzLD+Zb8xHyrvlRy1hID+bCaBOgpgt0SfUjduMWJd4vWeZ4Ws2uqxhSA/hPChhNmB3X3m+
mNZYeEiooBgDwxQD8TJ4cqXny7g11518f0rWmdIKAkyaNNhoUgGkv0LV4c/csahIp+n4Xs8rIrHn
V7xyke6ndBmaGOG3XaBvSeEQAO/rrUsgqTLwlalYpMCBG5XUcABq4c3uhFWmB9SPB1JQxEyq5Rvb
J9x52g6iAvQBtHuItOxbkjcol1OluKELQpiBxhTAkS4F3dQYjspLgCOeEQ4mpsLWN8/T98rkFBbS
n+S5FpREGjccOFb5vUo5D3KjXBlIZBK6bI9UWUJNCTHIhuk2wh8EgJT145aecZg4XoKJLL+kquBI
KVObjYfWBPpaXTy+I/EUm6E2zktIsDY4xRbm3Ofx33fBhZ/Xp8GIVY6fJ4gh2qps1mxgH8SDD6Gu
Q6l3jXR5v+U8xYyG5B2HiqjYWED0prP/i2PRis2F6ISv8VlSUWHyFsqQ6PlzPm8pySe1iRkT6mgY
lNtuZB8JgEmTehhtJ6f6+LOv7Zvs759tuF7YSK3t3cP4/0XEr7BO/DaXjsp6PhrfuJPrWikvYgu8
AFG+6B7PY0MmOtKAA34g2jFqd1A0t1Q8ke5WDVTCLY22BNtiGa/lzQTzuhWZaTOsF4yYjLgGecNU
/KK4jxurCFx3WZNFK6VGbAkWAwqhlwrawWQyyZbHMF5lI92b6h5mL1cRO+ltt7aSXZ8yVjMNDrWC
/ax6+mYoIiEPM9JF7uDVDMOA6Gv42DaciZFcyoIsaU1BhmatowdSwDg+irCZZrXhwDacqnM9h6/r
mu2SAqBuYaLEuhAriyX1oXsfPsh4spHFqhAe5MhpN9CNaRL6/j6SY0J5pmuuNE9dyOQgg4nxY7Yv
IH4MO7eYdEHua63yOEcYz7v8Y/DxExH06OEUQQEaewDCdy+sik32cnMUnhc1i1EX6sgh2NGaxl/s
c1L4wh2/CylQ0cQA6A0CuXjj7qg0TcwrEk1zgEUTWNVNPwoaMQ7Q+kzkPLyDPkffGR5wlW1RCJND
maUzWAhmO/8TLvRw7wX+FoDI1ADXx04+/91bMraOrom6gjuEcJ146xPERhJjP9+yWFN7Y1BSh/8F
C2YfHzGtixAqwf38/f+JJ3S0dahyk9BA1Mrf/qLtsRn+BIgrmyLuPFUmunWimCqvjMBlKRJVJPPC
GEMeFLgaLsuPtxotxVAa5VHxulvRQ3fErLey/ajF/q1ErNzZTYTgaYNaltqldIs0k1hUJRbycudz
JJBnUHWVgR/SY6XJlLKl35p25LbZttRPV+KwFRrIVphJyt4toMPcZL+9aZqBmw9+2vE2i8jq8YKx
9T/wEpVNnn3fGymdwmxgj0CGW04Bm/BoJavRonNv5bCtKZhta2mjy7c2FBajgPrA2w/40peks7S8
ahtUVq/i75diRVov2m9D+YevpU9OMcDOzr8yVwgP6aNn2guJ30QfS3+sK1T2CxgQGA3W9b5oKYf+
/Z3r/jWXsN4HpjGDlYw6Udky0yATYt+xOUjtOjrxP/RLB51D/pNtKI/9U0HPEIdnvJGVItcuzXKU
a97Myx847nzuwNelnFJjSHuDaX2h97n4txCfIK1vuSxkwN19WBHdFe6K5jP4+r+ROp+x8eb0E4ot
1/qvuu5Axz0cNacUgbOW21XcgroXhTywNAlQutqGiIY6Y22w0hU0oBBFtpIkBOOGtpQAg3B19oK3
WlIInjkUp2V+9JqgWxtnfsEqP3twiOfZqC89M36/91PHsa5rnRJXaf4I/WcOPFp0+4pHbDPKHD83
D5yzyHlIDMnBLFGllaQjGubXK5tOBejwvRhkX0dJuqwc0eFdxPva1Zq/iIlGggh4IuUd6z845bYZ
k4tFojuJ6tvXU/HazUfgx2dNf3PGRUKGZzwSrOWOB2ooG4ov6qZUVppGrlFKilWcDjfMyBqBI+0l
B1emKMtTqkC1zk5zLoZElBSAfbQ1t7ssS5mwLyMFjEJHEvDZzY984kfMnp+eRPs3mMERVNj8KjiG
8IdTjsTeDoY7S7jR2DPLdUGyXUTSb5WZUkSEqhqj5Y84Wjd+wraQQJVPtfsLrAQs17GHV1Ckbrh2
JiHEKK3l05n+qBrQNakgXYmEZzGKhqaYYIXv8HrXdAoaVIPEL42CtNdhE+x0XUAKQzKccGdydgbY
cGtJYOVPjUUv4StJvHE132qTTDOPz2e13cV3LfEN8yTAYSk/kCMphH5iBJZFeHufQlavKJPBoFcF
ZIiB0sfis5MHg4RLqYwf81DHiKhfacdGRvOLtFT+mrSUPLhFLqEzR6wwOTnVKaN707ezpitZK8YZ
4SLTftiQkjr5eiwurpIAItQlGcWH0QbcJuqsMAColp5Xi4eqEOjlyzkCKAAVKVOdWMCC8KwoMPrr
GrCA8Gdk52NXgiNHqs4MAEGBNjXq9qDnw5HlpYRWfJYPVK+eshUqFvfKZF5LODJ79WuufVNZAFbo
GIhqEfvZ6oKBbHfbpIs5Wwuv+25uiNqkgBDU0lXPosxLm5A9iGnvsCb0KfTRJrh0z3CkCMidN/v5
yX1Mty+JsU1TMT3OB2FsRiKuR37zArOcnoIXWKThhnLKJrLYo6KFMQB/SvO1MKNEfxaFS3v+8g1v
LvztCpM9WARQyxdQ+LUuhlU7nJwumZG5kyklnlohql3b0fJ4VU4I9YCE88IDfDIq41ODEdQ5BxTa
hIbEV+20YJf/hEc74TfKJKAw5tKuhIEvE1LptcEk/glqFQYqfo2RP5JzsVw6VpJVRpE0Wobjprx4
AhCIBEZMru39JEF1xQWKfMJ7gwVBreoUkhSdJeieuesf61fRAyPnaUDR4BVytUMKYbx692MU1H9R
tNVsDyvoq5dRTLDWW431zuE39qzHOX104+5NQD/zb0YFO6S935xGxqhMr1q6zhqzatfdzJ8exkJQ
4JEpi1XeW5CfEI0haRj/b/uY5Ut8Fxns7fbL9rrOvuSKQL1yoNL4YQ2BTRHe8jCX37KNFZlOiESQ
M6meGZDYw670OfcxWKYa3xhf/UElnHE1yOOPKA7grapAe5vIYg9lOt+oSKS5ImaszE/AC++yzlao
KtDiwEWZyL6lCLTvCuc+Qq1It7jnK19VgnuVFomtOsgeV+b/CndyPnE6tAFbHg/jN3QSrTaGU7WH
qs6gj3qf5ZVa6O7ualipjGNeJFq4T9hD9h2H0h/+wvrnCrElmozlBfZ52jV6mU3HjhqbUeirFTwf
t/540/DYoi368lDF3XAh7Yc/yTT8EYhvsvvt6sqcI8xQ0db4Xpge9JDMKAT4SRzkaEIwpH/Z3i89
oeM1Ft5nAIQWkAoSr8Vu2vz60aCVDJPE2Cwkn/7B4Jvp/D5o4TEkYJOH4J7MRWnNukaqntLtQv97
YYSTjqY92wGGYfCy8tSLIiV6wyonaF83BJ+JKCSL4heUfrtLOkeSUXjUPjXin0vjoNR9UcIXNRtr
9ooU1TNec5W1onTCa21s0yIpX90lbKYc1j2KvT9Di3ChAfSOiy22L3SHDvJmel1gJuQDbwY9GI9x
9HwMQ0ozveXo0kEDsZ8443E2L02mZDg5qyjCaNIIRVbN3qfn/l2ekzMqmsgjEmrAyLOnmgxdPjjC
761EMrNEcVNZHtcV+x3hk12pGeEuGrPXMbZRt+TnRdK9GMypT71PEAzs9Pfsw6T+F2vx2HQa8ZaO
tAxWAtvl5SYpmW9dXBsWK08xwss3sZ1zZCIS2KtApieabF85uxjkXXP65ewToalUOGH2mWSj1GqQ
aU/tu67iamIv4GV0TmP+L53+l+h8Uyxc6PGRy9/eZqE0ysVHnyLLdt/FUR3O4CNn927OxIZqAu2Y
/h7eXbONrOKvGhsBGmq9S0VqLv9R15l6aOdWeis4MelRX+RFgvx/ZFGjSMtAaeVZc0GFzPQaZ9di
KljYesy2bIcthmJMP8DmkkEddS5kB9tiWJWZK74xjYC7BAwJwXEAlfJ/8hpBIxtZFCkTxs23pHsF
ishYcPW/m3OfQUaAHC7Xg9i3ko9b5Y2JXNsedcrc/libGYAbvFugikwE2BwiKS1xiGvpH7UaQbM0
YkHB40Wq6CL2Fy0HJNr9HI8GiaISuvWX/QG27iIJUdnvPudrFatQYCl5etNeF1KEYy4BQ1ZMwOZQ
bq8cEd+tgPlzw19da9YP6tLgbq6Mc3VVu6fsysj9z59XS6jtDYPh+Cm82IYN+KnLSXWv38xNhzLl
kO45zbnszv4snWGEpe1h699jn9xqiUgshTErcr5KyTkukyNOhnz8x0kDx5GjIUEvRnMw5WKoQ0BK
B9BOtrBTUQMa3zvg1lpW9vl95kOp2L0dmi9EdkRQmhHrbNpZHARQoVuTHB8uYHS7whdGqQZ99Atg
rgYAMBdXKH+EiPgHZW+XYK+Qo6tEHPOVgArOFj8gXXedoBLgRGuKzSIkQHCX2fCbWJhP8x8tMwN1
rFFwm2qizhcIFyS183OsJ6Lbe2Jds2gElavqcGIoLhURvQt7bqJ5xdnXlEDcMJ3N7+PVUuyRz5r8
KNY4NgfMjheMb4qQXMML7T8VpkG7TYpAzJU/7kIXExMja7S0qwsQ9sn2kW3kNCSLw/qEaKf0eVWu
zBIo1iHfN4bL0Fa+usUjF1xqtE4otjpPm+WjWwV1wZk5kpFIDhO7eiAr7Xtmy9EWRQkQaNMsG35j
ra9VHcKRtVZ3sC4CWz4VY6pQkAl9qxg4rLjaVYn/kHDkgfyDJBIAAR3/tESHaKpHE+EOctOWlSKJ
l/0+rGLcruxaKN94LyEjV8MH3vii4wISZnKe+8SMA/X366vgHtgAboZy31NFfgFqc5ba73zlh7Kw
w+L07p4mgEkKZDVr9Rhj8mTPN1tDhF6dZdNNADo1aNTFzFQsik9xkmwhENYVQteOkToTlXei1Vwb
uL8H0KoPguNEXC2hLDX0gjFqUdMaYOHzCQQRMT/akhmxQQXDdfdrv6LAghmpckVMrml9PhPdslIO
FDHCg2heY1wubLfgd7EEDEN0cbMjpb+OKXw/2jsLMZ2F5VOclhKdw51CqdxaDGba5Ea0S4UkGkek
OaRVwdm/oU5UxQeRqe6MAwOwDHiyLZKTpEnlcp1YzfblZSPjMEg39QzddeEVMfESf23b8uaCeKMT
o3oElzKx+Pw9rrl5UhDYARLnCjo9gf7AeT0Lr/6e+eJs7ZqcjsLENgrRiMcXRaCybt2pWC3HOqBp
fkPa2TStTuhev0qsy3lGQm1wKGQIe8FLj9rQJXWSedR7oSNU13QOuHb/abK3dWpkgIVeYDYN3V3A
gbxc0Y9TT67G6fjjkPoZeZtY8wVpGy2n6YgGdDT3vIHCxfH1CrKSr8DEF2/ztVmohc+4wyPg7JtA
gwUAaODEtj7X2X4apa1dNH5To66xPP6dAalEWNcWnJFwRbirwJAcjB6+WPXrk7bYVw8fORF4N3U8
ybdQ7UiS+j8bvlL1Fg2iAuRzQ94eCOn1IC8XY0LdAVUxnu9LtTpYAnJb6wGk4uB7XDMIBYE+Bjmr
/W8yy5P4uQFy5hKIQSR+Lt7Hw0LgIh2UfIfdQ9iexBpdheWogBAp/jYWBWdvYEzC2YRDZmoTnri9
egfFdlY4R+VLkPz8eV5EoFu0NHFwA2wy/8eMCeH4wr5gB/EyELydkDVaG4SdNXe1zbph3+IHnDB4
bVUZHyAeOWVm4+EwosGMhl9Qm3umRWomJzloG7H5EnSI4F0zDczaVu0xBQMrAQlgY5mAQF65Va5z
sANihotsC6GcICnQUT465vnFfC8QoacOMTXE1ILKemvv1+wIaNG1DjsAf1xV5dw/H46V/I/kjbtS
5VyEKD2EMzYYg/jlf1S8sIGYzauWpIlq7o2nQaVdMFVX0gfRv6K4O+rU0AbclRMyuysUuOkzGSRK
VPmOqhaxobCLNzEkK2hrU9atbCd5JPmei1W0Yw+Fk/rgBL6ULDYX6QKQiV769NaaeEzBLC6dntq2
+XVSNIgsTYh+uaBZi5+ISmavUHstrMnwvm/X3/jcGmP1z9PG28ftXKlbTSROeIAiEq0DHLOf5ReK
VOyf5kE21MudmYHitnDp1LwVMyEL2YvX8MMRkdTv0EQOLbbbgiiXsiV0OIP79Vgr53YMMoDuv9co
lQrjkQQcUe2MDXbgSuMYvUzPaW6hh5KCvURqlNt5H5bPvs6ZRAIE5A1uaUt42dwIeksgJNit+Wa4
MYu8c6OQQj9c4T4ng5czr4P/lG20KcbK2DS7ORGe0H3uw3kncvRV0+U3h+Hqbn5E0dC0vTysiZgJ
CweSSWWRD49exnoIXhy32k/FljfvOs+HAgTZP1eTNVfSZSE3xupJKxTW0Bx0bx4ALCPgPk957mY0
ILguZVtTDyP36CFpGoYrDBrEW1MbmU8v5WUi2OFi+VAiLOBWFlODLsrcwIaUjUJFfdAz2WQg7+mr
SY2N6cBI1AtiaEOZnd87JKfNkFNHPIf10n15k1Uw9sbZjpB5Cxasb1priLUaTlghXWqrclZPZ1xK
enuL3aYbIDoICyCDhWQ2W7h6rhzXzmwMa+XWFv3i/cI2KerleUXSiF2fcMOWkvs0GlNdnoNgjZ+v
S2zIQY4RoFMDkFqfz49buBNmePgCRi4CcIk5+EBLpLq77jcDasSdJ2Db5Rdhd+hz2frV8/Bi3pPO
kTAmiNwnYh+fLKeE1Aho2LwwmX8ecQhkaSPvgZxvnuXt5e9XJICZeZGIrQFLPVwGv4XNQUbMONgk
imTodDgn0sQf5uFEgatm+toPsg1Hgwblfe/CXqfzxP3qyZMFPVpH1aRTp5Qqfvym/2oz6OZUxtg0
pFaDft34EiqGkV6iD2uWHh7hfQm3dujpJIEZWMmSRPw5ANDMRK4maN+P3FaLCWnoqsLDD1H7bSXO
ZloFBpQR7iT4qjRNXvpDFT5FKMAk/Do7QwDcp6+iGnQ+5Eb8zPo1Ehbl7cYWCv761LFsBLmx6K7/
m1pNK5ESrka/OY8R/xg7gVlQOc/g1iIjjJRcQyR7zQ9wdmxuEXbW0mzBzdNI4duIK1PhcQG1B+Gj
Xr2jKAdriCjzpolb/0rPMbV6gnWHSvsvoe5JSpBYjJ4sFMTcEh/5R/3UEI7PKmU6tX0SfFrM0U0B
AL/zFeHNqEqajmHCgoiutSIVV48qctTV9vXroBZcXtuAHk5ZVfCP+7S4mshTXguD2TCjgkPT+Rnu
ybNW5COQIl4Cue1qn8QHNwhOiPK1fiq4AcWT5pHQjcxTMx3h36qLlHZpfQhoDzCtnQ2r6A3EJuOB
cB9myRZ53f2EwctkZjI0QDNZhwNkqf21vc6EPOtSSF33QIOArkU934Gg6bKi6HIDyr/4Yict/jHP
xGAt/fS/dZbra7YymmQAzwE5fVROZmL9aeLZec5FBO5VkwKbAKFzQ5JM6OVN18Ql6wp+z1RsKNKP
V41Kdddp2hsLfiQZ2MGlBZJ7hUtLpZsUmPn9PV7B2vowm5hszMkBGzM2kKNHQ6x5ONpfj81hPqbf
tz1AzEtFIxL97RQR9RKUl/1aUAvZsx2l/8YfvFstG+mQjUL84FDXIVqiTEXX95GreuXmLuATkqWJ
1X4BIo8UNoeFrCSLn4iL3JTjQB5OK1tJQ6A7fiWksu5r7BRq8+ufkGT3+I/Mvcbp0audGjME/mab
2mjmtEMsXCWFzuOWmmB+DostRGRyDIAlFM2g9GnTEcRFO/yTx7aAMvgQ1lpE5u7zp2D6ea4OEYKE
RNgFfPLzyhR81wkizUwX2oWisBKvhlvQG91XHXMyZEx7WFzgJIT93NR/veDcQ3+GWTVTMbD+GhTF
sWF3y0v5C0bQ33I2etw7Aq4OkpRTV3RphF2pBq7MrtkSA4kplLtkJZ+Djeuh9BIEGripgErNvUiL
l2pgU8psDpIKh73zggvJdl6GHblPdH7J1t+sbAB54A7DqmBpUhM2MLML7qT6AYdBdEpcFUvm+wIa
bxitrsIadMTyH53pDTknkHlBCE4E1ndMJDf1ET11G4ui0Kmj+Gq+usXJbkXo1mLcT6dZNPAcaR9O
Lr1tx7Pfz6YE9ieSedwnW5DGdTp91e5G+6niIPQkHQvNKbCdQ/qzZExEtjHCsLphnLOKBOSTXvJi
avPHMdv2SYHLuMYuucL+Sol0KtXvk/z7BVQb83F7pOifjYMaUVV97P/86D78/JxYawE5BJD5us0y
dGhoWmigO2bBmmEWdW1qz1MT68ounBYccbonVV/Fg1YcBAGu6cDj2EX+1O5wdAN+V7b8Oggs2prc
iFTIfCtpjaYj475fJhpvb4Py1UiwwsCOq/jxNaEgS7L5xEYnPiUCN2Dc1eLK9lhpbreM3RcCirJd
yKr80Nkxalq8pxkt5pdZa0+NWxI2T8hCIcLSC+WFWZHFZabmcxSldGgOirsHcbSasRmjFfr5SQqL
YTr2F55dVCe/A4+DFLroMJUtoXf/LNmCxLa37Hk//iPb7kuDTaBjfO146Dg5NgN86g+l5nlxRM6T
s0lrJ6Jb2Cu/eclJV9cS4UVQG7ouL6xY08MDF1P7fC5H6pOLCRPI9Vqwxh5FKUD/djslAC9zfxkg
3aVcbh8Af4nSlIAVumR5ArLLb9wa+UWa7povR4bzaXnob1gDDXU0+aqylC/D88KG/YkLi4gbMorr
6GGOGSTrOoCXa/Q9IvK9FSBfs9UaaB21rTbegkX6rTlNa1dXSqtTNPJ8QQs3CEqhgzX/6Y8M8uBx
a8xLX5pGGp+wVqw9PBlD4jlRIx2Zsfm8wPoctZDlax1nwXHD0vGgxjyhy7DgSekc94Q9Ro7vLWKG
j03LrM2pL+7UlAjUmGuModyVxaJ+E2TT070IL3fLisxpby5h8SrQUb9jTvntInbpiJGEOlHnhaVe
fCS4w6FlhE0NeLYTZjcAaiPjZ4eNW5WLw++jxmc0WoixTJQPUDPGE67p9/BTOtUByKNIpxlGuFAl
E3PVG6ZE8y8k9ZpzsOGt9lyQ19OI69jCCL1p0AA1+gy8jA0f6COO/TLdEaMQ+x9qD59yvZDpfLqg
xC8lRJESksEYvKLF565d3xy2JdtSp8wDLTNlBFkWmjREG8146yZpR4RwixpJOAkFuPsECgRb62k0
MLFee+AvI561IAhCorVFfe4I+Lx/v02L9lupD6Zh/loNb4hROJtAtQREOD4NILoLN+/KWJu7MiLz
1LF8soMJAEAE+QOogVpJ13jP9apr9ytkWbQi4FtZFoLvMVcHrYBtoCQ/6jxiWI1EerG6oA+eMTQq
/fgLd3PMNgNhj2bUqKejuf/VPyqorYj49M1vObYQ8aLfCGAPRBGn8JoUj/nCYIAYRAAEGoWZ5q8h
Rg5A7T3w/J6HUxmjW8CITAhdPhvgbu7zbzI/1z+6+TPPwXYZCxhRq0d9j0J4owaEcp0ysIVkDptM
1RzfzJLn3IJNLUE2ILOyRluyEd6GjFptLu7/oCyJzO5LYcNSzC3AJ2S8RH8Fk0Qw4FydHzI+xn2u
ktL14OebY+fMwe8/lKDRecO0CuE5R1sPzi6w4TPtOzbNJVo782MXluBRtr2JgExpZxDZHf+7+sYm
ueJRmR83DdeNSNk9EvMprL5oENw8+OzuXD14O2/B3g8n05sMM/AIem4qDezrgVo9Qy8bGkjz2yii
3Ph+9Ho4HKACpUZTgex4qviIkAnG/CY0tVPXJrDyvK8+1iWg2WMEbonf1E6g0PT0H09FPv3GRkh2
4dm5P3w6Wb8Wf65wan+ZQfES0oSQLkyv3hQX9LIO5XUBUWlwkDYMxjVMRw36geDs6rPvBqYnAS5L
x4SruDAtW09oftznIdQA/SIC+p8jasDN4FvkeSu/RArvVEw2X+s9Qfxge8ZlRUQDiD7zqdqD1Xn6
e6rs+Bh+07a9ohzf/4WTM21EIYOMKd/9mVsbjEKs52WLNMkKe2dnyocobIr7JF53Z5/TGnZ2pdNS
sD/LpCtl5QnFS5aRnkQWjrIgG+HFQp9zm+ZIgTklT5Fh42Ctt7TMjiBA50uGjPH0SuRnWPG2+Cbj
AAAn3zf73fX5Tp/UkdEs0sqIvGpSrJP2w1+tuY7004cPxyLgE0h5P5QngR5OEnCUuQGWMIsH9YG0
Rrka35wE7fRGlybW/AWx11Aw3jyBIeM3Yy6nu4Uy6b/RCt2Vv34C1Ml/l+9owmxoCwQrwuHouh7a
erxXbZ+0dzTb3LxQrofAbHjmBpxG5SgJmtQnDp+PmAMynWsefY4FjBQivDIKYWQqkdt9E9uSR9Qm
0P7bmE3Axq5IEYWUVgUlP3vH4N03/FMTcIk0JgN2IKODaYZEw1LSudZGPzwkRmBkoemuAiw43Q8C
oTbI1QAbDzRDB2ihMnH7JxGTgLc+gtv2r5N0J4RutnmJUBOfTmoQl1KFJNSahKzFn3WG5fcW0ftr
kZMCI6jyCftvm+SJc6Q6CkDhInJEWd90rPjMF8crOI0oG25eFRzXm3oUGaHSXPez6lmBmnQYjLed
9l9Sf2N6fzxnIDG9aRwH05eLNX4DW3PXquxkrUpqShtc4iKcuv/0WMFU/wiL6lpCZ/oX/dDGqDCk
EGtrFECOSR/6b7Mwib1dFSU63wPcO6Xk04jv7pSwZRIXrMZbkwWC6KWJAH9lnwAvsZwuZv4wIvoV
tYnvxBMna2UIJe1UGjNq3k/SOZ7MOqb6gm8/iPmD+LKvN+GJ5Gpk/miBt9CvwL/UECng7ng/Kp4D
wcfW7ATIQ7tdl+/a+AGfukBePgiiC6bFv83rsPGDGGHxFaG4EYRbtjn6xEfBdajUjASsdYdu1NbF
lq5J1Bzgwqh+ouTF45pAokYOX8nzuY9YgZSJJGMWADAaHkOi+dXZvRR/XXZ6+RGMdBK+/jvIabL5
6l0LqLpq6PvWWYwlXSZqCZjyXo3ArFnXK0h+9m7IhJWDNt0igzNfbAvS3y4DZp9Gyj9sRy+n4hCj
wXN9eyD2SLcOqKZ2oqoVbkk09Q7WieacfMkUxS74eqkmjX6Tz7CWbhmm4Zvjp9IMeqbnoJknDnnV
keaaJ8a7+3fH6jst1q3Pk959E6UckYZWD2MuZm8jRAzq7qnhSO24xjO33FqCx2RnfI8P6Dn/dTkR
YMfiNFSHZm74w5/TlP45xbcq/1nQhI6VE444YnAjsk1sod5CxYTF5plDLeeziQvG0Urnh7EEmNhI
KcIuOzf6btJqtlBw5kTFsdwxbTYu0KjnT0X9iZh0IH9ccXNbJ9F3Cty+tiLclqY2QYTE9dIcrv9s
gKZdFtZ8UagJ2iiuaBmCyT2om6YYEI4pbJvasvb2scjecZy2y5zONmV8DfYK+HIAVtxayMlDnjUH
h0KM7vHgwwOLvZZcrLD1bqDnz5dFO4oC3akiTw59qcpre3Rso29cD3UOPSMgRKCWzoH1FcnL7OTo
FC1VkK3Y+9tMSaVKWStcK08vM2Ie+y4g+LX9xvOr97vhxVFc/g7wAl67bNs9MCmOR6UbRDiug8bw
0VKtPzsTLwWxIFv5oGt+bd75VLIIgkoJHI+Z93kxgrppk1L3OPGuTnfaXtw3HahdxQtDIIAdblPu
I+q9M4YKChSRZisSAqjKoZW3G54J08m3KnCyFNn9uOIRZNPqlRULHQHWOh6yOwqXQCX5fKfy+bWK
3g2hO3O9jp8c/oj3cXrvPthYAF8oOHyQc25+HE8rFV1tw/gCJZ2MLyJObJRcp7vxvgLob9GaPJsR
bJQY7j7Ju/khjdWZ1OLuhRRUJX8zoPnZ/2BDf342D2n5TQEtlGxnI8IcY23FYm30MgszEg+rntye
e5l7hY6R1KFWRJ4CgC+yOs9ooeFN1W9+PEvXwDxkbhBC/3KEFLO6Yiy+YAowaNMD/pm5khcqu1lo
YMtfKE5qfEP5uZa2WShTdegYiCrdWmMSPXDlTxAeYABYncJdc+jWK9zS69AB8E0vRZxaVBuzw5F8
hW4A0YxAz6TqxKqMAK3SYlsuUTLaDx3rWo94Mf2FcwGJvgsPvMrnOzrruQggb/JvM9hC5hC9/+eu
tDs9L/vYlYPfJ3nL5m5cyTrijHu6tGiYe8Gik5jHDetEqLpbBeR33qeUj0Q9W83odqzyY2Wcm7ci
q1h7pDCe419d0fcEBKNfLt0IdPr5Xc4Rqc5LNWxd8QGC16G5QB7hs1XrBgh7D63IZZGaxV1ZpP52
n0fQWpaWykk/WqECUVLL3pUOCKVFdAyddXU+JtpNCln7cxdRTBnaP10fg3wS9teYT9ggcQNdWFsm
AbkfUK1z/zoGu6NdAnC1x34BC5o61ChmrT7jA8k2ktOIjRBWN90hwEgNP35mityEeHeawGZhT8wa
HePOUYzLHLlYGMbqg/WDsatBe/8K1HZogsgLBEY/eDoxKiM9G0WsAJbNpq/G0toDOSEzg1pS+aOt
E125P6/SmhpkzlHdVndFO0dRbMwxCYjlZLlYXizsZWjQOgCLi0N46VG80yFXL5/tjFHFEzeOgORD
upjq5QNEcaCtXWTfDqCqRTXHREdGPAMeFuroVe/8SR1kqwVYebQxIqCdjcES3E7h8jSI/SsWVyh1
skBOmdLb5ZVKRWnuWXOyNHYeTyVSgBnGRUiiHZQeO45djRAp0LEfw18CGEB8rU0nVywRlyuwKoUu
dMFxZRiEaikxV0v4GJTCDXX2xMFYwjQqrGYEITot8UMMd9c+hvrrzFdGYbN0f9SuvXpgelTmrFXE
h9WxFLXpSdBnfVUrEQCxpYKyCrMUyhK1TVlfv9DmuwI2HHS0TXeUQf+YdzfjnCGQeJ9XBNwmNckE
cnaaSH1TJIZqA/jZkJOteukMgOJGvdRQGO+l3e370gULgZjMVEc8BSDhTo8naFqXiPTR4jX3UnAz
3NkPFcwy/NkEsC31GAo72qv1tbFVSBz1MgcRsXKvMtj2mXNHGxWgjYSf8PncWqNV8EoezAVVqaz3
+TafUU4Av8SOKzKjsmev0G6ptk+dgCeJvcNGkCA+TY0/rqLLHoQWVs92/sRtrZ/396COcdIbyRtW
bjgbwCqzPUh2Usyj+Sk0QTandjf2WilKC1c2NjJyCKF/uXcOd7MZghWAP3PsxKgRALaxL6sgyzOP
s8vvU46SarjxaRxx55T4T/QWSi9MPE6xjHLxFHd8XlNAUvrg7glH820/ob0xvQOz3I+U9uCKWeya
KCHoWlG3xwTWkyMoF3t3dymbVeUNF0/PatXSqoDjE5rEHnHRQqQTInTvqP7LSYhaXZr4ECgwUeAl
hG0q0B0XkPTCUturi2v2VsRlSMeQJiE3FkCRKkbJE0iWl4GOo65RJoOalEYCLXR85Gm+1wWpUH+J
I58UGsxtiJ+p8kRrxozkxNLw1b9KsS+xc48zwIcDdZCLnyUCVDBuKG2KAU1CdBUSXVGqRiS1giAw
ySwcYFrjfC/JUmeiLdGqMawESKM0KrHMzzj35FwjTPti4rK60/dzytEzPrNiHlZexy+wt/UV72PS
NMh6eJ6wahVWv8KaXtaIhiY8vNRgw5AcSdiTv9GDwBKytwdIowOM+kK9sQtgE7wdkjaJuz7AlaYX
YfeR3FPwMnfNaI9s9XYgQ5Tf1HhyA8sIs+b9JjpI9fwPLFj3GjeCst2df6XKqvKNi8CFLnF2zwah
P5HfGLXuRBkR4V9JQUaK5wGTPi9nFu+Cyrwdh8CPaENiuSWmbfkGssc2eWBRpxTXOgoWmo4R/LqR
3Tzm9vm2Rp3GnmU12pu5Vsqtkbf3SeQQSStVjZvmbBw3uM6unePPMMdVdWoEBcrvL0jF24yQhhDP
UqU+Vct/iylkYyBfWQAMb39knc9W5fhDSFg6DWJZs8HeQgNQgEgVMFirPUjU9QIRUCjWZ+WjyBWu
MPdL+pt3vNu3CO7pFNz8U6ZCDnq5ksoVWgDvbx1RFFKNIBVAl8oGwEO88wClZEt2ki6uCu+iqEX6
aL+DsJJJPDbqVKX0IaaLHcqKA/KqfiIn8YCJmSKKtg14ijBQPgALFAiMwCK+v3jL0VF404DgLFT8
qIyqRmIyjlF+aL/3vPaYUZrKPVWbBCfCT7MSfOXYahALRhCjuARovYZ4LNDlTyQwJF4RiL3TqLvZ
q4vCoEivzazJbWgmrsFKGPVVhAiMPI7OqvsWfNvbvyPH/XjPyVjZDAs7BCQoGxlKfURcvA4m6atO
WGzJNeSh9m9j3D7ZRMTtMF9UTGoIrFAIHXCk/XhpGJH54TBHNLBDKMe+Qzyx3m9D4a13vpbZC8gr
TMmzz1XsSz281q3L682ROQoNq5H+Dzz85jcsDqhQwu09rrAuLC9nNUisuyM4N0mSZSK6DgVDJC2u
pKxWWDJbfvMiuUxKsDSYPCy1VPyAuLAS/qHKSLD8DZo98wvGaO2G3UBFl5J1iaiRexkIEoBPGhHO
92j8M+WIV6u8wm4Xwcq+GTAyDoiZpj37pFRNK1xvCtwDYVbXs1+43prlB62iZ/3kcur3nhRJtGfg
3f0Jz3uTRn9WyxuUnlSY8kXIEfoDT9l9s5ahoebI3JQKZ56La50vr4LRa2JCPknMon3w7Kon5CgR
mv5rgkK8b2sPRcK+9phOKDNrcewFsyOkVbAXXLEU+B7qwUCFFEESpQD9xicovlK/ypQTdEt3oy1k
v5z3MdcFfUlds+VlomKt3uomhulVDUtWpOHP8DENJMkYKBIsx5Ohd9rYjugx+btLRIq0Vb4LF4Ze
2QLjBonhvmayOr6dHTFgnOU8Kc73dMDDzjN0eDLxZ2IKsjd54mVHn3/6GmVm+OycojgugyAFN8Bq
TSUT/WoOXEsBx+mtjaShh7oHA6Wb/I8I8Y1OvgzPuscaGPWQyWHMOOiJD6HMB5Li7m4iHobkkKuJ
nQINCZ0nPWr7Dep7YmUKauxjkSMgyQSCOn6n5B7fyBprFG3DrkPH12d+3lzJc10S58sg0tRbDTgu
kg6B3Mrb4ZoW9zYV9cBt4HMF1OtXpG8kZvUVntzPqWvfEZ9WOspLnVQI3Exw5M969R5pnrKtCwyI
AbBec/We0sjizFSxlmLv4QagfTamjDaqGcMON94AX2Ckkt+eLoHYlfVmBgnsJAXtwnMMQSJTW1Ao
gjsXdfE/mlOIs06gSdDfDcqOgdVASVdy5xtjMukckIfFriWm1zesByrj3eqq23BWsjEoWqNSEk17
i9NStwKfxsnJ3FZ5ri5I1P85ItllqYSWpvpwlNB3rFm7nSSRaMDAc/X734X16Q45oF/OgR0Ap59l
5lVNa8YOm5xoHsTx/hS5EO/kRp0leTZS0ju64YjUaMwt42gdP/kfehcVAKFmBN2ztaBeQgWyYkms
UqnnXLs9qWer9ElSaZQEf/EwOj40JXtP0T98old8G9yLtAG84pY2NCh5jYPsa79E49AQ7IhHaFHm
A8Jp2kLK+dsMBQEMUnKmIEz/Gqqt0JTtb4Cno1S/u6v4uIjM7URtAM87OAwdGAtmJzpJJaLtWCCp
rk+WXM+GQPwYXIx1Kzf/nttiu+GqM6xgaUArRG2C6yy65gGRMx9sjunkMYz3GbY2gn43fjdAd8HW
C2ZTw3eIzy2zDI9rRava9YKWq7RWc1x5X6MpRI1ubiZwNPVh1I0LPtVSkrTSy3uLdIZ6MQehQOJE
YcDZmlt1J6cAC56A/cA8Ukzwb6oPb3ZwLMY17p+ZFI5nWYdUPQUwUPrt3jmf4C1Q4tVeNrI9IDnI
AEtt8/6/hIE8+WImex65xW0TyEbtWIDfP5UXFLH6uuz/R8zlFWLoFftxQy4z1TSblOMIZPAQ0M9i
tEvKjM1NHYWzGPvuMpcuZy08V+yKR23hx8Mo584JzT1TD5hsmxeWkZFMVAVPEYjeqoBb841djMYM
0XZTNYflgZlukFssLwtgQDev7v3jk3MOCCfKdwUky4YaPIkRpeRZuB0xMI5zMfhH3ycNjb31eAP+
4eO3mQdJAKosvSSuSu5PosxxqeUqShlHnnPz8S8V+HpdffSnnwvUzez99GPQkNNSo9pYTQQ9xduO
X75AsfDPyaSBQXrvT+n5zIzPEtrIkGlWsNC8DhNpq6OsQvhWZKkXt1I/Btxmxcg8HH/fb1+wH65x
x258VgcX0kPbgOr3s3RK7D3wfKKZ3Jt1v1CTso1GPLwalaz/7wnbMHseImXQNv2eQOginXAdCKYb
sugssdngxa5kYr9l3BQ9ebG9tUPYVRi/sQXoYySFH9eLPq1uQQABn8Df2GwtL+Lv4KbgRfoLQB6S
kID5W2Vz7rr4vBejlhyolhOL4V8KombY7ZGwl+apVnUGklmfYMLf0gl1VGP1897aA02URXkVxkuB
ch+pn6vNUffQ9rQWUkU8ZDigJw1ifi/dMr+E+ozmSL384uR1bzaBRhSQ/twl6H7w9SzD0spLErXc
rCpY+eiEZOugeU454IcgqEemEc0+hfTN5zrza6Q+5ddO6NkdUL6RGKiVZmRi7KbMfq7iri1k6Z3N
89ARa4aMd11IDNYBhrTNgijTnAXvVYcmRf9UNnhs7j81gMPWk5bJ4zlBszC+AnpuHCiX1UtZJp1m
A2MWeQ89DwcjTvxx2vASUWqLbx7d7RbDkbVZxFXIYpe7VOVBWjj/mGF0PY02Fn1MHddgkRSRwhrS
E5aYZ0eEd+V0YOiCFLtxpmNC8tt1VR7/zHyShB6XGXMylUds/z4uVP0yXgp2fPDlrN6KRV/uf64x
KHv5zHal8Ybqs9DBxoqgOcShOo0vBl89/yVQ0hxDmAXufMFSYLyygQ7uihZsm9YD//nP+QOJ42tz
iAneIXesAXuOGoT7rTj1aThr6j11G3Wlem7IhLX2zRXbInsAGO18sCjBN6yVbb5IgGcZ12sObLlf
+4p67tiIgf53NyU1VHYUFC9trKcbI9qyJaCupR+cqPwHJC0j5H9JWgHFe2+RFBeFPn1tTttSEXUQ
mAHySHxX6hOkwiPS6BlVc3637fNcPFYVVSMJ/Ts0B/8EmfP7NXbI31Mgd6aE9MJyNjH+YgWY7bFB
9IbP8R+7alQiELpct+TwozTioKhCxI6AgNVZtHtVNJVJyaDrhRr5KcIIzstHWmOF8Bm4H6R/tbls
c1E9Z5vc7Z01rD0l0rBhIOHPLWsXYO45/BFJMhMOYKDqhSXn70DjpHPqLb7DENtJ8FGQhAUR0ruI
efkJ2qwdzJ9UQPLpG9vap2iPEakMVuoxfnJM9wkfSa9PvWoi81jjtzFoz+th2Yq5ULiKG6zFx4VV
P0upBj+G7ogZGSUg67u0LlU1v+dMwAvrLpdPJxBGw8FLSjC6DjHoyyW+O8PwlLatfLzC7hPBwZPy
2vW/4UyGF/SaVxRPJCeOxN7mq+bK6/RJewdiCinqdlDrXyXiafp0SEZTeHjuKIbxdv99kcrDKDtv
lLw2JV7dGzETJnwoOLZLG3lsG+rfrcU0/vMijw5QnnhpIoohe34dnzFY9X5mVcKDezyjagtnNPUI
qepq6UMXiWmbiwFpK3wIv1jQ7rtZbzYD6Nx4kQc860Gf50JqQ4dbMEjHiCYHAdbsOl8EI/Zr8plV
EDZv3bxQJn9LsxPjdQp534ZOc07tAz5QOPZOtH1IXKF83RwN5x+ypIm1haiDBrj6Bo3S2Ehd/pft
vzB5JJ8u6WobNKAIYqzjIz99BQ+kKXJDf6jB4oTSe57L+hyt592KlOuVD9ilg4RXyRHX6WhwPTu2
VQWaA5dy9BehEoY5k/Vm8YkaHidT0a8VIqxa3V0VwEy/wC++eRcjUcuuilSYyzUyJ2lRfPZ0udck
xjWGgAgi8haLjEdqN5/LnNcVRQTlNY39VZIUMfifOW/pzzH0mo8Eot6yEykGrRvkfZ4DI7iLqbtn
Jp1DMnB1y70Bh0GD2uiSNemCYE1dpn6gKm+J3BByI+UgLxmLXPST5ieXnEB4Exzc2Ea48Ph18cva
lX+O02yQ1qLNh6FAhMtJv2aGXWbSXv3iby3oXwG9LXHEAZvp64HCAnutKhjv4b4+ICfBi2ZmsjFI
4yKZlmIKBJsAzisZy9l4X1JYBSVN9JELqNmS4/WxCz/odOd0p3w2fw1tDzM+x6LqaRL1kD8dDXZw
K/c4jRY9/9MvdsHRrSYmIMxZ2rdhc1aE4Uo5by+eNox1WTRs4ykYF9LbAWUyTDwXwYX76jEY1un3
HSaQAAjWws92CBhbR/tQZKDoNqrJH7rG6l7aoqJuc59Q7AC203Upa9+Pus0SbIsR9A90OybuoByC
SrMLa5xuZyM2MEyCHUsxpcfZpbRbP77PDlcrwB8PAH5AiMl0AOT+XNlSaDehTuI1BVsDT3n5aAoF
zOs7ZPpL3LS37sCO5Z0YTa+uqIf9IZWVb1hbc5HREHshIh5wIB4iEHE6h3aiAAOER4MwOE5MLf8f
cOd9LyRRXsFuK/Vm1AV6eHifcPPs90d+XfObrHd5fMTc3NraIwwL4h6lNI6B6L/NslxGWeEmpPpD
K9dRz0P3mUM6+9HWrSHIBXv2bZk78ZwZxERUENEW4Pl5HMpuep70lQXWlotuJm6lR/G/Lj5KbjDl
ISGU2yDDQ0rqSHLVO6hySyhAU8GBb1+x/F0zyijuz1aQm6IGm/zzy6+PRFLnGe4GOh0qQuPyjXmN
v2us14x5zM8vNFE1zZHvPIBFCTdQkmvcHn4vnm1imT3ypu6WkXcF1/rnzhgGBNFStyuKE8T8C4ve
YRk72rgHo4BSdNl1LqpZJwyvOxNsYnjFEsi9crF8cl/tMhE6Rkj1aV6FNMppDU1n1cXS1rB3ddTO
GPmZFJuBsdYK5nf38SR8X5HI1w11bQRwhxhUTqlqHbuEjwS2/3rjL+5SwsfMELQZaGGMgF1yu6PW
R+wkr6ekkt5SSok6l5LxGWGg7b0y4XJgJvTfGuDzBH798MOET0wX8ivgiiVQ5qq3xa4nW/vgw+mG
HoFFqnHIHOZOJAEPASzUiHavIAVuWsGiFs9Wx0xCOqKLb1F8CrC9DeJjgAvcMGHLRQ4BvBewIjk5
7TRL7kAgmiEKULMgaRy4DE8C4etgExHBTmP5423+OED49RxSdKiYhfATcz+43MzvEv/V+uk2i6xC
28A4DTIfWKXMiGTZYWKQSKrVqc9dokVhJgUdSA4kTJqK/v0mpGFCU55Jbmx21x6UolmK5GLr0etC
dBDSnSnQc8wGNgc38wVH16UxQva/awNtMBJkvJvfJaUAPH6J0vlWD3dqVI08Fmsouk8sW41a3yto
65UwbaG+7cq9n4K40NTL0Ervx4PlrM3cxPVZQR/+gm2lbumcPs7qZbKlaNNhQdvkjrwfSWXrNVEO
9JFkUMh+t2pAc5CfgUGgvxALyFLu3C/lld+YsUh6B6Y8vVlYwHqhcbW3sC1CWgAUUw9g95JcN741
9RR0aA3qY6qRDln9wDReI5trDKwmhOWH9CRCotyrfgDmc1A8lyry5APo0PpJcH0yYbyUMAzUBIef
H8HBQGmh2sAxnmBewsSccDrnKXv16xM8xzK8KFYMRhPVO4GHL1Rdzq1jpIlNRe9L18ogcpY4tpuM
5FSlq94SPvR3SHYB5gttCvAIdGfJ4arTEJTG+828Z9T+TlDwb13icLUPRB8b9Ce2yrKatj4i/Rs8
gA5HZtdlWYOvIdjqtFNAFyA8RaMEyv3+o2lT1/9GA/qcX6ZrNs3cyQUs5X0Bb3rI0caX7Mxv14Ge
1Jj03b/PSvMZOX3s6BBNWD600lJVhONF5FAR2byTEWUQ5qaom/kmrVCj1nxKtCWHwO9cQH3k/xwM
svIjL7Y6WbEjA0uG7Qm10YwfdTT17qBls6XlmjKiBxu7onoVkSIib4vtxNfpuXD7rCnqUy0jR2zV
16DNzIX6jd0f+CCVdydjdCsF/+8iM66v9j41Pbd8oEop2alQUIOLjOTOlK0susV5PN6ou6PSod5t
VANBwNGP1xx3BP6ahsX43uAO56LG6zXZAEVxVAAz6CF3NZOy3TVFQDIcWCev/tlY7ECJjnZeLAn0
/jY3SgNqFWD6pz/wR+7jBjKbYH3pej7FVJyT3OzuRpWyzkgEwDs4Dx5vEQIFmn8ee+sIByTfUznP
Rb1N1f+JLzlMOYce2mzHQOWh2AU26uIRP2POpt/SGRW3mrmHiMXrLiM0CSigcorD8tTjUeN0GnTb
hx0ifEOwkwuHSNRiZSEr/dtarAa3xG+CsKzkNX8Nu8ijO+lawyIC8DjOaDlJxB7qrA8du8WZlevz
5QCjym7XHOKiZ1r5Tai5MhRgLkzxxdJqHCyQuToBIZCwTWe3G8BDoxLbiybsumO7vtHo6JZjHcWr
dIZIWeOcfHc3G25eem+P1SqNW3+ln78HPvOtpjZwfMCphFb5bJ//cKZK6IjSRdhYRURe/EiOs0My
cYMSY1eJwfoLlSODIstcjRHEpS+vwP+kcRRqSNs9jyeHFVFYkIUu2HCjphPUgRHfOr5BRogQKrF8
i2Q49VG5yIb4yaAOKfrYLN1HivRGJuZDDe6eJowa2AX/1QSMBc7fY8a8QCWQiD+2aWD/r6XAojyo
KIuz/SXYHyTCE8BURVwMovcjGjUHc7DtPA1n5j+Dl7reLrYXKwVxFse1fjv4DU/vN69bKswil12t
oXaen8IQnKmY2wtTzsDvBi8fD7abZUVP6ycAmxd49jrjoOiAGHIgOW7QzXxdFix/YkzH7onp8jlJ
BSXbc5LCB352kZUXafsRHQYSU01zMjuurp2wbbW4TOpX8YySz3LGxfgPkpLWoePbq7T4lfqhHLVB
fE5feioYsZ9vyzzaFTHBQiGhC+5c4fiddRWbsjEa/dgNC1SuB/enbwDruPBzenO6/OrfSR8cn5+J
U3aTZIydoIN519ZXxnHOFvqKbUT/+kaJgGxIBkLR6RxHABJFlU5KdPDULBw6OfONFCbcchOK5zy5
rvcg+xrV7+RKo05NqmiCHmPOLzpdIbNpINMkIuMJBOqX9pVKWwY4V5U9+WOGRQcpPV2n/8PBniX1
lVY18M9mVLSaxiUB6FOm9Xsf42vnpOmjp7qW6kZBhmqMGU1W4X5RNvo6fkoDsL+Wui3lCHLG7yb+
I1YWcklJwbokEuWVRl8Gn4AB4UzyJvtWiSvM8fFfqEVVDQF/xPkWSEI429/SJtD/BEj+GFMRn0zs
qvCpBYUKUcx2VP/ZvzLVHlG1zkqp+qGT38ixNt3SbGx3vvHLMepM/Nmj+vfHvtjeOKZVyEoPRTnM
2YpH8ogw14sq2LwbjQtN1dRohTdUv7/vSSY7o3Hb1CjeRPH6IB+3Cj5ABSD7SmZyKGm1O6cVjwe5
NL4N+0D0obFaAKaKsMONCGB7nTbxu+9h1pGR2QQv2YSzSTRKVmU6CG+DuCo8EvN7SS5FyD3BoQDF
OUdnCJwsxPqeC3i0lmBU5+MzDY8RV3RRwOmv48i5s/3GB3PW/SoXxF6/riTtHqWM4zj+/UvvTnEp
gLYQP0wSA2ooh/9i5FEp0dW/ruOW/QH+yznQ3hRNPfJF0yrt3nyEwsRV9Pag2otF4TBz0p9TkJnI
wjrcl1TU/4nhFynug17vuV3jWfrmSq1avQDTsBE7ms5ysA0jAxCCQGGK62mA2XgOBrF9R4s2N74Z
FpJIqSMWXFCT677gLKRnv/LejC+iNQ1+IK7eqNQqRjMembGL54LgJZJggB+OXoOkJ33gK61e1DEm
RH1bv1J9+ttI+s5BMLSspd+FCVJaGTLHgDHTtnSe51a1j4NmOLOZTkwPGs/MqN1qLZRX8YoM338Z
p5lPxpJwhmbZGVd+5OvGAimdAN/Rl3G4YIc7tmCFcbT80noljxF5+E5e91wXzoc/Mkz/1JbZikwa
d4lJ8Loo32zPL41zuVNLSU8R06JaEu0470sUdF+2vppLSMBElsQbziy27ASfsIX1DkwNqegeKk5e
/Jegq0pxpZA4sU9jbBLbLmf1eCB3ska2K7AiD3jeWOzyDDbo4mNkwQGOwZzxbMniG/tVd6ON3xW1
h+eQdEHoZmGEmy/urgZHELYCmUU98gDbwovGLs2EqRTsyoH78WzXfYpnsKyatTIY5u4f+xSrLhTD
HAdY9TVyGBjkS7dMlccP9q1AQI4ZK2zr5oiGCnyU0TofqsZQKDdgW/wGV0Rh7nPJgBEzDsllEOsd
YoHbo56m1gah7ZQmw+MMOpXE0ZtPsthw7kD/nPMAhNlnwkT7KeI1jRsRWSILF3d9bHykiTkb0Wa9
qOYQ3Ztw5ZQiTWGxuFjSFaFpF/z2emd7eUw5hNxUit2CIfOvEI5s+h9i0qJ5C3A2lY+5XMUnyQge
XeWnO7UXxpyAZg9i/k13hjb2ft56D2T2vXWWzsHENuUwYtO0Ddl+uI2QgBKPwAlP5FEvk3RXKfqr
7uab3wtVsFZVEcdWiPIruufNn7Uw0zA6Fh0v9jdLA6vLG4YLfnShR8Xmw485RAS/lvNy/umbE5i+
kJi+FjCgj8BnBf5upg49740pVK8JTG9Ufn7hdEyUGrZKZ69DSoJ3/iL2Ou/D1Y38fdPBT+hVlTKd
nvBW2kw9jL2B35YWoadvfYukl0jzXQ1fiJyI4V+ngyQnk/P8kxouHCmk1Dn6yk0xMp6ivY2Iag72
D+lF1GWdBv4EFrzOaWIh93qK35g7WSytuX8h6ADGc4TzSXjtwX+xH1+w3tRJQa58A9Bc+T4Wsmkf
6aGoQgFA2OviAbrI955VZwjeLVH4i3DBhYGXLEONEoioBxFxQK/H82ojELTRmRjEN0gyVBfMrDYr
7FbD6FjsRMf4CVAKfTTV/HzE7fCJ+GedgxSZ6zOgDRyy8+QzcUw9KUUhd8JL+s0bCQIEjvtuVsAl
tiYca+Zbl15LrmEhIfg6aeQlR/ZV9BBIv1enhU9GGSUskGIB2FgXlZ+LtAkxhILr6i719QHQNAk1
dxi3wYXxaLF5el5ayY1rLI5blpjxsPB585NzF4jDKLWSQsV58WwwILetM7bwfRsLrj/v5iTFH+QL
/DdvXGVJmg2arPVUbCqMImUQoDI6qv+JHn9FKCOqfmH66xGrGJNGe6raHBRddLy3eQjVhAHOU45Q
PaKE/S0R82SwUWAlmqbMLEt8YRZquLU6J4/+0l0OSjHqU63wFeO1iDnBB2JRWrwJxXsrz+Mx506t
3ZtNmX9OcQtb4BJGx06xpEll+fZ/YmP3FQLIjd0jXOjODiJzuwz3mp25rYjVP11NT9oa0HNqfaWq
k6BvTFR2hAXM27JiKrgDCs+Te7J6xPql0Qakp5G9jr/V6pDOJ+8nu5kXBCZT8r+WeZrqAxvSfSor
+I4L56bRkE0PAxp4mdwThaWB3hYK5vEI7d9tWQrJqIygwoVtKYzLTHjLyNCl9W/jX08s0+/NIyde
lPQAZuTmbaWAtP8gAyyACGIdVQyLewpU7EsrPjoKQVKRH781Y3t/8ftgX/wrHuwJLJhOOX7qQBZF
XPvUvra+5rXZpRijrCUzDzcoQAHhspYPiMugeBQm+G1hMsloNjzM7ASHVgLyTNQZCjyjo1xwlEBD
BbzOg4V9UqYE33qTh+HhT2Mr2CO02/jLGmjzSNHNmQ7zCMzTJ4rggdYE5kMoNiA8QqR3Li3nqeZY
/98wNaC2EAoJJc55j+pPxaWb+YrfejOvK+gQ5OgkfJSrLPEKVgpfp49/0cP038Lq+vowTOG0WN6g
4dh3SNKkUnsVikFS20RiF1i/JPYMEz+GZOercpTa/SFmJNNPbSCPxFnbu5SuVfYLhS2qSIFuVOqi
5Pprh4LU5AtacBCE2LRB8BBK5IF4BOOTQgo75gbfs6I8Bx5xokc4p+lM+Vroqh4lXzk4bq2vpaAh
jVjGpWF9xjWrPLcKtpZ5sQ8Mabfke0wGkdFX+qYu9A5HqJHdJcNZnT/L/rf2c3OHJwEAsi+8F2Jd
RFlUdgXzZiafDmu4mo0FMBrR/xi/0ekiZ/+u2N7z8rx6SFVneezO1LGiTCxCUL0F4gB1RqllvwxS
YHyi1yRaSLIfOgw7kU9ZYQngKfpbQUWoA9LbvIALzBf7s30SpsxQ9CJqedUVhH9n3q04J9tcp5V5
ZFbWeR7o48FbP2B3akxrAedJx4A2bXyWrrC/QWQsEyfAQnpm/yJll6Uqua2v6xIqF3srrMEuPozp
dbg8kQz89MFXD43kM7SqGSxpKwVqhua6EcJFdY+uXPXCIaVshCo4nT/9Ql7CnIwA66Gzw4JBFD5z
B16VaNwUN6HjfRbedJS8DALwxgRhnqjUBC/V/t1shnJ3rbCMAcpwJ1q4ef0gTFQwekPWSgX6p2rZ
F3bIpDxAXLtwmX8/ib0a0OVUUz1O20OmKMSEsT4l+LqZrfTFoBCBQfP2EklNJ795CHN7x+cRUc7s
Eh62N/GIaOoxfNETnHcZk9ziemLKOx87DaIWJH7/gU+s45myJsJGoLHkT8Nq3NQgLlNOt43aYsYc
LdEge3OzuDKe8Ox/3Fg7NwkpxKaSHJOAnLPQARFpy6zSYwZTSB7VIW+3WV0zauq5qvgJydqjGhlL
szWnreGu4EV+GGo0+p714SqrKjrdb5veHmhxCfmVkjvvqGCUPdlIYnf8yeM5ModkNkJpOojiS/Z/
sMC5qaWbJvOT3dsywAj9m7Wv8KuAG2Gyl+CwTQ5yEdSejiiQXdn5RSpVLyAgQSYwSm1UtTTxXCPs
sbzHT6rWss9+cSXs3p+wuGxl0wQnZODayQxc9iAWv8q7E04jx4Qjy5i3/pBSYq/hC9STDQV0PKPj
O5h7yvF2g37/GkJtTYwyc5fipXdd4TYPYTMlW695uFWBcE/A5lRakbCR43IqwUsRLbY9K4IEV4s2
29mjDeokIxpe2MIlw3ZSLXoAn2nzbGS2oKfHxyfFTcNO3oP5FvIHGSfOSUpgFuahkXfkY0m6VMsS
4LzS+7WjvaATC0c13z1C/hbGw0kOO5Hq9KbFzYwkLs88SWPDLbX0F4fTzUwe9X6hsdOh8j9p1kMZ
L1pW4clGlfacBaanQv1TJbdaeNh82YptaZP6dEavjuu4UWnTDIfPcaEI0epm6s8DuItgCbKyrkR7
ClHUyKir4ndF7EKvAglCF07KTBNtUvHCOc96ZYY7xSA0M4gOdxFI0cZuvsB1RCfP8RNiz+qx8Him
hSi0VKC1j9mR4KKMK3+oAtverUiaLTK2+VKSFTIww4yF4G1VdS1fg15JqHLRpqMog4isBr5QIMOd
N+UdFPoQYzncH0c4yZ2GDJ6q44rw+DK7/ELArVPlqQKXumoYYouNbYLP0yvmeQwIQJVSiNtfCVZS
f9dCgKm0IqCz+1WYbeiWl2v0OLRBKT83sgWi6qoPgn+JcofPZXm4GOk5Dgv2tSZj9ucQmTn/vs1T
mRSsWKwxn5Iv/livfZoYDASyAWTCySXYzA3+PwoQPkZWzYg8OYs815byaX8v9rUW6uRDe80DxDlz
qGJ6i0f50b8a0Vs9Qf5uFDq5NcDgIM6ph4JAwdT5xALFxXICah3aVnnpdPZ3vExltaoE/0DxD2fg
k7SoV12QSkjsGB84sM/fAKi1qfG1nAj9r1X8XXSuDAgx/vbrVKzCIhTNbNVaSH0HkCFFrptMVA3F
4CKjPRwKzuOXJvcUa8Qg4f3FcgJgWDOkJ7HYZErMn36mghmbFp6taKfPWeNQp9rd82pX/4ZmG2/i
AZpG0bSeoPtH32NR5ORYUhCHOv4ogHJTa178c3wi4fXAgpRvmvKiRzqCx6kcNDhlnQij/ojFozUe
HtEA8PibDOqERO1Rc/r0kSx2hmdmHm0cgf6ntEf57YltffheBYhgQTfHoRzAIBpKmL1pRNh1VGHS
VdA2xKwEIyOszRskBeytysyVgnPbeny2w6UM3bzr48IOXlL93rIUBqf0DBLF99easeK7J/dvap/l
nCtRpc/JDfT2aWLGiXZnTRWKltZXm/nZ2OCBD/1BpIjLtmVV6v7hKc0FEO/lOK3IIw5qNeX01NlA
v0jJD/NZeqHKKxP0aI13Hz/RKQggRiesahNCi22sKRnMq+ieBlW857qdmT30gK/fH9bb/vggLtQK
JQ2H6EuDHuFgLk9QDZqkHCwfFCqOHBtAOA30uSZK4i4Q0d/9KzLHsh0bfx1EEW744cJ2ToqW/Nf/
WBF2jB7BQe9QGWYCpvjnr5h25ndYwWqt3IWh6bGnW838PsBybj6ceYmhIA8YRTvK3F+uE3KrHMAz
g9CpZovYimci/7UUQjq5G1ZKRC8w+1IGNXZeghWAQwmdTothUeObnmSWgyp2ZJaJKC5sj5Ev5p9d
608mxjDGgZKEO1ESZkRJoHC7LyIZhBBZclvBJX6YMk3hsTioarbcJMR7srmi87zYjsF9Xbs09STZ
9GuSeRjs2Huh8NbV+RQZ8evTw+2WfwhRpzOsPjUMhEgL8vFzXgWHZiDoSKQpEUMXL/uztarVcp96
Ba1kSJWQH7z0aHHIgN2JL/5MKGXX/2+udTrWyJpScDw86QIfp1nt9IIL6Mp3b824AONG+TnW86+i
hPmDLDbcyl9nLfaf+aqe8FsrUzl4zkqXEKyyn+dx0N8YiYUpED3aeKDGZpNfc67/UpyRoSjsfOkr
T/srOZXI9jAA5Azgx5kY5cx2M1RJgiEZSLblVH/UD/vrI/rZAtc9mIAWDoMZqg7uSHSczFijH6Oc
SHd9fRWNevO+WNra3a7XW1vPOZZMXLltqh2SgOKSQUANTdw24koSMdLJKCqvSobyG3raCZnT1oaf
sdZJO+IVc0vMwrmJL38ouF8Q7GKcSHG/jKYoddECGmk0kLghzkwU0goyNPxw7kt4Mt4s60cH3xkt
kqza5+TNxj8Yv+DwcpGeCRw5Nwr7BRLWLZedF8JJaOWV1HLnpbf1Sj5xFgSPFdL/ddYpK5wbFOo7
J6Et6G+5RrL2CUcAr07P0/ufev5CiFYTIsL0EDrsCQX6RRDt4RTCc3xtnaD15WTkBE9J1KxoxSZ1
ShAjmRYutqlAhuwxKANtA7Q5/lb2MS43vAJWVs0e7z++37x7VNHp/ErYD//KgVnXwzP/FGQETC1O
tO6oDdZF/tQzU3nh/LlyXUL/5zD1Of5Qgc60sESDzR1sc/p1i0gaSCCRRekU4N4IIrf4UzLlKno4
WC014FhjA7oX6kd4ftK2mNJrJIJFSx3/c2/QKSxf1Xtnu/zxtokiyGWRZoXoSeltrvSShe0IBHFa
WxYBTjs02cFtz9veKJkKWnjhGVJEZqRKVowlOegaZ1isN15A1HW5Cs+eXcRo9haK3u0fKy+efdTH
M1mNLa6x5IqXpiTmdq77oPDsrqUB3pCwJeRlVQHWY/bMIphZJXjnywUFORl6BIQEPT+MOXmcLBxT
1Sv4OngssOrIjIC9crQRW3fThz7XuVQEOLi+4MV2SQxzITuG+GRmQ+1+x7xdHJF3bidyVLLffalz
Myb5f4T0ja3RCtKYlYTN/cNH+aX6l/u7K9M/IZAov8HL6opgGJk05t2tkoVqqZCb63h2ng2qLMsN
Jkm2B1vxfzZgKscYXvRzDlIaDJCyoTeL+j2QKXkqdxHW1omaHYP1xRUNd6ScKu8+Y5lEYvpkSsva
0dRGecyrusSoaEKbNABID053ixSl9M1FgCCK0Tr98ecY15euh1EFE8qYjychtgJxvMUe89A1ttAd
DRLhfcmTXYMM+JWoZ+bYqGV6PPu49g1VmAPHyAskGEE0iQCxHXbm26uZE79qzECtqge/KmKA1Tcs
jUa/rt7IeiGRVcoY7g8Wz0FfPwf09iTudIpTGNYTby25RveOlfF9CaJjn5Gxnkhae3N8ar2bNoff
Z94pn04Ig62opLkqBEgs+esqOCRVmXfYVvql3hu64U6bnQIyND20+wVrqfjk51NXnnfZ+oVY2Qm+
VLphm/bUKhGGdoky9WkUc32glM/FUnbLnZKh4tMfwYVvQu6mqt8fvh02xt5HHOPxZroimUlEtEf8
RwYOzR1oVwpyFH1JxvfVuVY9HolTDYwGQDposrhBmb5940BlpcvlmBd3SNt/ep92wTYt9naovx+u
vJbGyUdPuICuXBPz4s3MWQ8Wp9DC9ohPCcKwaWhBrgP3gKInQT4end5MlZOI3miQZc47AXaNKP0W
htvS/567rsY1fYakBNuWJfNYPt922Suxq8wkoxprzfgk/j8og1RaVtz/dAJcvv55QffcTG7TbGSi
k6X0QOJDbhUgZwNXKMx/8SaEFPo5VrAIauA/+LGBS8yRxpoqt6kd+WWCTUVLoDRNsdO55rASAEqJ
6or5yLNMC8r6KK0O8N9Lj8DT3tCa6SLSZUvoAiINKVb6tQLLtvQRSEKlJP29QxnGKULgDcR3F8Gc
UFOaNiVdQ3homVQ278J8bDV55v7DeDd6nku/q7M/M7cOQfgD7M5Fy6F6lWqYoqxGnQICdODFCPg+
Rx3uWcYwxYILp0cfvwXCVqcjCKi9RutwhGFSRU0bymPLfPeZrAbAHLcibtHvOZeQN7oY04GddM7v
lr2E0RfTueVWBQs/+s1y+a96tjLGAoRzQ0amTiWKtgkRHR5HbAsBLBUoxHSnABoc5/HJqHibReLU
3QzVMO5CDbDCBPfdCexrkjNkJn/zI86eN5NP8swEQIliDSTuiZc9c/uutHAr42tGT/neUbUOlMyD
W1xYZCms2Yw4JzcZl8qFw8M+B49tYLMSTiNtWy1PAyW9IE0ryyaKDhtZsUso8fNymy1v2HbHcVAt
dj3rBOs/qQP9CyLq33LPrVqAvTEJjNrPgelTn0ldyuphbONj6GCdJ+doAY+4A9Ri+Xq7Lm7i6xFf
MKOvTnziTYqJ3+3MWS6LD6ckoRqSPKSGVWyvf21htax6deUDNur5lPvfFPmgIU+yn60dBJ33sIV6
nCh+/M9kUFFbt6dIjZU3Mr6KeguC/Ivq2n+n3YbnxWq2e6GSo2QncL6079DBeuDeO2UbosUC+znq
0o5A4LiUuJhAKdLTdU5ALFjNR5NAG9dUfDETJgnIvgPlfQI9r1LZ3kDzPA8xwLzY020oeVnLwWJy
/1hVav98IBgwnSfBV33n5X1CYpXvT7lv/aDQi+g9RtO4qD2BIcNYSI18La7vQB5bgKF0FOY9HTU3
FiUWm+gLN6foYBErY0RWaCZ5oDQwMzEUaynRejDsoxWBBWLyBSLH3nLeZ3FBHwqs1o3YoTuXMkPK
1rBthVeqxJQG+U7amB4mw0xiuXC5NxZ3Jx9YoCcHWxvxKNYZVQoLJELmHXcM5pdkCLmd8ZwC/shB
b7dzVEz1Y6BX0YNYO5uGSzhCaPjDI3+9ufG6Opc6c9j2OSjnx9eJYtWi4b2jJWlqBJV0AT5oSEhy
HWD4/CiNdQ8I54xkE5COsRLjR1ffY0/8pr8gpOIaeXp+Hz4zf3s6ggg+p0T0/ubk3QszwR/LbP7Y
YEaCnoE13pkRV7x+dQ9Fpp1ZGZ2HuqYkJtKyuyvLSVRdav1m/m4fCRPxsqtC6qLHbKkLaiPVl6/9
o4vcArDE4WWyvYUEFDuSvM3MvphiBYMq2+pasEWsPfRr06/kFCae2W1t/Nthg+TW7XtF+H6lQt2R
NNhqsrwwM9AzIL8piVH0hJ+d/ZNfhsO4+MpsOYq6e80Al2gpx8J3Tb6PAIt/S5JkFjDLik+27TTJ
dYSXEbaD/3L/l/qyIrPXS/8agilW3vAXyKEwuwQzDf5BwmM/BCNCH1bc469cVYI3UdBiEOD9u6F1
tPgcwtdoSAQn+53DQaNKPwFhs8B9oQi6RDF5P6YgVSat8+wuQmqOuBwE9zgBSvHtLK1ovaAux0nF
QTM0/YgcP98yo7MWA0YM0ytgFolt2oMRgxsTlYvUasUbNHAqTjO0k//R0yGEMbnKUoEOJqlFd550
32Dvf32+eFYj4/vrazhlu84VpdJP3Ou/dXahBs3HGu1FZIdMxBeMHO9Jj1jMevqY1fLbkBdFEkgo
NBxXsOUyd0AHCgws/T5ZngGnR1ymzDSOJiCkWadEnMryg9eIb1lzt23wVHXKrtvQpO1pNwaDF+PC
Mw7uDypBW0EUrBUl7fRB6mpdMb1klQv0EeF6QZzILalLhKZzMKloIlmzLKJMZgaGlbAtDvLDrBkc
lDH9yGl35vdmB9zC2aJ8lj2UWSxxv5YreNYsGxa37VVa9olMIVQ7lLEAm9L5f3PPQ2/B37DFBP4O
5VvudBMCBTT5YI2yompDshYuqj0mghtSc9OodDxojT7PRX1wSowGvbbgfYzYVFbDYR46hlgFNyok
HOK40FduWT8Rr4BOsTtWJoqDO2DovSIZ0YrZIrYv7ySOYaIHmiTlySaj9zMGfZTFT2+PF0Hl/ZBg
5wZ5BWLf5LgWtzDPRp7SmaKrfRDZJbGge/kL5lb2C4TZGTuolxdDbrwFBG1IX4f82JRUo+aK0Bm1
v8v2ox3Z6kbgrjtQhU9chQCvvvyblUYVueak9iICwztuspIkh/D7er4YN3boYodmGEo7kAdvQV5B
aGGRcsUedOUxmrVctEKpoI6Pky73MxpLisS520cAJDN7o9YbDNuWuB0lA0MFMkL/ZtPTiMaTNxfO
BzoGqiZ/G8vrq69dJmZJ+XIUDpTkUpsRBTuZDa6H7aePaH5ZfiUNc/1Rrh9I3/ODfu3ZJGOyveKE
iAvhiEbj7BPHW+S5KQ2/ti+cgR88uz+3YuF1NQvrxDXpnm08sudFRhflQVJbxybaIoOIJ4bBHO+F
6h3rtTJlI13WIaIzqliAFDaTFwM7ryjlvlDySgy/DVvvTkEy03twgw/ebJ3ImdXAeXMTHfhXsHe8
jbbvtl+v76WV2bOzoqDc5vP+sGZPsvfzrqvk4/K9xNU04iSW354fhqh8+jpEAymuEzRxQy0an1tP
Eu9bBmU/lVPDipdpN/K3Q+ZuK8gGchE41s6rLxUzd5suc56GahLV6nT1yrHFXBpbSocjdWKvCqBj
fh7PmWKoTE85dw3jzXJFJbBVIoZ6GGbd+wHexU1nbJPkELkl0O8ecLjk8LxiMllsKN5UK9zIkSKe
1VVnrF+UR1Jz7u25+AjD6nrj5B2qfbTtDKJB4N5xot34SWj7OijED+vwS/cH9JIhkj2Kv4Jqbnlt
ydoYRNwaUHrkWf0yM4QubrDsDyyYcj+m0GXkd8C+F98WdTtgLXVx55nJkA72ARkSAYpWI85I+/13
V8l/S+YUJUS8y3cUslQ6l2tKIUlEnLha/sX3IJSYB5qIoekn0iZyEi/Gz7eAQ1mJwNKeGnuhYqZv
ecvp7VLL5uKzwQGYKbYIlW3enSbhB5hrGHGHkPWKvvkAL2vC9v+kued36Ot4voBKnm2QsPnT+DP9
LwHxXi6wpz92r1xsL6iPlN0LHN7ZHNZY3kAVFUlvz7Rqn858z/h8CDHjXb3HnEo4BuGqxsTPfMuE
6JuSkhKJrYNgDtpMg76v+F9WBpVoRw2sFOPwRk1/nv9euYqiCiZYxAqDn3UF1i82bitDZBMvnXVO
W+pWsOC5iNPPi/UCGv3w6Vl7xFt3MeTnWCh6e5f9NTz30mIW5sumKWcFUaMbGlZEOQOvCyKMCfYW
UHASAkymKeWq86HDDsjNGgH2pjG3xNLLi/FpXq/YL951yjvQcIkJ8nDknM+nFwRUOR7h3Dd39rjZ
R0Hr1NbCTQZEXEY7J4OC45sg12xdqsXA6ydvvXgnv2OrI3sSNmjxjKs6Sm3WgfFfPustX+WtlEwZ
hCW4F9JpLpzqh7bYWp0IA5UX9YFxiXMsxzplRHhGIHh0M7/IMeOCh2mg8pRPUexU+agwxRrmEKiS
ZrJFq1fmsglsPhf/F4229COWFFhhdSQoy+1LvL3XJBKdPbKC4JlgVmKbyIdoweskXyMeRxpAUJTJ
doGqjZXf6/KmNkMrF75xTx79Zk1a2NWQMZaJHwX1+rjw26VpGtpquqZgnhscrFJX0Sg1msyI8/vm
n/eybUDV2Pqcl2ACxq36ibOyJ5JLoOfCISiskFmGdjqiu+B29B+H/zyUZ9UGR2/Y4le3ey16o4hu
OBWHQrP1zK2bKeghC/BQTmtE1JBzi6UFy6V5To7Jbjbw+tZ7hrlYFxDvAPBBcJR1p1baccJzmLDu
7xyDQ28MIQ7DUprNMQnUaJNveXOaMB/Lci3FUsWNh7+ZYLh7DcvCqwM56AsEcqYjnjWBIFeo86LX
JfeKZJ2GuDdF6yjTi+gNTy5WPJUrMmcubG0DkzcNZcwYfG6U+QwEjlP0xn9dkaQDPuCi8WpkB9hd
FPLABmhy8vE0dCe/lQSSe6zcDz3T2RkuJOtEwoydah/mYhZUz2c4Qh6RnZQIZG729O7o1qQH6COf
1rGs+zb/9mrMsBgRVe55hRlFrm4RT43v6NU7Cw3HFq3JewtKWQcLB7iztliLne8I6XjGsZU8KwgZ
cxicY5qHTS4QFb0OzeDvYY94UwEK0KzvaBu1YR1vjku3atpRxMkKpQslGGBhJXGbsBwORoot/6v8
v7Um+8W7wSXb6BYV+qB+4PtYEGoFHiEyK4SIaiqCktL20+w92I+dkz7lnZy4Sk6nzPqoTBd4Lt71
tJT+N8lpzrPRNFvLbRYGyvWYyotnA2zTf3tDu3CIqFd7zSyqqultNJDERDEIu64cgCVsQ1BNgZxa
sAO1hnFVgHs2ceABa0bmdIlGKYxOlIkgV66Ih54IgVlpx72Uh1tQH92ZKOV+Ekz8PBCVmwIV0ilz
kc33rvBembP9CkHXY/coPyRdRK40w3tD3hlxXJlzh0rRVpT6ppyqLffVMGOmBSEn2YaJpBCeN9sX
nHo4ioy36PSM5B+iUaAGn3LEBVYkgJ5Mr/PzS4wlaKpmR2l5sCauidrX1E575Wa7jKA32t6wwT2J
GtR3IgXOpq76wTz0vq/SKJ6Z9SqnZYr/wBJXM93utYRE9yL6BabB2p3K1jjafOPRY1omjqH8NwF1
egoZTb21kwUk0bk2sW6HUxWPlVBlR6azZBA1pe8PFbQEK1tf82vy6zJJeqG+bR6ui0XeQsBxsFSp
6QeVbi+8hJxMuFDbBxTiYwEqEkBJzFdfuBsC7WsNHGjKhnzDS7w7GgEPoVZVFjOiRac3zGTSzt/c
+Fg3eSOywauNER5nyrfW3a5SPfcfRsGtL7xeIPrPnc93h2MqcUte8byWXJYQvYqGvGSuHm2qWk4o
uS8UXLUyzg5OLGVcB+7FEqcwhRQ+6U09BcKnCkio6/pQcfGscLodcHUUsLCMGoW1k1EYGzShYaSE
aY2ksV/LjajkyWiuPjrkgxXWmUX72+i1lRgh6Ll38pS0/6gjvcIWT4bsdjD+0Llmdn1XnLHOo7Ol
p8j67+G6CmJ05JG4qRNappOOEIKCLrnCd2McXOX6ybND2hI1BGthBm8x94cA2YjaCJ9eSoEA4aKz
EctM2hkQF6bq41cvQAQoEDCREq7LdkAmgqE1+zADLdmtVU/yKPIqXRwDuAi3lGaR0W+Bjx/CMJPs
r3TzVX40vnLN4OQ+NT1NC/b7ZfBNOpgbvu6OWsBxeQ9jXVicN9Z8MiDIBqeMdsb2N/PO74D+T/vR
xhEaE5tCzbrU+cdJIdNPZiK+mwT6HEhIS3qhJhWehK2ZXCgpnQKwdu3amhXtYmUQL6vNIfW1yC13
p6Z9IjaNyn0SosNA53Apvdft4Xg4lss0ZAQzwYMZTLfIvR9IHylkSKQWGIL7eJr3k9ftwlvfc8vN
pL1EYZxx9c+MdIDWZuYDU4/67WOx10DcYVHdnko1zJmkfbFIo0WqJdd0ETy6zKKMvk4MfY4HlXo5
LjtB+TtKXXYUqjv5Bwf5Wh0AqQGJ9nC0hdBewPW6J1HT1xPxqEs6Iez4Uy483hcLtP6zA2o/NV3g
SS18L7AYWUrqXRNomHZ7NwUIZwpYone1J1DSH1TRYDWNVJ3FsKhhG/bqoapTV/Y9HrGXee2vFIQE
ZiDXyFOIDMhX8GQjzQfApz3+yeyYEHrSrQrItfnIf6ZsfFgIBKO2QN9FyC2AWwU7hM+ppndO8EDz
cbAMAIM0lVviZs1C/wXFf74c07CSJ5YbaMT0GCDFStus4DyaMDWR8032xTPIe8Ks/1BUAiBWf13e
iun9w/NFNKGshpfwIbbm2DKeILUnyMLeDFg4TTmXQ6wDYfrVQRhRAZIU2/jT8CV5Lq63G3rRmrAk
k2pNwgSRtIX5Hnm6nV6izoHv5fXwpLZBc3mLdnbwKgZVH+a47uWzxBr+nvxXHa4AXpV655voqovP
9rTsX5EuCSsr/ICCxtr77+Ysjkr9nPbaOIF2USoEdZ3y8/4zP0R6H5Ckk6uvuX2WOKbUJCqnZLxq
B9Q4SsTqKkwkGTUmQM62FhTggwShdyV6GfLtLHIGF6lbLR8a9ye0JveLiaWiAbkqCEGRp57CvAng
q9Id0Ip/K0mHUYd750eEo0Vj5MGIKVtpYL5jTO0QNGXUEUemNEBydAKTe5bPuIotm+eHn6i/E5AQ
dBlkd+dYGF3S81xe0D5Pa90vLDL/xSv7NlYh9mAexbvVMJ2wjCgbd86nnpRbtDOKVox8ft5lSurK
fZ5ZheZNr5GuqSSnRvEYc9t06nKax7YqceJ/Hro9JaaG/vk1n6hZkOp+S9NHZxt1c3j/l6i4bSRh
chYuw+6FgKcoQopcLoQJjCQPkopZItolhq0ml8IgXKzAaPFn94WHd+Dk2zez+ecxuOa4Xgxbt86n
g2y1iNW+IxCT3yjoS3Y3E8ma418bKCxARf82e4uoz5od+oWyBwVmQA+xIEumqh10/AZgkuqetdev
7mTjkFOTa59y3ccDa0ILqc3OoluEl5tXPxTQ0VzWBpODYZPfy7qY8Udz6JINhr/pfcoUi5hmoPI5
Rw6MVm/x7Oafym+ONcrtHkim5gf9JVUB6dAH9EPILSCy3TiJphg7Yjp9hW9MGFIatTazjY0K8xOl
VnTHESx+6RJRxSd3tNj4gnoPDPMmwP4Vzxst1jqNkwEOCRNyWILXuUJ1VBo4VsWiKj9EmyD8GKtT
1aLJXwg28toa0rdLj7VKRkZEjq774oqbiib8JxfALSA5gu1VrjWJmULV12osuuYhTORnrnoFKnsO
Y1uu4HTgTpxCAyNKPz5fEzBUG7aw49fm+PpyIQ5wAjdLwXvP22Qd2blz+Aixo5bD0zz7EjalY4p2
4f5e5d6oLQLabMpSshja588C4Vn5Epq1SuF7jFmLM76kf8+EpAe2bzdvAxS8hNnl0r9VliEayB4L
7Io2ZSp6B5bNmUM9RDtlMjXZCZMge6GvO2X4faHJaM1WwehRbdX5OprJZ/HwOlYjC0W8Y+pekF8K
FmK7p6Zy5T3gdNTkUmfdyMs8LYSBmETTOJ1PIBYDHQ7bYme8mcW97dEgms7n+I8ZYxiH/R1xhqp1
pV/gFRrjDHDbgP2J036rBjPnBQi26KDIBSnQXrTo70Oe2K1UZzraDF1YXEfC5fmoWw2d/nkbVTwH
A6uF1SGhA6brmjEBDNZu56xhHYv/eCrgg7mnM1VccM4bDswud8zEiCty8n1QaKrYorNAvXZZVJeQ
hNv0bqRpxmSpWpbLTbNc/7D+S8hHuyWYb+9PQuwXUxOIbPy2EQ/sbbRVaSpkNvVOUN9+2JBIWXel
tDAPfaonn62O9qNYkWznAEX5+e3kNZr/u7kM+KV6YK9oRa+3rkpfBTblPQs2plE8orPRgG+Q7gyB
QSBwZ+V48VjcATYCkur8oNIrUgrHyCDu4t+S6J69piVYe81UMdkVXezH8BX6BKLFTBE2UOChXl96
f0rmaMlrnGXDWAm9yJOAB4GciqrDtA/fYJMk7+c/c0UK8lfx+cIMI9Xw6K7/0k+WYCKquPjRU5pU
uiAU81zikNIdrv8gatCLHoF4RoZaLc/ed7RyXscM7i2gUVxrm1g/PuVSrbq6GeWEUt+lBTTINU4e
3/KzFRMUK/jPcJ9p/n/wR5VzKv2WTpHjlusAf/UjSL6vB2SkiiO9NTyl/nqq6Ky7McF0sjlf8dkn
0aKWaASpT6Yotadtqr7utJugSmxXtnbxlzqfXXK1QR8wxJGluGlUATOrRG/TzLc6pv0H+oBmA9/B
ER2jxWd8t1kZR0Bc+lE+L76HGaUyfkWXpjtjt/RFMIgZBZgItjv6Hnh7qUPFh686nkEz9HhTH8Ih
gHG0DLVKyS+RyzGMYjSM+mjQUT29FusshzJ7+z3dZS9vrNDQqMY9ZO25coPF+4bYMxuB3/hzGAwz
a0VYQD9MLKALQBw9mCYMBNz/KQWVYPaL9h30cGZ832VzmTFmVjtP4WOq9rEB6nNK3c7fk0z7Y68a
C1R/dm/c+c6erPa7CbgPE4ftZJEB5dgrQ3EbP2JirX39n22pay/3zRdNgtuEVIlqEZyuO5kNYFwm
iP2bdpC99cUa0xZwtuvZQhp9Mye8hbBNerZOQT8DWgLqAgbpMft2/IlUk7KIlvk5J5Pyh5GPYRoI
CGV35Txc/4tArBnjfEzNIPFubEGHYMBfLxHgFowDa2tH6MNFhYAoiH5Ui4zdnUWTv9QLcTzlp+it
UT/gAFIeKj4Ym0lgbCqHLKekLH4E8nPi7QEoCnZcjtTMDxm+0ijEG+gdt72naCNuJ30XQBVCsomv
kpagp//uTeDsiEYMsbg6Hs2R0Ljv/95CF15ZJ+pAjExqkxipry27wcj6dKs/pn6Puh2ovnXtOj0A
SRDWCS2qMYBXz9UQI6WUg9tYi/JEQ2+amd9zLjdd3fF9ARN8ZHA8Avu5717nqKHDtYVrvv8edZ/P
Nq2mRuP4SJUHT4Ci+OEzTM0bZy6tRgcVGZnGNd4vrN8FzzYjk2oU8KdXkosyXg2ajGLB8YE5r+Qk
GYHpAaqAUrLLYdfye1BRjYUqoDXma7tbmNyn6qRm6aTxp3c15gCVP6Th4tIPJ7Lj08msjpUC6Emr
5Ttm3r82ZOWDfilFe5g2nM89Dw85hNtBKVllgH5mJziTkbpno6sjDE1MoqbUrLoAoOQ4aPs36GkG
sfUCAddlLd6CqW45usuyhprGlfX+ZBk10LUqOnNTpznhrGAbJZx5gJ+nRDMEQFNVSuQEtz6vPGq2
wTUdnI9/zXtPYkXJaI4FLo6iKyMCuj6grxnLwdOZdvibMi27XptyHvtXKnJC2MrUuQfw0vuLTOak
srarK9kaJcfjzLxAhBbAgbhYrv3jQGJcqwshbexJVTip9ZxpyOc8dALgk+JgE+Cxiq5Bb4a2lwG9
eEPROjXUNJz+OzebKib0b1vbEZGjRQUciFzq50MaB61M4CKz+yXaKhLAjSEvx1oCTOznbiv5wcCK
8L07L/Byjlj/p8gLCoyesp26aud8klcdfqjfGydWgUVXjFShUr7XpFqi2ELZMefSJzW0GRejDWO0
ewwtloTlW79JvsV7jIB329yhM/0TNxmD4ozKDmG8Gq1MiB52hp+KHX3Y5wZKtMBa7MXlbUwB+1Mq
1lPgWDHbgmgNSbC/be0wOyAnIdo68zZ6cdtQddSKFc1Ybyw8FLpZCi+0LC3TjzM/3lYA3xhIe+2Y
kqx1ahedKkeqq3iy1zLVdEHzVwT+spvsSGWONgiF3Pu06jCT6ziLNun+q9OMt2Vrwf0jffvkgJU7
AXUP7rBDwNt/Vfn9mH5t1xdFDWhCOoU6Ot86ZoqaSJ/81jdrYBsFKaPj/rjJKIUPt92oCO2/50hd
EuqsmLWbdFiW6K/BhoIk9bzvDN4YX7JqsOsFijp3VEdYB57T86mACnLUO7ccQDmCvoJ84Sk5yks4
a0pOK3+NMR0qaRMhORB2HeWKQE1yR/5Z9pRYQY2pVWa2Nz39PTw2PSiNnJBJQLoxvpYIA6gFTW4Q
8Za9a8esZserzJIXb80ecDFuDrIS+mOsqwdy1BNOYg4oKejn7sH6pno8O+F9/z0Khfbdn2BFXwP+
pkx3S1jHYV3hYCuwBbqS3D4q/TOIpV3e9pMzEBcRhc+xb/K0ACWTNp+qb4XA/t7DEKFlbZAmlhce
8INVuN9QEd8fe/x7N+1IPh+5WMFta//BEZa95kiqEcEQKHcRSoUm9RbAH6wu/GunpvhNJhl1tCY0
cWb7LZJt2rmFSwyX/Z3I0wUIYpFdshUc9sUs/Xmw3YRT4biQ2AS+4j8MTV8pZbyBd2l5RV76kYSM
K92nPKa3PZ/0LyLGcLi94IpBV3BTJVu+i/HkcDEnNpBKtSGWCyxjRE4UkKQMM7FplqtYUY20hWTG
Fb2H+q90I/lvnCKOK4NWerYKoDuSINM6DZqtOkofCqfYdNhd2rwYuITyvf9rogb94e5ghLhcB1Cy
cQqyLvLr/2+AKEjAy5PjspzZ7XjPfCH7T/LUO1Sw7SK18YowxEmHecCxMzhFVG0xnL6J+a+mTqL1
JT3x6pr1R+cHrHVeP8wZdzcslj+kc1a02vgpKDeK1zGsB2m0JyrnY+c7F6nnDEmT/hxToHCTH+6c
PwKno3EAUBEA9RlfGKSx4kibrpNz7M8lo/+ylcez5M+UBliaZZg1V5fT0S9huJkP+B9bcXOtONQZ
8qA41pIumFCkb+ENkqWQ4iBtVfXg9810HZgmcxnX9rs2vnb5Im8f0IeNRxkqsKtg+iliuO2gQ3bE
Ta6zpwln7ko+tlCKRJZCx/36u1QhT9PytJ96P+vSEiqtvrt0hvSV8BLQjR74AQ0AyyeFO1+QxKgW
qEbW95oRrOvKUOcP2qhr+JBtOKcoZQ7pOxTwjxnEGqjtwEYhgh1X2EzA3q+/qJ2LJe0NwyuT+g4q
WtxnjNC8EUXTiz8dXcUilDj/IX4UTs9tmTHnOZrVgNk0DScjkRY+843NbZw2t5ixfQULUJ6GeNDd
TVylIHGE8JBoKu0PPaCFuQzimrWi6uvr8HFeTo24epy6bXie6a8UiFiWx+MONBcUkREPSu8z80TD
/n+dmRZ0Aw7RflA/3SDKnOrzphaqMU4sm5TtOi8cB3uw8LnGY6xbF1UHud4PbnuWxQCg+qIwJZ4h
jk3ak/lc09VrjFWLGLUFmvk6/yvmRZRLkPBU+t7uQzRZ0E9cMm1Lza7bsoWAt06PZW3HAdLSnJQ3
O5O/PmdZ2VGWfqg2Vm4FJ3VH1a+GdzLIUiSjsZJN9kXPbLW4PcaG09gFe7wk/olgCHApJBosc92h
cIaDoU2ONcJM1QX24IDmxuFF9Wr2WKewmy6aefJDL8mXK30uywfqY+pkPje+j474z+uYwnFeS5y3
ueoHqFBq0+xJXL66Gzu3LDjOiCz41jFfDwT22pBknRAeq0OM5DTs3kzrqaIA21OVdC8GyPCC5L5W
IQCiKov/je6wJy2QU46YCBtEnZR7rlTDFjSovozwf1HHYCcA39LxE7g2Pqkp3bkz68RLtM3fpaJ1
1QLeXtH5VB1Iy1GxtHve19ETr0OHMPEO2hZ6WmnmEJ8yjbWnj6bd1k7lb2vYInubBRWth8r26/pc
xhpP7oUpDXzKmLKcGtFJjdMIEHwJJeFDGJenHTsDEe9oTaibQfofS7ImlQII2wFzGISe3/XMa/wh
DQPIouTeMtfc8IR0JxffOQN3Pd4JMS0rCRAF614MzVbdnC5U45XDmnJW0SRuzo9J9mqdzIQDaJq2
SYb60R2jZArP8aMuqgmiM3frx1vMLOONqTHRj2FaPdReUAc1zebSwwn6FSs+1+ZUBk5Ir5LAhVvX
NZ2SRDDhbIdI0DYQEZrq4Y2oBJ70Nfiq7z0ZMGMEBJvNacWdRw6+owv8H9eyNCXp7+LuOiCTUQ+k
eo0wzUVNK4byp2WBA/+90d9bR6fh9MXPxqfByHTNp9MwVXNVoUguoECOu8XUG28+ZmhkvI9umZVv
oLJzti6wBgFs/ZWT1PT6VmPHLBqR6o+5GtsCnV2bSbp3EtDNc/V8zWB003uZj6lDjz4iIs9JRKwE
P7KZHlW80VacZW4nHfxn90/FA5G/wLfnuiwXGkfw/XUdrtsNPYWNJXxnDhizZQWBQK1BXgrcj1n4
ScwsZgdm6r1WTxa+z+bKUvWxGslqyRlAR864gsO0rhjUE3osqgNHV/hVyyHlCQBMIdOLw1EiVk+c
5BAxm6qYlvOgR6Cv8iBcSow3DrQRBYNXIxJLD5riZshi2fxJcaHffPIsnt7pD8igOyS6q0Gfrooy
pfuW+uym8n9d+ogTCTtAqN67li3iSHF/Sb7utx1WEs1nDRjemjTNtqUmOFtDO0cBxU+r2ZpBJAVG
XyBPMf8RXSy6/z5y2wWuDIN59pSb16y+Dybx/9h3R+nYKKiFJBlszxeRJi2kBbp8F7nhoS2cqum9
zWiYlscxvrfC/CWRi3vcUPK7HZM2gcN9hk8SDM4UqQMrsgQcwKAQnUfjguc6PflK/BzmrS+pB4+I
Z/4OKcuZ71zlPAvLklb8IvCS+g+qmVjn/f2qdxh9kv08bdOce4P8fQYqCfrFShz3Ula/Q/PG6pVq
a9vRcY69J3NDkpSOml8xdkBzVGET21Rn8feflMNfBPyD2w1+yGmNsFpUY26YA5KQB0xACcC4rttJ
sPgJaOUZCaw2Cftm+eLUQIUcwSbfvsCHrLsYOy/S0KwA5dvqR6nIz5paX+7pyD/XV39en9Vjhede
ROv4W5crAQoUOI9aznZCjo1CkdHORIiezb2Rp4kcJh9+jIsnJzQZnjWOclsX7sM7vhHcy6UUXQ9G
3ChALqoWLQzA8DnojLbqFC5GRjUIi0eFROvVKOsQkCruPw7v4sVzpoBPeud/+YSCYZlE7XcirBnp
kpep6LprZjBJ9vPUky/hnSFA76QKkn9afiRsZ8piwVRKRsKAUYdVDNgfj2ZJmjPk5iID28KvhdnB
ISrJ7z53/NWVusJx+g1TfMMpCDo4K80zqPVRBHG37jtM3Emq3EwmAn1KbIEG0YJk6k+Zdi10Vz/d
sky0sI2ABOwoxhmBc+8hi7sj7PjaTpkS4ZNTjypiLOTf3J8qTUM69NBheEDH61OgYTmSR1zVxPvi
yoNOH9n734AWQIv27WCl3+KjupYB+zUbS5DAMNZKCFzM7Xc/m5UXd+60jgaKJNAkvVLCjJ5yLElA
9jjd3Ckqc1NDVRWAu7quM8Q1gUaMcwDrxq4B6Kb1SpiEyXCI+HYokfW3GLGjHDGxKvcq+7X77meT
IrRajK2jA/XHD/6D7uYfEzWuLWN8uAKp6R+0LmiaPaPDoI/YZAy4Y4RiyjhvpuObJ7NLsHejuVZw
lszIKdaUMLlxa+NITsleNcMVNFVFrGCV++TZwjF0inizbUnJcE+ZcK+aIGhbwkRcKCjm3wFtT9No
8JanQ3BM/fFjsOVKLkeZsiEYsK2vx9TmljSOFNJd19VhHewGYwfhGX2/eQJT+1kNIwTBPm5BC2wC
8uaiI8IJLDMn73xTcsjGenM8oWMm7A8aoZy1YiqZw+YUvwpw6LDFQPwJaplzpGTI2LhGj5ZoGms7
3xPCEEGRSEI8bCGtl2uCxy6LMPUAem8NynodMB1+If/Y5mifSRBQO1AllKi9cGEjcpcriw8QXkU4
p5w3TeUx5UtiiGApWUmGHX+ElAmcKUrr5KX0UZHsftgYCxEQ9rXmXwZUx1EyTnjwaN4L4r6AnsOV
wwtgyEIdZyjmKuq/OJOcdFbfiz7ANo3GUzhetmNo6wd25GUks+xutuvgQAEevoCc4XMGF0yj1dcW
kCvECTz/Ep3WZoPE2UA3USahVCAX01TkVgEE41MYAYtD5Z9Vr8kzEOhNDgpNDXS04fy7l7Vul9Uj
9RjVWqnXC7tdGb1jIUdK6KA9BGwbxot1/vM7tU0uXk8LCuAHfoqDS0/Btqx1mN2Y+c8LNYjpomWV
deSb2aKqhWbDejpOueA6NFIzDFWVFGAoi+ARI76f1b3eLkbWbr+qm/9DBArM4eWGogJXAhub0FDp
dzfytHaCm6RTw5BXfp37p1izNbSRPfkdq7VeURJMJdDlXENxQHv/WmCtgpAnTtlOT5s+bauP5oAF
db9enJDOc0BAGGY3JnA2pcLsoRcWgztodBrbxm+PfHZw2q/DK6Q8z9IuHhh0oQS8Z+/1p1Zef6WQ
AsMR+0FCBavgyQzSxJHRNakHvjE7QMFJnSFrIhLIvHgzOk7CuQcRsG8lTt6bziQoDQtzcXA1n/X3
ye4aJWW8RK1Z6C40jdjfzQCW17iSeBHoDfbPlaLXQ/B4Ck+Xeb33P5MiEa4KGS4276Gd8MFGck45
cffZTrxgcbwtaq/0JfCZFSTAXtv36RZAyJusZnpyWY93j3MQFvMWSl2M2H6o1L5HaUABaopwageA
tORw/wivMnYLwjJyQQRnJvPukTOp5xIL1YxwyJ8giryyI0j9MseEp+IdAqIHEX2zNJy/X/PgTZpd
CfdCpvZ+ygCgZPGUJz/CRxRHNu2lcHk8pwnKD7EcF5jN6eNFmHFkK3cKBKNhavNgsasMmvgv1TlA
0FGC3koenhHpUtxpVoGAxL4kQ8BYPaU8B1WCBP8adoDdjCQG+VPMs4pS01VYi8g9xEDIy46naqRc
eRegip4oPLM3R6liMM+F+eTY5ztb0npecA9nR2XNlgPU6VJeYF9U+YM7F58o6C3iO4sYqEPFJrO1
LKt9Z7J8x9me+fU+J3I4EUeSL5fHNXJlIOImXMzvQ27JFz2u8ecT2DERQxGdW2vqD0R9gXZ14Izt
fIp9XMSnyjVixw4TP2Xmdk9DwgfNHK2g4YBldusweY4AT+Cq3dPDdZkDYr5q/378su4iiNFYWN2+
yDuJsoFYAyrMi9Ww6KLlK7tY8RXVppsR95QmUriDotfhDC7Crs3T0Yk7TGbPvCci5pYEM3i3xQIK
BK4BAbLKvsjRUwhBIFMKzvv3Yea2ihvTfp99s18aXb/fHDvLX7zSdPUu+Z1AB3ESZVawb6ICTZyr
+9GAVcMsb7ZsqrzyPRk1vWUy9irBrwJlfzFSwPQZ3GBB12fsdzdE8Pioz5DgUntgxrvJeSCYnqtE
YTuVAOIx6xmudnCOFsMeNzkbfC7FqXPz9q/0n6LdYyFeuK3ER1QKb+B59lUioi6JU20MSL/yP+64
Jhq6pHseinHWhZnd+XraHn4RLwVBufsRnmHKJBjKwJeXDJ2HhI4jsoKVTMcnWY4p39yQ/hWNE3jl
/kgOauxa5ZTygqmdKwFd/psO2XOizFey/h8uq+MXjK/5XCXPcYZTZnIJoAim0vlX3S4sBxTlFWCk
fd1RzBUKXL3brsmbc3ZuUDPd1/3vvljTHobfuHxpKM+dB9cxgpMoraOuZBb3kgFbrDo5T74CAzGB
ScHs9chAgR6aBkXyaoEUmqLpwbvOz8cpjv32JJHFG4p2v78RodxqJs/d6DXEZrte57oYK4lLp8FV
w1x80Ia6tIfKSCl9YTD5/AlIQeBOYhSL11cuer1rUAXgxw5AuqxizLoxcNtNdMPqP2sRN9VasvGZ
Z6e58CMT8xWib3frFYEQTJhlQNR8WciWj4wLxfP/oh+ljw/tCCoQIxKQCFZr+P+QtB27K4LxdcWF
ZdJxfeBixNiSc+/eRMvhvNi230F8yGCv3FMfnvimIl/bGCa8Khx8aCFn2rfStIk4ooUVA58MspA1
v68BHmgJCtL1IJ5x4Vc8b8vIURgqgRWL5iuNMMzpMyD+4tbad7bUbaw8pRv/MElQHqmSsuyiYUXj
QRRpYuHtOd1WhfVsGTG5tS3vV4ydcQhjI7xIDg0jvf83n/xKwAZOqtUZyE704THA3+pS0hYX+zLp
EgRfEmQNfJyDUx988ohCCtArOp3ijOGUOrIPdp/1OlkUTuYIqRwbELlWq/Gy0BhZq/Wp0GuZiVhU
fGegU0+OFFdeLSiqMVEGyOwA8iNmjMUKDWoHnZODEB3xFl5YYauUn4qrB93CQEsFC/URWgXcF6tM
Um5+lCjRLK7ouaeQ/cHOwbtdfy1boTRzKjfwr2C9bjOFxU4JBUSiqsbv/YQH8nXia6kJAbNZIw82
5LhKJP6jbbkr2MB/q7VhJGugyRa+uHO6BPTmR1Fd3PNxdyvrMAgoJmylw2q+St2FEtEGZ1KR73Jw
BUoufuFr5fDfdohLQFvuBAJ3CpK6RNSk9bMP4XnmVx3Dmsmsauxga8fgkLNXrWFvzXGG6si71jVE
LV34SuE5S4AJqSfcDYrHhT9md1UEp2rrdtHVD/2Dewz1/aBijmDSoaRMazzw3q+xlAe5Xi9RAx5M
s6Vvj3sn0aC+72xTJOKWYRkrPl37ZpBS4hrjrxkfwlT6CwVXuu5hf+DT2Svr98crMgBfzFcyzror
deqfNhTAaAgDiD1QieUDlrRuJjYfFduENb13LAn9Pu3l5kEhJB8fWMbudtmk+cXFJK0TXWflQrJv
ERZLzGsTYdeTRWrLNVrwSrfv1P5IB8s4U8wrT/jK8k5ApGkkLu0Rwlz9/fNn8dqg8oQyZDgJX4AB
su1eUzoc40zCsW5mjzyDwwFaVRmCAhtSjn2wmy+VMKMu3ZUrlUxLviRPxsmDOYdfq+hxOfDeqIB0
Z502jdnd3Yl2sMM2A6hQxlfQblMgGgM+jTd53d0id0eNFEHZEJhXW/egIKIiYX27jChSTkKwWv65
CM4LBow2c7b6/aSrm4UCKPXtVm9VbnHgQKtUHZO+dMqHkbNrt4nM5783ItmMAQKxAoCZa8Kbxo35
cmwp+ocwQvM2WyMrIo0VhTiacnD6qu1xEQLXvhlBEBaPalYK7pUAsZ49bwfHvk+mHA8i9NGQXtjb
eyhn2sf/2PCoXDpKiKKAmCUvnNwah2tPtLoygwuAfIboHsDeMGw5mtdoi9ByLNbNVJ7OGkSuyoT/
iJCkNoISuiPczo5Jg9DeZaMyTfz9CpjrurM/79kNtGY83fAUkMXe9NKIbs754gzvhDpCnfibrQtp
0h2YGMA7ZX+tvYWLvB2Crr1BjKfPGgboN9SdmhIrQFmR7ICuLIgMMrCnh1PvBu9ZBiu41B29DdpD
JBT1RDVvToFxLW2EC00h14xgYJCBlr6i+YROwlpccLRH59JcH390egw3SgTDceR3Un0JCwxee2fl
32/ocILl5G/Kkl0hh9QE/hs+cVjugXlibqmUwtfIdnI3QXclhd8k7WZflFti8RuE9J1PlPvaoXCP
E/Yn+w01NW5j/pD1YaU6cRzqWW1Lyntlsm2UV7ISLcBSbjRRNpfkqFq7lDCok7h8mTDGFAnCGCs+
hwFIdKSt+DHzcFmgrngPI6cXPKiFonxqWvkCu3enGFEuCHbAchZ9EH/yP2oI6Y4QZ/kTIIXte/C6
/5PkJ/ZyUal4KDdSpmTTq33h8+pP6W1inPmmkpiGnIFWBx51R953Xz1+K8Q7t9I62eDsO8NWQfTk
3ShWj22KfA6Wm1n/gleyuyGumqP9gB6Gi0qLum76HMvy5sHzhtAW8ykIIRzxtn/NpOalQQiwzWzB
Hq75CGOewguxczwfYwAf8+CQG1GfXCPViIB2lPUKwy48/zFM3u2cbNuo74+cauoq3butjmWktAiH
nzNKv1XtyTvcD3/d+HCcXPuZ5PhMh3w0P/c13zGFkOcaKTq3vsemAwy+hRarLNenShJCgsZPyHZ4
dWhXMAO652B5VgMHBjuo+GLClhCDdttou6fslzI0ksyg0ha/1KDylrKIXRYYqmnNqu1PaRh81MBn
isCu+Z7HCykwM7HQ5knWDy+t5HXUKBKP8WO5b3ASdlDGTtL+FNe/2caTuFlJ3U7xFu93lcZW2Do4
AhZeMEqq+sOmGik2Yli8xLa/u+8vhsYGEbj2t4cGqbtD0I9RvmtSwvLV0zN6Gbh7WEG1WL/VZrps
amRorgM/Wz+pOacsR2Yh2BMbu4NDHKLoelHGnB8UfC1bk9WZdB1lgWoAwUQghpILOycUOf6p47O/
outzWTfTbPmyAu4kLOoM1B7ApksImr/OXTzXw1tuxcs/YDdsewDzn9w+3UAOiy0VyEyIR5P4y23l
j9djeh3yd1/xmMdEP1EL8MOgk0EGN8gizCm1DnugnIbWUsSW11dHoH/Dz54vmF57yr/N5s/UOjqB
r/D+kx/NqWaKoUvB/wtIpItLYksrnkIQphk7kPQet1UEsZaZlnbtJIVjzomaaW8iLDgCHp0oekPZ
O7RKJIC5cxfSgAEi4MNSWxt5grhLptYnbckVx0WiGjeak94cG5sZ1Gf/pIWdOnKLeV5jatIn4Pd0
/U4qdiY04kDOBnz2GcxINPnAkdA1FBx9BCzwg7grNa6XsDKMF+at9UotbC26y9H5/XszeA2uDkl6
Df/CDJhb2flMErF3tF3uAwWaX7BV7q0qnd4PjYiF8rFT2VMWM4JuDPFbWALqIV0EaI8O0LAcaiU4
xnDyFU9mHqqRQ/3OE3Okv+0EJFPWOOXXnkSmdHf8es5MnjmYVkgvkAgGAUgG1M5NppB+18J99P6G
0RpCSRvEjJzKvx5bgwlMu/S2vB1Pw17c9usBYHvEQ9cktcJ4uVBj/ndNfF9jrxiIHSMeDOHmv9wz
PFRupYkVhS550HZnntIeFmB9srS0dGs4fGh3CASnEw+mcgqu+zWnK/IRhh9G+OhSXpC9V+U+tesY
GKHF9A++se6IiurC2LrZB6ANWNFM9Al94fWSB4amOTBpLFlwnf8EJ6nafRy+mrpFXgu55hFGR1IE
opBJjn7tJLDRqI5bwE5nfrK+91CLtFjiAnxL/ojmuD3zo3euBzkLwotMB3gfZi0KJwrzHmoKnk5/
7OpBjam8Wxy0D2yfQ543YUjxYMQypRkaEY/D9GqmkVMe3cQxiRAxSJrKBuukNfa0mB5KVq66N+2D
MN2K/M6X44FQNl5WGfxtuXYaAzvUiFCLzlcsWS1VnSP4vCH62ITRg/8MQZI79eXJBOK/GSNjPZgz
vzbg9EEI/9J2EiBjhrCwFQVt8WEte79swoLjBgzW1RsnJsezKCr8uNWvkxRrxaadGFdcqq6FyImV
dXY+oSOyHHyhtIowXC20s/p2J8gVINTTL7lzDIXcx42repARjYRjgKU932BIE9S/7hNGjoLy2dAX
Kw+kDF8K5fVk4d68Hm9gm60fQzCO1zNXTPa04JdZAdrHo4Jgzhf+qk0tPGhINU5HVz/ooAsluxja
v4jeAdpa7zbACTti3bKFMuwpFNIXpkzTreDF0xSvpQAH3GAOCsr8ATSdmVyuiIjMxiNJ11oyjfPg
yyZ6+Cp5qgp/7qTdezc0NDUBzJMOeOBCRaym1IoIeGH8QRIGo1Vj0a3h+FQOF1BNEtfXW3Hc2gYX
9qmYhQgs/0PwEki69RxB82uGhc7MDTLgvzALf4edtdyXMG5K+KjOD2X8YRV5xJZlo6moCBxlOdwA
8YQR5KULPFiD+dEr5dAJT7LV/0sJYPS2iSFG1M+gP2QFugX4s76JNLhnC3Wj6AAouPTKv0qVEO8O
9p3CgOMt0HAT0HsyGpoi8UoO06gAtjRZcnSi7DYDWSuReEm2nSQn368sjCqf1d5CrnOFFTVRAk8V
gs8SJSgK5ElO+xW2PeoH7UIX6PSOfj8QTARdDpSqb65+mb6qwCs1D+hIom4oCvqHi90ckkYYPAb6
eGKvK+BI5gFy5STTAoTyWArFtw4IrCH5AeOZ1zxYI4VzAzK3f5AZLQEaOIdWMJY17SRXO3XEHPB4
WiS6f01NEHFTHJsVwSyBOgjFBFMcf7zE1h35nlC0h1Z/AGUsJiweHbZVX0pn12ubJTAUscoTADaq
fZeTFMBO0szXpECzkcYVIREGsKDUfkSbwqGhdvEFkC9m/W5trJwCw5uxXWfJU3PTGg4wpSwYYpUf
7MEiqIBucsbdN7B5ALqAPMeXacK1IZXb1vBb+fGQ6TZUVqrWC1iM4QBzbxpd0Ast98UDlivLKeCQ
mR3Sy0Faq2RbAQKf52VKyCrKgty+Z+4iS1rA0p4sFFNg0hC2lnYcE43Fz2ju3WLuj70ccIlV1VV4
idEyUIz72WOkCraXNzLsrG56rUZd86G5zG3A/d+0I3PDm82+CwozQ6bPJ1UG16qSKkgOX24stoXR
wSWoiLo6LsQvRrTmI9nJoSPSCP7keYOOS/C99bxDFKIJ6uVc25sBbdpgzGVlt61nd+T0ysQo01le
11FWkodFwLDPso42gNcK6md7PbPdwcdKlhNYMqTFXEypoTKtl/g7aPmonPkiTbTztsszaVwtAdf6
tO+6zFr7hNTvhK2bND6vYV+NDZrBKTx+9EIP5GLGVSnXDwT1tx+Ks47MrEvnce67dO+CmIBY/wZ6
+Ic262hzLQZAD3+f8hvX0ZoL8o3rKw2WTdcTgZ1ol0yHTZ+8Q1RwCqD5nZowW2sIhWkl5Dnhrc8y
ZN1obdW+IA98BmZ3UfyCTJBHXimPrqwGYLJ9kcHBIGo0QM6cB7YAQYohwfC+LwUMyx+qdS75+rFL
J/7acD5arD2un9e9F3i3O4CXP0t+//v1hSU32hSKVBpQzDOhZUeed9zpjMoB5CLog81fTi1/INDZ
eeAxt5he200+4AyFdvSNmjLRnr7uNTGNlNMp0HkxryinD7iOec3P+UEQwVil+vs8J/lTmZ0dCWPv
0Md9gV4FDnOMs4OF/2GYHe0gmf88LFKetW6hi+qUoCfKsLF+BhLlfrdxzyxPWQzf0Jw1IrRapigQ
HS5A85s2fw4JWHOMhyYbqrVi5AM9MGZglffPZpSMfQFun9AfjlsSjV5A4SaSD9+k0kqjSMr7rwIG
F45NDpQeRm4AUuXXWpVixgOwpQw3NZTlMFfOjM/C/6fAK3fnfJcWJrJynJcglaCqbit7cvM51lw+
iAOu6xhsr//daMk10N6Tyv79bKNDDIVI7WLXUVZwXbMJykcXfz/wNW5YrRhJBBeyPsAQ/hFvCzMq
kHJD8pcVp/Oq10Lry8cnZf8fMzFIB74fU3kQU377hYp898wWso8jGiWerZSdvUayFHiQRzwg7c0U
PL8VmV+raUCpRpHcLy+l3h5Ofwza/xHcDZuXiQL+mKZgL98J/RB5WM9Q2axvpVRxBxY/W2MBr39y
+PcL2pKrOPHM4jkTazU0W+qDDDxeehYxc2RWMVNNV2UetOlIh0OmY19pD2VM52mrCvsfU3eNpJcq
LQtrAGt+KunsAXVx1YaQ8NXdpQlLprV24r1/hwP/nk3lJX1owUZmL7MEBajGadapqv2QQFiajPom
O0mGra1cUB9b3qC5U5OHfYASDwyHCXyCiAUIeGkwQHMEA7XC19+jsRO2arWlJQTk0mL46Mf23O86
+cN0Ke63ctISCfaKyDm8hVy5jgEdO4YjpKzMXjjblt4gzpm9ctCGZpMbDiQVtLZzwKUfEIY5vbXv
r3xZL738g+GIMMphWN7INMdXvc8VYObNNwz+fDUlXXdY65UH4GgmCIy1AkyzLTiODQNjLSPSxmlb
VX2jpEvSIP9X8aF612/76/XHuF5L9aT7LiQqt2qH3AdkPxYgNGUEkLe30AuzWb7GZB0evn4IShxQ
zCBSJbB+SONoozS5tJI3zcyNEg8646wmhiOsfD6zM1uPtFxdnRwXVBUUIqXInw78C4gLTP45mXJh
Oyxx+swxJhUa/ZwMWPfZ0X2pLi3bIXA6d1B3vbrtDkcHRstma2kJKKbcU6o9PdbU/v/hYXuZ/Gnd
Ds8QqB20hz68Vm32mInCVlXG9UUlrqVcFcx/iyeetfoGGyviQ8Pe+r5N1LRevECL8H2Vgi2/v9b9
EbkcVygamdQ5mC1LNqfEE9aI5nksFGGg7rKlLGKv2aW9hqjTtwAoRDpKAzQ8sUrj+7Mxo7dajPB6
F0aCx9yhCzbAT/Ajlwn0GMXmYxKqVjeu6Jcm2cVHWfJScxc8poiRw1Q/1XuYJWeni1q8Z2AYV0eC
squR1a10MM8Bp7OTD1GYkXNglVTxcu/+6LfEBtRWymx6ZNfFHiCNdWj2j/dudch3DLUmy3Gdi7EO
9EE4eCyjOg36ssPvtP6WcNkQyKeOjEZRYmKhWydxclOLKvf0JH14iRRbL8/yXTa1as5gKLZXknS6
UWbB8EsLYKVdusHydvtFXNVJuwPbzvdC685mbmY6K890njPajXmR03AfWyneuI4pMpAfMFc/1csT
IOFDEbyyiBZcXVlT69ejdqEh9+6xZE7Vvp7VfDwHYkyMxe4xW/GvuWJqRaD/P3MBdTNPMmGDwtTy
+xDAP3F+NYW+9RMZLf6vimGsndpvmKT7KegSkckZ/QRtFF1bFdMH26LY4Ly7B8O+JEWuhIoluGnI
6zdXRcV/H/mBIIfsZ6hYC7DTePMc0IeuEahcy6HbLW+mn3vi/r2JEdip+pNoT/4CxPfBi431H03I
hyqPsKko00S7rEhUgTscI+P8kp/JauumGCBxm2TUV3Nv6cz6YdQRs46eXCey0siNIB3MvobldAd9
yxOVeV+PPzKCQuzDyvZEDyhK4Kc+9g844KGN8GFEDNZ9yALiaT4Os+ysCE5KvMwvmpcvlC2nP7eJ
0jcezwI5NcD+zIqLnFi3FtVvAJcf0Wlb/Iy+qi+TpvBDjeJDXMgMFYXj9MHLSvM5GzMD+H7kQROC
UJNyOfWsduI/FZ3az11Tzk3o9WYlKpqKNnYDEl0MR+besMzDMDglTxW+23MAjqyJ+I7u1iRDk1gz
hLWH2DE693ae+bGhdp+BFz+bWaG7DlChBcezr2nZa6DfMefJhzRNeU6LPvHeEnCl5NCCYvknKI9m
QNj3P1tx2VRH5iVMSWaQS0X9/Fq6KJAYdCE7gPABi6FMcIdu4ZU7Cz2Su/BwhcBcX4aWoS4GZ6hB
/YRGLomZk2VrQowl/D0gXeoFVR57Tg26BznEnUO8eE6Gebj61MsKfXVWsQfnItb54ocP0UduiLX2
eYA16Q+5b3jfdhoyV04M29NJwUZFj6fQwrDBPSysatgcz0QroIObgHkIBRHR4pfUfL03wuO2VhZU
02tuq/w4suJldhZaM7P0T5ACr0p6stbEuJ7ng6dADe2LibELYE2+p8nttRQDUm6d9m249DKcbrNE
plPkFBLL9szVTy8KA1qmdovVWSDCbV5qWBrBFShpH4COEKUU5Z4Vi76UaBhMjY3wGEaWxc/GnjyC
rTl74G2gstBpdYIYFQX6lPX/V/q8NmsoTCKRwoF8hPzKBMAjA5Ja4pSPgsQw244VcpkA6nkIKWOE
Rq5//fQhu/kPTLxtnQF78ld442sR3i/c1TC37sBKd1bbr1VxhBU+kJyvwDx0pLGQLmiNpcjBxUOf
/9Cy6X+dgir1atr5GfoOcaFqUzqPUWoRRY2vf7U0HVapr8YZwtIgRcyuCH1ZB1NccE0uCDxvBwia
aMR6q5sU64VUvTfBnu26OxsXo/5hSqTjnbWZ+W7SJCXk+z5hgeuVwGPVuuPZvZ/41gjtu6AUvJ4h
uhZz+M0e7mF6Jih3vmTUIbESt7ZDke0gmhkUI6aCRHRa+m2ajNd3Y9tyLO2raCqvohzIAsUOa6G7
13PPy0gJBQOlB6XqT1qJoiP1rDMliaEG6bdj0HVo8RqblWUBfYpOkngPqymNex070olYRpFbPWsA
HZ+HWZ9kwEENn94AWwj7iSEUbPYvhRB1zEMUlLGtgNnKKWt1xQGy7uw5tjWRjq84u3cVHqkP3Q8T
Ee54smmfd1gNPDofTtphP0HPOXvKf/1ixr3dnuyQwfRqPc3p6m8wgpXI+MDkvbfTQEwNSFrk7hSx
t3uO3I5uaGooViQlLBdeWc5c10EJLvzlUg6jEZcwA9I6cDgDc+hV2jXyHAy5Pe52Iu4tfz1VImFp
QhRFDTbxNa6nsrXKXBOfQZZEQ67hWNVi2QA5Ec+SEbbRiwrAMtWLLqpVIeyZ2WUgkCJEcJiPS14L
Qj3PZfuT36eKBxeD5fNuxvxmiIEHbN9B/PaO1661mkawYOb6KoxW7kxbZS7F7WfHWo06KvR68fUO
DXfFhqL5VqfWoZr1jdtVvr0jEDawp4zWSN6DxhuUyvRuUiKONh+YD+XzpS/GhOjVfEVylQ0lbmkW
luIiJILsOfc8fJF0j2LM1xkm+Duh7dp9nuCbbqW/JLPJv0+DjLUTId6YQpMLRjLPaoc/nXpKdHkC
28u/Iemv4LAbz7lYn9X/IYID7GxLJ1HDl9g9BkveIkdlvS7vJgKL3l5ZvDnvUPuohtq1KsUslREa
bW4H9TFHsNdViEJFiYCcloVxrXiTH4KbbEL4SeffVBUYTacE3ZD2k+TPRdxf1nScqWDULucrFCpG
aiLFBgqlfGKtURead86ZI+y6IRUmFqkbjeOvfgU3QX6gR+0Ug+MPUkTP30lsm6ctmoK546X1r5Vx
swsr/dw5TGkg55PNDb9veJDoHgDsD9qBc+nfVPmrwHJmWcuPw/kmkuh6SNJarG3UkEFCtUiF2ecG
SSGOTjQdcJsoP9WuRaLLjfyegiHX7MYgNBi78DyzxqznWOjU57zSvbsUWg3F6TEPZDGJnpyvKVaT
TJCbHWZJobzG90uzuzr/iJSI4hiROMZC/M7Uzm8wLEEN1W6MCrC7NSm2rf4YxnuokMHkrQ45o9pl
EeIKbU94nbjL7GSIdzoLX3g+B8MdpNH5YbZFEQedXJZh5elMarh+es8RKkmT2NpJzYTk28ivx9RY
Lc4PVNejFC2WxKJnY/ihDncEMjVa42LyhpU4HhIcTn7xWsvIRUCWkyh/x+8Y9q1Y/KPbtotQcTAA
Tee00tEPqZsdNSMsvtDy/fRWrAeWOZZOPDk9qj+IxldIpGAR7YLiL5ACf0mOvkxZcQg5IL1+XI7O
ER5zpdlZApQN1xitEzWj1UPEMJOWIyvB556q3tVwxszDGPuJsbbjcV5RGC1VRWqUNbXfDBimKO7L
a8kcSlMQaXqiaNi3mtdXgJkglbLkCMvK7W5x1nVEcOLVQa/p4ihMsRbJW9mVR2B7UQlN+VTJqn+J
uPML0m/eBxjSgbSDG4m8eEFzkP4BH12TkseCFovI9+tyRXW4cVATGhUuNgp0eA1VfBrf89cpkzsv
119Ucc+awgjMsHJiT3DmqQhP2nKcdZRP6FuOqdFH+frPuSUPuqGF3CtDk+rkK6RV041Ha/ON+gff
sBJToJ4aTcOvmymLsKaV9a+g+7Is+gUhkgY1z/FugcKm2mEKbsLx5m48eT+lGqMUhkuCSkFMQr5H
3gFiusxR7RWWsiw7uFyQC+bd3J6ctLEi2ESZjzxHp3p0KUul7rSTlC3j2b7iOopYe7kb9UN/5Vwj
SpamCRqQK5wVbxKFTAsxYqF0P9G97WUIwO8IV+f/zlReGwDARNaOJA7iveuHRWSrTXvmYnTkgj+/
0IqEgd66PXnruswAs9Wzc4zU2fdj/3gVyNKr7vriaTsSJ0PPoc2+s3qdB4xX1Zw31LKeXn/EtSHo
D7lJyOiRUrngiN+cC36His7WKrDdsQZjodu5RhrnCFwl//tNsIjeqn/vfecBvh/EEbQ9FPPeFE0H
wDSEr0t38uxpzBeuCxu3eIuSWAAwcUJFFvelEJFPXPsXrJRbI2ZS/VRN4sWkpwa99Yu9XIpvUhLb
xie4EepQQHe0zgPnmJquszKyT5tn3AboM725bnxbOxYjqozsKy8FHWDxs7vIE2vF6btzgzBAsSNc
byNbyX+scItXGTpNhCSoMyC4jJlKUSRbCCMsCzwkpE0cvMRTEXoeNYtiJy08LOZFDUSi+cgxcqrH
w4FP3d5GotyziD6XTOAOPvhGmSxHpL1FtSLSzYdxQwWEcaNq/7GIpcLD4ye19/JFuPAXY/Coxano
ln9AgrtV1w5O/FLKcGyuXk20CHQpJvKN1S6UPQBl5SjOWVxhaeUeHlJizQSmXV3iERQu2Q3dID7T
gp0ehZ65SHr2vNuor3jYq3rG8I9J/NCd8Y3Im+p8tqLzqAfoBQ9DYsP5CdutYgvpmUVHfDgPUSSO
25uoEVgC3ki+ovKuHvgEfZadpqJ41cpAFSDQ8xHwgsc1oczo9Wg2ETWAM4y1OwE2JLxVKMPldNxg
5t++qDz6vYd1D2o04E/bhQOenSpUxB60IDcbCfYYrq7ayBpoa/v7HEt1K5zAi3uDMQ+omsz1pn7A
ARrOTBY6g+Xmla+IIDq4CIocDwJeFzPsPKWsOtp8RKQzfWGcIEr4wojBD3YkTkAg7MXCBkDNpZ9l
jAgHYe3RS4TROgPNmjA1U4pIpLPSACAZjyPy10GruJOZ8GbZdIEuxeO0NniskaztbzzTgl8N9UXb
MCWkuADak0fDNt2O7FER+9XpNxoexviA4ErPgqO9E4JAOQpocFqdqQf9AboGT847thKhJM/zpA74
D9cKiH3m27D3CyJuRs9hxgmOLcEEsGtBRhauVADYAu+ju5QvFUbUIQnuOY+OdShfWXvkILIaO8XL
e1/4+cb/l44zWcMwldHm67ata6mHte2EpVh1lLG5SboTV2MMBwQoOm3x5xfgzvQez+ZJwaChshHo
Ks7K+1ADC9AYz/I6wXYX8o24gjI0jsjWqrRQxyXO1wUPO9GVXos6B4dWJnqbs8fVRhLrm36OWncA
hqNJo1I1dP6uHUTvsNrRUNrrTxuIJNQlgxM2foaU+O4icO/3LnMvfadeoWSkX9FPpbLF4EljHrSz
siW+WjImKWQSfZlInfmg1h+tl6Vb9O7GBgqu5IHWjN7Y7u7tr+tWiKlpfsAdqkEy2RWN0bJJ0EsC
P6j+NG+1d2BoMW/90AruwuBm/NuuS9TY17Aih3BHvI5pORxX1eJN4TNwaJ37eNC2jhGPuaW/LdIO
Nsjd6W9XIdRxNPCuRMf8UEk4uwi4/qAG0sIk5/NhbDQ7jA1kOnDMPbhif8V4rE2NhO3BmQWhH1mI
5UaaCchL3+bHt2yRdlXoNVW/K/owjtsflKXXVrlpO/OXAdeWTzZlDCo7UBhUXTFru5lOZpJJpzaE
4ShxOUr+JIcrTJT+xo8odPwKPYXhIWJ6z3XEDDHdeWNGO90PRkdv33NY4vUmUDoYCuEJZzIPz/Tw
XuACnlqs7BX5+qixIo7XfbQo024MStIf/qciZUkhQ8ICRmDQJAKOS9tBKfvHRlxbVikhkyacGJV5
6v3PbJlXVAUjHtWqQRrLqqUT8IAH4CoO85jstoa34iC5f/2jurKHV60+QmiraYuSsajyYK2KN41Y
msxH8Y6txLmp08UYHi+JD6KqyjY9Bpy5mpo0I85vJ+CHuIAKc7rq0zkArQ3TVbk51q6a4GcOLBtZ
Lw7b8gUFvjGhzHqSzKeAo+7ZbeO7Re5Y5+TYkHensOYL8DbnsFy0lW0KGCzDlkL4E2WrRV2oPfdR
p9ybM+r9vO042xI+62UQUTtjrobeMy2sKAbaQvhjrKXjpu8SAjj1KkqYQiJwgztNgTTX9WpBTSOo
ubFEOeqfAiVQmOSDsBO03RIVxUZuUN1ll7kFKToVPAgthF0wLokNa8eRBebD0F1f1emiIrQA+JOR
p3TvxAra1z6yiVumozFzOSkjnpv5JZSoCo73gV1/Dz19nuri5t8waSLWhoQyj1G4EmiXFiNFwMlP
0zvs0kQmOivOxiz36OseWUM3M1GKR+mvdRWeW6n1Nb+7SY2fFPpQNrj3ckh5mJqqnj0eW17aAMAc
mhM0sMUSm34lUq+axuLU4ceqpmwqxGIRVBC5UI5SvmWZyYHd3KrgNIDqLlLyOQ+bii5OXCp1i65K
q+q4G/CEGY8KvL/EznaSpU29i7WmrEDXD7nlMAIdRDZvXcpe/MUe2X2T+zAxKiSSN+dUp8S5OYF7
TaYT+TGsabTimsyV7EXe1bhP0bcWfPmVNTH6WONk6pA1hZ2BLndAcALNtPnT/CKSIchxdvYGDwlM
ab7DfkSg9YKASdDVpVx9HiPKYmthiIrvHlvf+AUhVrBQ+7JPn+Esln+0WIGrzRlL7/+8LDBxyVrq
hyS5Bbjo/lz+pBzbfj1rvh+UB8Itl6dfBZ6dq6hqd/b0J0WKVDfCJwy0t53oacAOLuNe3tyRo8NG
qAsr5BIicZ4QvL9qfBT/FzXl1fCMASOBNmutp54Oigh+QKEEir9ypZXpe6FsxT9yojZgazGWuYVl
vh0zcBdZ5aknXn+oQTN9YocKaSlp2EpTIK1QY7arhk0n7i9+aQLgdXyfN5R2NeExHa9Mr4rOhT3l
nLdoQaWlktaqpy3CwgwFSLDrzUxRmbsnxT8iii7G6yqNCrj0dOiG06MQfLZVarqCHJb1dhLaY/EK
Eu//00WtAaEnBfflZ34mV3RCRzer8NL+hwXR5oeobUILWeWZeiE2HrlQkYMcO/9Wcv+wX7YKLseC
wHVhyDkMLI4bJVb2es1fTsYvDsI/8TZyabJf0bSJ+Fg2Qb9OOU4CsKULg61GX4dubyD+znd07Ysu
gI9dh58sFYsHyhdLT8myMBHhhPE/+xgd+Kgz/0tbIkxXG6X1ZHAScmfga+UdRbuOcHCqckeocVR5
otJKD0JJaZa3SaokxYSa13YvCkjbWxOg3fFIeCxyzYThcDEc2nmxP6F0VrGzLTg5vnxmzb7HmE8k
mWYENkDJHo4i3elkP3J3EF22F/3oAzcufk00i6Hb1+L5Dtf9RR5HkZm/l8bnpE6vhJ/aTi6D3gGC
LoSe58c62px6RTOQX9l1luS+N//AQ5uIf2eGSHM1yeNo6HgsDuGu6oLrh5IqSntRwMw+TNmbyIk0
hBmPxGUXS6vZckQORzCk7YgMPiJfXzDWJgspK95c5J/0S/33VTA8RaZFIvpzZ14VtwBWZb9C0SCX
ubSlKhLo1yOCBi9wwJ4NJ6Ug0XGR4vfTc6Wix1ENMzWULg0ETSlO7l13D+ZLB98Mglb2DdxNi91X
3GJyJf7up535uwFmqkfCk+Bs2HmMlDB+jmKoFS2F6k5nGR322eGFx8Ok77OgZ9oHg3oBKNZDmTyW
uFvxzRzm1UcGEmBlOE8c+Tn77WqkjnPdTefuidZraCLJF29y+gfFmz70rVU7kH5R246J9P+URHTM
CbmMY5HXA+xA/PGMIK7dEs76lFKdk2x+tpFxPuU0VluBbNnHWIamInYflSdrgRz8UAlnXtMeIEGk
7U+M0E8VKnYwsdBzGXpcw9NRjgF5A2g9NowshMqXpqJGrPUPZo6deUdTjnRq2/jFbxaTEEcQWLFB
bPmL9HBO44G2jl68zZi50KFbNBpgmXLt3Dxna+oGgpZHJr6YMScz6n4UgByAku4sXANdxp27nQkc
4mWz9eK4xmOs6ecj5q/60+DGFfRJ4/XFcdTArcfjnTGyDWEHwxC2vdpL1VOFRC0IRmymp1iGhIFS
3Gp0/UrGB+pzJymU0wqsEqybh30blC65a4F1LhRDSx9kMAkvm1iNSEpfjePrHABMRc05Na+gFSog
kC4LaSVENpz55kuPPPHyyho2/vMhY7j9RdrEXp+AAjQJMzLsj9y8ukX69yGFfWl8XrjtswSW6k+N
WAZ6RjdKc9NjxKN2KqG9O15hIaO8phB1vNE8xBRkseh8CcztrQu+jlVuJAdaGwCaf3fsd8/JeSao
mjdDeidfzzycbGsal/8ZdyJISEgGt0NglN5MS5rak3txzug+07Elw5ipBErguxOkyF1oG8WFw0E+
Rb63nT/kaXCLgHE1pWXx7AczMZb3GYOOYrkPhiDEb4qr6S64SCas6CMRUODjRIlepxPi0BQ1bXgQ
hn8eM2xW4Hn2J0Nu4WPUgX3+MYU4gCTXpIk6Dt8VPiKk4XrctCuIBOcjh3DjI+Z/HCvTdyJvhgnT
26JDzqsiS8Vezl4R+mu0zHJipwjZXxeVJjgayq7FplmtJaTVS0WZz4OKnKG+29kKGe+GBR2W3QGR
osupYFubFZ+681Q9oxTx3xr/tC+4J/3EY6vgWFn+qm82fYcaFPjH9wCR7dZnxTDeQyoapqooJsPu
3echQiKTg928xE+dNBaA9GdEXiLI2/FUTQNsBEdrE94aKPCGQW5AbsLRPetyvoub4XEtnCB9tVtt
YERR9uegcierHroRRXv32iSKriedYj9XAbS7sCShnSpULJiWG+4oyv5bvE4+4CEVvhfOMJA9E5iM
3jdxpLgh5mt5P7W5cPcas2Xb421Ee4PZaPfVyGUAlUzWzWoKzwz2ljSDULpnPduEJ8y7JpWmCe9P
yUaxJYDrbVNbfag+vMrWzfrWaSMgmzF0xJtU649UAC7S57NcnhGb66iKr/5lTByrXHtVMdukgmoH
GTGi0UNb8EmYETDJzAstBNd8Y0ZGlFoAWu9GeEjUBxf79hLnlQwZo7kMk6Q+Pb3klrUewA12ntNE
G/q6B2jBwhTH6V60DUDPQC8egBTgo9Sh4XwImuINBAH8jirX6RnsPnJItJ8jTCJePJKxg7tkRYIl
VgKwXR2Pr4eNCJMcuM7KS7BsgC9oiOeQjw/9C2uV7o3fJmGnYAkmmmzRBSimoDQFmF8E3+xM1Dhi
4ALBFJ+LutzwPF6Rmes2bZp8r8fT+ihQ8zvVWfuSdFMyAtoQUue53lcYHSeq4JEq4f4RlAwMd1Ej
0QGYyYW3tDy4f2FU5i7ZPRxtyTOh8MbNPFhDaebgUxB70dImZYF7jmk1WpIWKqPMRENUJ1PedS4C
uPF1PbOtQRNw2CbUu3LZ+mq3lLO62FRZrN9VPqgscBuz5xCW/7b/Z+MOOCA4NocbNEJSSNkdZW8v
wT9aYtz55VvP6YC9ahzQrTe0i4XEQZoN2IEReAoGP6TwGhaKkumvTY+JhWh2kjVfjKBe73FRvTQj
vEw0CQkOUYJQsMhrk+mtqYz4BAJILgA7RP5LP40GwV1fGeWGK0cbTxl/X+/n/r5bh6xZAuwmmn/u
vt1wfjIEcp6oKIqpn1lErf1w+1ek1uswYdlxn5CgVBl5xX2pRiGixs2AdKj74g87FW8IU4/9WMNM
l6lwqhMflg9SeYP4oDmMtNhuOixv9GvZuipDxgNJhbDF8sH0hw3b0sJenVHsvh5RRVeVv6It+npf
KB0FLGlmEKjTN1prsuk7yARD79tFKZ9txMZR20uRiqESLwVKbxuz7DScGlre/3cMDw9QrQF9eeoA
4Pz6iv0vN5hVbGFsBzfUFwFpfF+8RyBzqSeZ2GhbNw/2RPTkV/l5qTMDMo6V9yHxvub17pkVcYua
ftt6F/j/WZtvJUWkZ0WOjtMXe7wUksj17ay3SKQso4domE7v3H5xvBSHFpSezZ6fsaU+D3UleL4O
IOJhPBp4Vfp4nHgMSfyq/hhjmcShIXlA43+4gTxZR/gAZJBQCL6AyGl12SMxs/TpmVV6IsmzHDGE
bgxlOCFrVjIw5SAeU4nbuY5MBUSvE0aLTjZe8f90Q/C7agX244PLfFOMCS262W4sGFxOtG9KNtjT
dzyQUQAasAEforMyrXKMgN1luclX/8eG7PWRD6744uuQrI6wrqGn19GWFCLiAQySoC8S0jehcMIJ
f9jcAsXJRP3U90ng51VadCIzAY4bXhTo42JlJMDVObDhor1JtLaFkS0e3apmD7E8tqfCgVKWPs7w
+tZjgPpdAS6xOF9XW8vLkHb9FJ2w0tGBqDqWBqjq/Z+XLpmKfJQlk4q998wnhxpjW23I+2oE5aCr
6BqSXxOJ2rkxyxbwBvMN8kkeLRBKqK8TG5rsfHbq4HZWLdI8oe181X7GFP80HEEYgiGfWZ6Glp7j
VulB+h/yy/j2K85M5PkF+CQn/mi78Dy1Z7fYTX6qCVgJ8X07jd122e/pqxHv8VuUX5s98G2nGiGP
/Sdbb3x28Uaqlrwxjqroo8X5VQ+HO5u1juc5xMa885JlU1MWhQMf67y5OA0DN0SK8ob066shCPCM
40k8IxRh1lG/Ial+9Mtgo5SKQvhiqdSPZ9uWJyChtaLEzbiza41iSCxxbgJzFjwh4Qz53EXzZ72a
yXSbMIyGebyDkMoTKCkNu/0HNntMYS0ZHoxtuzPZ2zooADguQGCdisBLY0/ij2lVlxaHiZ6IODaj
qcSgCMXILMc70x88K+/81KdIcmtkETgR79FClqGXYyLkafpDkvwXOuLeNdFGVZezzfWWfFEqtzg8
mAgZqciANiATLrWiUqUtx9KSoCvhJbCG3lk8TJb1P+rj6OBEDeA9OjXk9K9cWhukTN8ELqAa0plq
coJB97/ozXQUHPx1kXHprWwYGg2cUKI5Ow7HgTzTwnHceqwyo9UScJjq5cVdQU5NHzCnf1QWyVR2
aXxlB3Xux0cUrzpyWxUO4hQJ4TwHhPrMIHZuF/Q05OXMRLcJ+De+kWf7PQzrOXVr7n71/nm2r4sX
ixvmttMdLv3M1IM5Xwq5+Q2c8PbKeFSQzG7/dmmIH6M5IPmH9gbLguRtocbKl5ZgfZDqltnu3qf5
vrhU5/M0zmYoIsNbFx4WflIbfxFwmKIN2+e0YsLs7fMdPmsbd6Axoy+pReuKwh/Jhxv91NFM2Gcv
zEJ/g5jrbo8r7apq7pFIVBwD4zwKZcC591EA5FsdpOTHxDpU/F2rzplABFm3/Dm2kT2a6nwLJPu5
m5tEUmaCGoLPca2dEKi9MLO28Ars5KBOLA1CeUNDoDk4Buk47qJFWYh+YKI3ujX9pxuilTVXl8eR
mB++Jt6kV+v55Ma97aHVnODl/I6nhbqikybZVMBYZiPa9uYUFF7aRC2nR94cJbbvKu8xh1O1W7Ff
re+gaRnZQbNXQWfGUmyqmycEqoq0k99SzHziWVWuoe56R6tek9bkysZShIPS809aMBo99pBQwrb+
SOfCchWOr8ZHTY+ctuV9uyfghprxmDjeYdt2LF93p9MllH9l3ZmHHwxEqvll+wbk7QOCSqj4af3R
M5AAS53pYer5XhWIORmoAZpZVYIPryasTStDIk60ETcjQPMIJVKVExi7xmwbAosJkNBmQpTLLcN1
CpNxTLBfNB3EWlQN2KWSNuSDD4a/YMGzRUvOBdICQYFeGUY3Aqvzfoyx+GVwjdMhaN1YZTCCkdgc
4gzL2Gbclil0dhiJQC5NoJC9lJsdMuk+fDO/F78baumqZHaXqfCb1ScrR8u7uQo3okUtjrVgzqly
HD+BJJkFNf/Rr7WDqPvS0j9UVOwCaBpSyPTY+JyQHVv9zCQJaYFvwX+JhjeV/CKRNrVqRvBi96pV
oOOpZp+BVcIKiuB4UzKbOh7OYpt3Lu6vrwp7blvV9XmUFwJpHPLFjn27RYEZQhVMEqOawmIBZcNc
nwLV36MN1dV9rtSI9njlbmlIF9kGR/86QHjf7hO1HFADhPbBjlVIgHXLMgKIcZIag7Qt0quDcCSK
LlZWWoZnD3Y+T9uR1hfMNXPpbebLKYBrgIy9p9CzdcWg4rF2Lilmfd5u0ihwW8DTqo9LPa1p7x5+
orBY8FhT4pD0pTssKxowScozlJYg5Xc38tzQrsAxs7vrlUbfj+oyTE1+EGJJb/UuC+jXZqnLCywK
n82nG5dFTODLDHllmqMrwU7W2JjZg1DKObq2tdUmkxZm4Ikn5dbFOU4lJT7+xDF6VhJNaWZNI0dr
srAl54plU/P+3lqZVk06FTC4+5VuElwg6KTo3Urwy7HlsCpe8tlVSI5mw/kxOkQa/mMhDFaOobWk
BLwziHdQGT7PrEMQ/ZfkE2q4bJ3l9YYEo5Vrg6kUa+o0WMVIReJoiTReI9eHPjFeF4JdC3v6WS91
mgE737mhFx/hKZGIyzkVETSxFScLDL0beYmyROZT2t5xFsAiLwc0OOSUkPKLfPaUuALlwOvATenl
zPYwW9XxvLs0U7BSMxoH83g6ng9gUfj9/RRFTCF0yuWsKqpQDn52riwTjJ53Cs8ctEhaGvCl8Ib2
5/1uTND34YqZ6eK+K5gBW97cGn9KDCiNKkCnvqL5fbNF4M1XK3rUvckIRzhl5is6D0A1HoZ4tFs0
1+95W2w1X/+R/UUViJkBR2EEGOTN11ueuyP9EnqdhD04N6rLfJSjERDFwnLOiS4/n2MbZrKxnNhX
KzMZxdCdgeOlLJVREujXFjAc0qfyPWYrdsyDf1y7RPIMN9ya7+IsOm1vt8IijHs3WraAOYkgCCd9
0k0Z5c5Eed76khIz8BBccfsX6A3MjDMJPWrNcgDY11IJj5E7qbKUt2gV0a1oHDgRipPmUvGgdRfz
ahtnGmz6f9Eyn1v7Dln6XEvRkSf/72gTvV0qtsOq1DhyQbpq3H8s+4AmbT/WnuF5b87tTjFqzs3i
cOE2+erozMpWe2a6UNnbrs8x9Unb2HXwdzfWabirnEFSxPkvSr/GE3ad3bniudttE4vH+Cn7s52p
dbbOxHljp2SgarGIWyWH2qpe5dq6Dt+zGkq5VwIUBNq4hlRxecnZxqB8v/VuJYdkNyVXpDpAtAT9
bBy4QLZ4YKgkoBtCh8t8G6iHej+iZsB1k94QViRpkpQdT8W/U3ZQjZqzSPXBZAdDLa/Ol0L3YzJ/
6zjcCvzAfRwQoSmTLDQj1PsK8hxoNV9H1TFsEQw2HJ7vedL80aEisBcYgcZrSrVd2LuYcYioLPhy
3IpAEONUWA+H+PdmzS5RPrcd6ULNUGdoaO7FX2uYTCvPQa7B3hkxOdRaig1vDpMZaHnS47MItTBH
fEC8Q0D8bGtnJqJo8VmXh4EXA2Q+XaVlmouOUpCw5rSoXpedx/eZSPBayynmnBJ944sZvDzyRKMR
c+m75o5Xfn1xHq85zFVYQr9zAtGAwkdNGaJ3q2p9EMTPmrpGenUvcolI8XmEAXY8ubfLuaUqX1Do
bo8UqxBYbg8NTN8dcrwaXZQsaiZKnc3lv1o7JgXxV5l8E19MVGJ0njGnUVdSIurIN+aZuTEidm+C
bac/+furPGm0i5ffiQIEiYtf0VOxs5svn7fohvFgVzYWyazYteBgmF0z2leuqKcVpOllH/4WFsfA
PloeNXdPf2cJPWp3b9Ogk1DvjwCSlGMc9JkmALeErOPYqA5avJzl9+N+PUUdX7AHAsVEZxFaillc
4mR5Hz51lS5ZLjgknw9kQeUuq6L9gyySwHWS+hwSENml5VvEljW4a6e0KiLqvBvP0aHQqUdD91De
xWErt9xcuuKbSf6EAmFqcgqzHZNSEgY7S22FJx9hMSNDyxrZqYvuDqbpFvmhkyyZQPrf4Bcn7TS9
lS8JE1RAgEgv9R/bdu63FnSHcJ3+WrZPej6o7lRPAWqtwvtHXJ2mi77okLON8NizxEFwKJV6c6St
gYC7MJcjYkJ3zP57SiSfxJTzjbzvx/dT12sYe6wwsF6BpDnWKAe+AxErIdvs75142A9/T1BOUszI
9iYI1wwYyIzCyya0KFZzmDE/W2GXNzz9UfKNRyBNainkp8vbxjU06/aXfdIHH4ImY68D+xXvym0I
ZinsfVG2X/OyXSuT1xoGPujloKdqhapWYtefGJxiNi0U6zdc2QHGLy1g4RmQKweVrWo8ABTuMwJy
FLeqrSR1d08h5e69omVqHLCnBjpukK8/PebOpVGUzMzBSbtnR7y7OLvkD4kXBJudECMUpd1IQmZV
eVdM2lxxjP7ZZqVAv10dvvp8qQOkOpZ3ehORB1Kyl80H6GyaCbRuqPhCm4gSfHCLL0bYL9/vWmDR
m/1aoj3IVrTEgZWQAyibZ2gjmpEDko2ernZUcGyMWRWpzDpC2tnSQYRye3R3QawlwuaTsbt/g4rC
yEfoHTTec06ps41Gx4STeERFK8d2g/BBKPcdX8B2wMdln4OB3u3Tp/P+P3dkRB9buj3Od93Wm6YH
CtQhg3G4h22d5uXDywiVyzMd7jKwH+C4m+PDpVGxC6HrDc3ia7M1zvZeYF8CIsaFxkjY02d9MaQv
FwoBTBYxIPdVn5B1OQ/gLyImIM5QK6RQw+CBUEHA5jCoo4UMrET2X2dkxHjAjn3qU1vqTx8mW4Ba
NzPARMIr+FviYqOEKR/HzB++Znut66IzbtSVHcOSYTs+ZYYuip019WgStWI8QfEYvoeIUSZcN97e
ndXrt4innVuBokJe8Ar4v5CUKXCzAeRQujOg8hnLZTAWdXRjCtRyvi1izA1LxH2pRCxrZdGNygjJ
ebIrB7rCXYpQeT9Enn1rioQ+k6EblY700bBWiuswIRGLqDq6DD3pen0qMhU8Lmkcw2Ox5g19Uuc5
mJ+SolK+WxKfmfFzcpVomEgqQNr/I5lnNAdspRPMuvIam2pKDhFJanCCrxSCtMiAT0289rxNS4/6
oyo5UILO/4ljbkGhfZvfJ+S38Dah2QOLz4TAzKMtVTThPMO7gYfIjhJ8HbxpHQfKTDKI3G8NtMKk
KwSNYGkc7JVzvb/qhWeG8Pahy6M3lw0N3rDxME+vc0CHkzViQi5FePQxKQxN5vqFpELtvLqs9Zdn
ao2ImHn2VT4qOodllaA/VatFuuNco/JAtJcV+cyqWOa5d5A/ldHhrpSeffIeMA54r36I0z5yNkw0
exyPsYXXR26pioD5RfHi1qetwDPPCQst6gPHxN00fd8l88Rk68G0f7qrI8Ftl9Qh4D0FhVcr4lKB
MdcH3NpKx4Fka8TgymsRuUwJmwjPXMnCzcESRQxt1MUMp2f0ZueJlY55ofFsih93OrPr34X91Vr3
Q33aOJk/GwvWYGYcMDTBGMR5wDr/3molevTFm0vmj98B5mQFnF3fwlhmVnpsfaY9SuahdPhZhuuO
1zRV/PpkuR9XvtvzU85Q7rhy2yoasfrThkY6UT/qe7fKXKJEGdnkZ+3mTsHL5WhKWsIugAZfLspS
1H4U4i8JICp3cZc1TTmFiPJbXNgg1SRe5k70rYek9bPJeMPIo5DzsvNhsW3OQPf8BRRUWIP0Tm9F
z0HkhSxmOA86t5Tq5XH23fzTpNx8uk9hypMDqDlNs4PRGiBFpsGL2xYt6Vk/Go7OvvJaaU5gBlLp
b1fMBlMcbf8r+N7zIz6K6w6+xTg7yJuhqdFi2Z3kngcj7zUD40FZ/hHTmdEuUgAbZT5K6SC/6aLf
mK5cKNb82aWg81xmBoZufjTLhfDE5khwTOqvrKyO2/jFaGHUEkNWoIDHTy4XQWAf6yXPNw36fIZu
pt8StRLvNoTT6qn4txKuMAzcycaWAYiiCVu5ciFyoIPcfRS+THeFTW3GfmHtwH+3/kbCapRrWigB
nvAUu09VhuaHwgwwr2Qeukawtje68wIbwg1wcMB1rSaOaeuIyZclR/ihpzzRZ3Q8aqlWQfBUOMkm
vwTEDoisRrkvWIFb33n8UuTlniRsQldy4Utu3netK1eUg4CnzWj/14ZNqhZ2KH4unNWI+ZGmB1ms
YuYHhtBsvtzXdCNSUWoyQux2x6CZwll0cXyWSHOYjF4OO683O3zShRTNy+ukrypoU0mKVx8/It5X
ldN0dXJDaQXS1qSH+9G3TAJ6TTzogHZ3knJTlhaWQQlIFzOixvzhO4B5I9WLoMGp3+zDHCk3xjN0
DOVE+QsjJ76giHr9oVB56dmQAXXYXPiV04cC9MOfTqq80Zpn65iguwPuh6RCQeOL3cHgvaCCN1hA
8BwIBRzFNbfk8dxseWT7NnsQPcsrdOS9zhyR7yrhD3px5QykPzRZ95andjHGDniay1BzHSU6yDmT
Hl4vGEcZ+3EExUGbiMoi3mNM9SdhFGOOmzHDajGfSt7FnwLLUKGOXQlBJZ9KbSGLphJnceY+0RQh
eSuRzFXtcKxsyVeDzPp/tARwOC/GB4b8mEFUlonbEXE9e9YIP1KDRNwfWBuUwKWxzm/wqAg/6ndb
Yr7JN1Z3G9YuWyhByNW+GSBrjJk4gNvIP9TU2eub/b1ert2ltpCKe6hmf/P18L4gRSIF8gKgsghT
xWWJXL40KkhHrG7m25JHUI/wVlGy8SxiP6uGvUTxiXSQNdmQJ94/6pjXPaxhiob8UR3q8GX602QV
r2ZXXsqcnFto4JnMjvheH8ZB9urFnqEjkacU0yPDc2nyv8XKF2qC9MVvApxX0Xjxvsu0CR9zuPg6
3Ge856w9GJP5E/+jVvlwaXMqgXMaj26lpQ6MufP/ZgMBQakAnS5gHVqFjKMqCQmXmSwawqh2jMmK
lMRD9cZhTW3UzkrKTvaEru511fJ7b7QM6UgxHCDoWI0V/1QFCkO6V8QRI8h+Ms2BrXezsx57egY2
X+saiEf7yXfuHRRSxPhybo/znEmyi5u1sZSOLshTaR2FuCE5gspDU+2T+I2wfGOTVMaO6Bb3Wm+k
Ku9e20JbTOy4J6d/dsP5PhbOynHwMF3zd1iQ7FQZWKwF21pztk3VqgGx/3LTIkijem2cieXlikUx
DvXu0+EJvPRRs76eSYEYOdwMNzbuargC5NLXuE85WVfwLD8V6tOtWAzLcDpF4YLWl6a9cgZpBLin
EfsHkEUlRXn7eFZ6iG1eAgWC0F9IWOgdnYibT1k8VhhdgEpxeJJFVoqMW+PlKYCGg/NKBrS8TeFE
6vpbN/4KLuWJqnY7voQI+dlH9KZlsJNaOE2Iw9PHo2chOZTH4bPRRoHPfoiwfhyIoSpmTjfWhcHJ
shTXQuc6TTpUSPLPP09Xt0k3zYHsGaB4j6fcUr/24dYdfCfJD2Z+hqY86OR9vLbAt3ndmfjFKoqz
JTfQbKm6sCrO+HJ+VdDz8qiXAtWSfaMZrncNmHDrjwQgteaA1sCybDO+TSwYgTLiZYYKsMzWPbQ7
UVJut63h+PkXjdaCzCneNy5Z8+KLDYSkA/LkHpgFp7prH3jnBbrd4zXFGQLbTptfyBSqAFbTPdHN
FVIOR1ZUlt4DEJUWbz4F7T6ljNzVyy9BESxFPmbe4wyiJHeot8wgqX0ofcIsl9bmzgZBJrbqyqsn
vQ3M6pKIgGLXBHvn1+Kvdedk4MfS1Krg+TDOCr7Mo7lXt35Kp5yv8wlv0UcSWbA9FO26X+bA3Cyi
8kISKushkTSeRIop7br1wuTopgnrCzX29jpwxL5VGUuZdGW1JygrkB2bkGp7rdIqvuC4Y26ZI+je
dDjWv2VYJf3HssrdrKDWap6rq/1Vl2guBIJs2+jUCPauHJO/JzY370Cm7O/xZK9BaBIzU2Lj/upZ
63HILzspa0J0VSO3CPftmBnwecmsQy85UBfl/KClBVEiKiPO7tJZNa9qFl1N+4IBxT1W+0HZSko5
M7dU0jWe2gd1JngGdK6hZqsjjP0nJw/8NO0QWDLKkaS4zD9nc32lv/uYi7JBHwYOB8vuao6XBbfO
+2xTNff6gzyrhbF3ys0cFbDPTlrTbXrMXc+NTRkRaYwaYGn/EFCN3ZIsXkA9vFjJZMUiusij8GSg
khkUy7hDggfZ2z0UcTR+5MzMFjtEp2OkbTYo4OOUVbGWPWzU5pps7mmXYq8N4QzOM0aGG8yHVzg9
GIe1t1pOfgDvoxBcAsmXN3kGAPFKbI2Nz4LHRNsciOe/9Z7eDsNhfgN8Fsd6H5P2YG0GQ+kL/bO5
x1BYjH+RMdFpbXIgWomRSG8c1k9+FCX2dali+DoZp718j1rRF2zTswKf7nMz0yoJtQVV/PyFxekZ
VgXM2XlKNyoCLsr3Po9S+eFiHBF76p5GhpYmcXGCxhoEw670zwOY7pOkIDk5WmqMIs76b94dg5F5
uDIMM746WHVFBLt6P8vpSxabou6TUlXII5HBwUfLWqSeB6OYCUUy4Aoa+aq1Q7ifHhT/85OZuqxs
Gs5MezLiuxDZc1VCgOSsBI/MH4bJ7wk1018ff34+gAmKIrG+DiEXYyMtNrXiWdRroq89BCxHUvmE
DceTW7PzK84yAr3UgcWRCaprSZ84EZpWZQvtdVDo+4nsx4dwGg9gL6se44vrhJJP6wJcXFM9xEds
Vtg1TYmp0rsEuLJuc5v0F3NZcai03IbA/G+PEKfmZjYfSduvS8Ybc5gdWugY3P1/Q4IVWR3MqPTs
zttarUim3rqCxsQC1IdtKgmAs/jp1/txUrBdd7sb46I7LRhTZcq4hnM5YCuzdb8OEKAt+VasREjC
kMYwWQHVql4qkkock7YAbmYFoNEIrGIwL5eq6oX2VIvUrWpvkuOufJs0M738I4sMxfDiUzYyDJM6
FPFeh3+3AQp60JRQJMitJBpEotc7rXhwF0bHlXUtmVnsv1H3/k7OYYEjB/QmnqtG14bkhBBH0bNw
abRS0+49aHZxxderjYsq4wVX5tlwT1OXge7Z55Dk1Dv2HdYYCbD3TXwE45BJh7+gNgdmMYR5rN8G
mNff+hEc0YBkfr5BWOkQtwTkAd8TjK7jYQ6u9oiZA8jIoJhB2QBRTptDIi0bWeSKHnJgDLtJYWx1
vj+ggMXUJu5Eb0hsxq2oMMTvLGLehznCMERL77QO173ER9FcazYmsTG6Q18CBLQHhvtPMUExwX4X
fPB6kw1Am8AKDoAj8NNGqWczI3/JyH4xDaXhFPW0AD2HEV2JjPWF2EmNHrBiIHpsecCb94DbDfjh
6vwpZ++7riMbg3//XIZ2CK1lH1lDe7Vd0f4RcPAhkyZSBMx64xDdQZdvAKx+esF3fTGpzYpWEwgq
we0dEpQRE/goYZaAChSi1Fe5DpzHQRWir11U+bDu85dmeQVPx8g2+91a7Le+CBuHZd8QX0FPoz0e
UUtuoE/88+WCnzyL1FSUs2Qk38icpebpyoZtDEOPtl3X1zP/AP/BS/baHTTHUvwv6b33QO3HOrL+
8Vyu9Olv1KY8P4L78CP8z1BjnMz7XffXltC6/HRRKYCaezO6FLxYlhhfGePizC0tCKr8s18wbVNj
tjfRlNGL5edX16oovvMY0SYE3MPiT7beemdB9IVJHbz1t/h+ctmphMhT++a3taJUaT1aY3cJ9fGb
NMxhPEpht0aM7KaZEhEWeTriiDqV6He6dwGt1gKFi3QvibBMEK5y+yhSuv2mw3nOPWHdmezmvWhT
vRynkIMbh+GayvlFNBWU+wO9XwnHsNhpF9O0DmKn5vbyrDHKDaLybdePk1ehp8GE6r8A/HHLFAQY
UP0vH8s03H39ADmbBDGbK/Ef+DvilrI5Xp2lqHhAfu0MzwQqFQ8Th0nStPHrQNTcTZYNWmyBosZB
LVDc4Y6SI0jWQSy3MVQIQctWlr0j2ywjsd1Ggr2GwK/Y/qhiHPLq5EJE+3MsemXj740cnc/6TpjF
t3xoK7AmEYs0ogYNrKi/XEufkbmlOvo06CVDRD60qWLA29/sFGlukS8Soa28kzaTT/W5TAc6YCCo
Kw7NUd6J1nfqoDv0BR/4/I55djJdWydrbFjrgZQ0owXb4elJuuUTIFvGQ9udZd8L/FcdiJCgb93b
yOgqOtpuBiclUKgk2ho/bNG0JU3bGqWuC7DL8bCXzCgwhTN+WCZnvL9Yvb5nJ/E/9NylENDiAkyY
cxcnvoZv3mfOsXqNkZZ26O0LBtewAzOEPe8ffTTfcIZHLB6odlzRxWEYnZeHm5aX+4tTI4IqSGyn
qhFe5JVWvSRCjTSOyez0tRHXez2vwvsABvq1xVbTC86sB7bgE+Uy5vXHhPuWKTBzOJEdDgCnEG7l
lbKIOuhgJpp+YZ8xQHvwi05npYSslH9uyn99Wby2NCJ9FCo/AUhArskwo9GmYbh+gs2fQ5QuRelI
RgeGbvDUbrStrVmnvuvdWrQxcG1Dn2qrBGEeBOGZdFXu69JXW3EuTzonP1PuNS8giyN2k7qRuhMD
aBIyDbHwsR3TbxkNm2OgH5S7FCqHQbVZqdfdW10VUTjVmE05xtMdJRiHYj5VvaXTKGEYjKRKlKmu
4c0xwDCR+pTDjzSSlX7I9KMrmRSw1cAWuNkksFB8NqBXKGcMhrcfETpfxzz2p9tM+GbdQXyKGveR
Gj1yr3XH+9nR2/m/VeLrArGL5BBKHGJ0Xjn01isMgXWhpbuQBGR485Rz5RZmWi6aw2J4uiogUUkR
/Rh0su4oDsBlyrm4rZ8y9Ty/84ohigZRKDIjzsiQHfF/4IS3UI0SrY9kyLgK8fqxPAB7ENx1l565
NDaUrs0dVqVHSLWdguvawdqbiUDCCNoagLNpT9eGAqD6f4wDe561Qrog7BnEtUMOCX/wvHkk4Lqs
H2X6bqwRJ59H8H3t8IeAmlS+VyiWzCuJaRt+bu9EOT88SOroyBR6KtjZWxWMhmVlkEQi5d7mvCx8
CpbR3MYHhcXTIjgCdslCUOPWZkKzLolY4YLBOeTXWWqAJWOuuvq1SLktTaz4MPfM3ItWgPo1Axfc
dXO7PQeY/rL6ihdHmJDyh2DzS61ebG+yq8kVz9S0Phi+dPnkbewqTpWcAqtq1qPSjsek2ZqHk4CH
7RAGaw88vEZBQbPmEvbqWKXb5DHUYn1VVPAogt+WBU6WWOelcliDPhftqCh/Lxek4Rq9uQPZP3za
RH3tZHnBJTGrYBbOwRxNTEOV/84ZH/XuRNoJKzww5wKHifQInvQMlh1hWPVpE8DGEsGE4vDn9Yzd
j+KVOUAySuIbzfpW7E+kvRthDefCYywat6CMMLXA42dxpPqxx27f0gmFH1mGdkoTSlDJidm1qE2a
EEFXqPI/9bu2E0qNl3CERoMiOM1L+LPxkIHqQZoCWdojWTRNF+FV2x3jxuIoKkNiLZPIvLlnx1Qy
ASycdZ3Y0paagcjpSZQFjIuYcGg50zIWoyvVHM3yYEOCFWm+40q8l1JijjZ56rTM5BHgKXQDQV9G
PtGExeqDPbX5i3vmAJ+ssIibzdn1ae41j9jKSiUuU3CSJjgSYzgSjG8ipa27Ue2aejN9wPRl+Kxq
RtVQm0urTuxOc26jN7PObN87yBix8BiCbcGSrJS83OQwMRJSqA25EotCNDkAWoM6jNBxa5bA92dH
Bu0iewKNlyoMAgQzV3JUMuEo/NuAtfKnPmaroYai2hH0ECEY6/kCwnLcBzakFM9+STPiT+X50vnp
Px2vB/8rlDnGBVWkoSmIt0O+WfOAKTqj/yrpLRungXUgeqPs2ZNGGK9A1lF49HqyzZCFXPTymYfh
UCg4ksq3sB/DYOIa9yVnxIDeZ8TpWTqbHD4vnN+lPM7Z+rBmCVaKf1z4zcFh8knC4ixJxPzmDJqJ
c4Wi1PX3RD62nOdgIww1BP4K6LRC6dhXBWm2iypa74nCx+kDHxUyHdBTU0eGPNi4fIjlqbW4GSo5
jy7J8i1sRTIRhAUtjQq25IUwVGspHMCRHioFeeZ4P8ciluN9wdgWux+MdTpJmk2UMTiFnRm5K/76
4oukD8fLjcGg4ex4O0vTc4dhWnxDuEoZ23aR1NWSR78lwE8dTsk2n2VnWyWiRmZVK1Pmj7KUM9tw
0suI8nkxaakJu2roQGG2HhnuCAQSanuNdUBEA0NNdfm8e5UjHwR3cUNK6/P5SZQARLbaBCpw5W7G
98vX2Z4qvUPF5zbmoxRUPo2tcNik345pR1vaXRkXGJRDLrqUQLGCjYeaUV+2Mnz2wbb/xk3tnLAW
iaKlaBgZIDSgoOwf5a1st0sj7H+ywFmwv8UagOCX5gRHbjc0itZMZ8U9SPJjutUfj2nZnrQEyZ+C
Kl4+uqg3vmjx61oH5p9RcPk0Y7YtQDxGvi2uFAB026x0+CSF14wTFyQ1DhR7bnZGvGN0eNZPdVe8
+KlEGLx0QtMmXhYEN0EOprgoSm1OXtc0S9mHVs6b8DAFDQ0jbK+kTgxF7ze5P+eq//thBiegfZI+
jb5kRjuTOLyLvaJfCe1ghSa2NJKVGQvlYBcNYrvj5oVx62981APPE1/xXDYk6zM0ll4FAv4GKnfC
qbg/yoIuErb6bFWfOl59OhHr8F5SMPELzKvEBDbuehaQUmJ3hRZF7ZgfisOATN2VWgaMoOHBtAHx
QWairMAomU5GVYGLorP+II2i3lDD0nOvLlqupZOloEVAgS3o97f+9NJtfduaqBf62AcMpA9l41Us
04M0HpDPzqBSl0D9WW2rKZHZeN7l5qh8A3WJgsXXkAY3okcNKxlRWNB/PQpKttG2M9DcvbozPpIP
YRKQr6M6WK8ir8Hc+N2k6sZ0ENKevnSj40fWS96TmCbAlZKXavilMwDEqn5FbqiRwwhBogZrdfFk
PCMmZxzsX4UdjXT/0TUoqDmMtRIA2YCebY7xId/08HBl22gBc2KIPemHJIa9mLrMOaA/WAFFzJhS
NC12Rt2ES/HGr8nR9dr3GVed2e3l+kIRAuSyiZ8PDjHhshDcZ9j0EROnwR7FQ+D9pi8Oa26+hK+f
gnoxmFUcBQ+sLH/wyLH6Hgrfsv+lJ+mcub5xr45eDwdLmh56+SE1F+BNtTYsRZ5pMCrNhJbKJrOf
QVMcqLEpoN6F2F88fvB5x7EM/5w/yDEKMTXH9LiJsioxDWp6EQkzVbn97W+mrjyx82Tr1LXQdR6l
rqHL8Ile9CdHVnonl/e1PbvgafSUBrdBnYRraGiX+ZR8xQ7tr7psUCXztlUn9Ds37skjFc08BhqJ
h60MzjN9aBLl/JlAZTfIPqf6coV1zKhjA41ZWGfekHOnzzyNxQL3N2AaCwVODG+Jyz+eta//ciJh
55NzItMJ0b6Ya43YH+ZmDhgQWr0MXXE6BzUDj0MswbRD0gDxZFvMmg0+Z2RHDAtONO8H6qKhnEMG
nhsDnocNIq35RYgWqqXsSxbggWZeqBM2UmFRvPCX/aQFaogQfUMQ3xs2My30VEDy550BXNzjBaHH
WRUVJCkAf3dUzDqG4dnYhq1yUZ/iWN04kbyzKpm5s2jXYbewSTW3ccF3zRI+Tqgqalo/XHvHuftN
KxcjtbRWGvhBqSlZIl154owN3Pk4tUC9Rt1Wy0RmjbUeMIjSkuMX32LPFg+pMVYv9WxHaeCWUuMH
fzbEEZeZkaL2uoh43iAwaDL70D9fzUVkorKP+gHG2NALT3tGQHqSJXRgdatbhWdpBh5wyIXHC2f5
03+In5NvNavr8cIoPQldoOSFcSUVoCj/pcfKkKtrzYnZ630i9fxMqm1TqHeHPiOB9nOi7kiKGrFo
i4gVU5QS9sTL/rji6Bqy2D/QqM/Q+gUzIPaaDdSMwPuCmuL4yImps976TFBbPb9S4YQ2RiTAVRFC
2wKvZHl8pzDrvQGW0ueMilxiRlMlH8V+QXRPz+W/1bLw8KbNJOfy1IuZTuirel746lecx3UvWiad
0jmoRvA72Eqa715VaZ2Rlp5gXzLZv3GjbdebJOCoACz+MWaOCEb6GYSTCze6BBmVzL9969q3fmzr
4cjx0EflObOZOcFr9d1YhP8ySGrCyuuQ/N5U8maB6WYT5NKJhVGMMlEQ9Rq0utHxwF4HJt0dvlrs
jbnY47EaqVfbY1YSeepLuoALtdrSVcWzhNbYgSs0PHcOLjOb6i40iXeWIpyUZHiwDN7A97HwNLJ8
HiaYmifaEw0pAxfQ8huzVMn7BavgPpuTlSwGQr1ed5BVZlT2ynSUsVLzebMD0jD7F2WCsrN3G6vL
TJM4YbdEMUADiBGQMveYeu+yEfCeWvvfx0MNgTV6mZLiUrqZtv5NpYVCrXshdfHzRMen2yiPps1g
1paBEUJkddvTsahdaL5TTQPMdh462m8C3yDYyTvc22SbACIZpmLDNp1VDqM6XRzPRevA3PcSr/Y/
HL1/5fkSKVDkC+Xvr+Ptki9Sr44qlUaiiKd7GrWkZtrVdmB3R842Jbnbtvd03QLkBmcxYB9RFErt
2Jdo2vxQ9TZx/fgv26844laM0eTWm80BJ0wJzotkKhaBgVSb6yF/zU/YOJxpETetx3qtxqJKV7I7
DhLWzoPQhaGxZmuwiy6pOXMhj5VFgZGFgMQSMLafAx+/pqvJZ2X5lLUe38wSqBVqoE5W/kSeNsdE
V9HxKEDqpQ2PQBgsMN9RsFWiUrG97uQ28ctwN1GPHCXOVWXV8Qcw+9D+uEpq2gPC8XoC+oUG/Z4w
fN6oc8wmH9gNakD3JymWsteV6ac649pW0Gjt6HyBzG4wWGcjxq7mHpItQTcnesf+McV4PhbXFZZs
5lHVrLJoSoxrgZHxPOnBrRzVzMnAvRiDE1eZWanpMVx9v30nAnZ3wZynRlGWkzhFdD+B10BY8PK9
7YEaDAGcAshwhoLkueSMbZLhiyE9/jbi1WzT/saBqPE5VyK+MluqArzrPMzzoVI0COGrbWmS9hhC
f9IHV0+AXJSkyXaSSdpNTJrXIXOuOkuxAKLvpi3LQj3OQDYwD1q8fAdcOrXH/3LBPHhJ9JVXACjo
jquAcqPoXwIswOe0GjywMJfl74ed8peL4fkLqgZ55dE/UBUp833nR6EXcB6cbWgQdij6twPbytAH
0k1qAVpgz57ZggymLGNX/pDons1A3peTufQH8+bRo0Ysmu8LrdWhSyRZ4PLrguNSqiJexll8Y8r4
QqFELI6LaS3NT1CckpKqmdIVdnaJz6hYqvGICucSjyXRe9BxKsQ8jKD3mZueYPceC+x27hLqFiHJ
+gL+IvMebdCTj9jjhnylLTV2KXDs+DXDpfl8iCfpybmKMXSCzEzBolwV9mYNHzgHlBEGTSN26w9+
GYvrYPhWFjGcH45nzwaGUX+nxjcgW0J4QdSX3u9hjeEBQfJpZbv4WHUK/dM8YHQWgdpju642OMaC
ehTnWbFNroGErKkgSj3vZBy1K7YiXOlnbf737VIXxfU3k5DQfNwKcHjzJagnojYGDDz5Bn5BT0nI
ZuZHYPxxt9vRMe3NZCbcsLJYeTXihBmjuXod11Q0jh554AxNAcp7532ZJBVdU9/AD5JW5mrVFXOU
OydwBpV9ON6ua5eyF8mccRrXgRfegJ2sfB6jzngMxx56y53uwaj9f+bkpx8LLSdsRy9qfrRiqRRd
YDdu/UHETMoN5oErQlK+mmp8VvvD21d9BBPc0RK4gp+ERWPx3Y2ltutGk1BST1VApFxTzO6yix8s
jYF9qinzoCGIpD9bpMUStJ0CRf3CcuhJNjms0aZIB315yAs90Q21sJad5DQfrnkUs+Dp8jZhfJrd
Wu74alqagbsEbBVyOkGEx14JjooAFYJkSqDIJSX9Fw6YoLpFbzT9n9txmqTbHhdenMDbrDrWrWuB
JMG2gYm+ZdoK0UONIyIDX8NVNGVcH9wt5y2NqHQ7wRFSr75N1UxxB97QIf3SVAu+ZLHjklyubzEw
LFWjsB9ESf8K17FUVOcKZTkd54Xmp6PPb0yuaKveLzANIMXoNGroy4KO/WwFd1DAjxyfGsepD8Zs
R3ityV7q7vN2fshMoniYiSteLp+PkgDq46PfZHWFlyHnQ/iDxbcBV0LDAdt0tQjftnf4K7L3UDCE
yokNsvGTfVt8kjXSsGorF2IAYEiLVbVMlZJWoKegfOhCxMab2V6J41jzD1WCu5IjazHa+gCfWu13
BYOosP/C+7Sh22vHsgssbAwOEuYV2tuppo274b5lGsUQLqEv+tWPAnKZHNcjLeHF6oC0+md03mvw
3BZcgGyHp3JRBfE7w7twia9yB5a64iooQA6LDUOGVUqaZFP9Kk44PmvqXItWU9UGjxvcrf9lLu5k
9nlTTes8YaBin4GCnnEJdIRvHsF8IMtYmtrtQclOV5IKJMRCaGfCmq5/sEahwabSPQQsk8qMs31v
373V9f3OG2/AGZqYL9OIzPy97fM/vXk+ygfpRONa1ZM8agiUPfqRai3XGmBMTi9Y3OHlGOSNkpws
ANZYVS5O512F+xMTZbzYO0iyfJfDkDrwDUOuDxFUFhtS7SgapnlCvLZJahQ3wYwpKAT2rRXYBT6v
FyRO9v+rsvnFqwNt9FonaXQEnhbp+Hsrd5qszIW1UBGqsuTWlqtiZweS6iWXXwyyGf7QzA1ek1pe
9ozie7sMXcjB8yxJ+Zi9oHmpToPKlmRNI7Zo4bogOe2BVyxjs+fXmM5vNdZ73gLIf4kCclFc+/yU
Xm61nfVKrGtikq88dl1UTOv7Hw2hlCJhq07dYxIG7RJyWP0CbSzoeYZHfvO6b8OcuavV1VkmhTv0
BbRUW3ZxAz11fI4torNtErOb/zGcp3Y4Xnoie391v8uJ1QE61fE7PO+KmhwLqkDVJ9nkA4xxqe9K
VZHcFwoHRobJSP3oBm2rfMOzgEX38rGqVKOpG4uSGfTps69bUpNIVeRbwaNg5cUeBDpdD/eVZ1q1
khIPQvCiRU3rhJyTb9WUQ+2BbV9TZ/PBpsH5InqMuWADf9SH1bDgUi9LGUhSJ7be00Qg3rEzJloa
6phd9GytS8hr8c9KdBlAaMjkefy7Ti4EJPl+2oL3UpmhbTXrW8JGn5R8aYsdUuXgM813LfE19sEz
MDQYfjoPXpSWmDVB/HjZGqq7cuCVBwojCz7P8U62mNLlIlujC67c3t/Jr/uRmQQRCtxTvwGfeQmn
3PT2lnvgkLPhfuyzhHNeu/4M7vyBgCN7zltP0lwhhKMeSPUejvbXI90m7k+xn0t9b7+rPtbcSjqW
u2YgHdZvkUdX3Gt3mZ73B9NnbAvLJX5p0jB+ocXPdyuj8bkI0Yy8VrUOYOEFAvK8gbx8zRXo+fZ5
9Ov9kSynAtId7Ff0CzJK7vqCpsfbuQpAbk6knQrLp18bsO2Jy14XuUndIAYiwRncCXT6HTDObZA3
YirWTUuJMs/x1BKlPaqGHWoCgASHtMXJIcHlFWOjAKlkLxNUBkkGhIMghBVseqKVvd+Oqv3j692g
Sj12Umdgqk6yAgtkaM8Wx0/K9pnO7s7im56msJg6v13GRVP36m2zmjIaXUS5VEOKz+wyyCX9cxBJ
REwunYmDbnqWHKBZDBujRjVgQQShk7sISxO/6TInuOdM/EAyd5WaxYkiSDYN4Sv6/onfPcSiixSS
P2JBJ6k1nCJA0iHt0YTm0npncXFdGaC+vmxqCEatGANCSJwaczzrQizluuNnnMH07csGJ7VOYAsO
5SqkTqbz80p5TJF5UFTNGQ2GzRw7oX+k5TCgAWz/tiilEjUWPWeQXiQ9ldp1suEunyWZe6wmBj3E
XqP601fYLl5I//04O+AbU10mqmZk1oeqFOcl11oMPWi4bhT9MoLDn7VcWRrViAf7J8A93+dJ+6bC
roOGncunKpGb1piFHYTsJEW8NCT19DIH6LG+fD9r5QaDmrxx/3mSWmYirtuPHlAM0zaCPc1wBxSd
t/zIx2CQ+J8Ya+O5Y/r/xrbPUUoNqwOYYxnynlDrA9gdKdrLRafGar+khHcsHKxhJi7lqd9kI68U
r3mEW4sVvUJ6qDujA0m4sLl/N9G48ofGEhdk1oQGmwdHWlqkFtQY+v7nflX9l8yezWNGN7FPMuB1
KNQC0jxBwUyt+99/FsvsDHo5r83jKRYAFdkQM+vhFNWBklxsjBYqfSCKjMM2gVZI/S5I4PJ7UYs6
EqNiiwCtB8BCuLO3+tP3eljmHsUCXY7P5G25wb/Et+p38TLQ3o6d4AP8ysQAb0aFWoJyQy9ZVR4Q
KD4H8kgwg5LZOm7ta62xFErP8Di7xKiIcsOmVjCSMa3PLvKrynN94M7GdGV47qoUWLszuUq9ZrFj
6A5SGcgUdfOrnl34240H/T0iFjrZ92hymuQ30YpbjXeY58IOKRFla2jvzihO6KBmC201KeVU7Cn5
g8v/RPhKSnO4xFIbHByAfNONFTSYPdZgu34abXz7V7ep5gWKRJAH1tlMFQp225ekHdg0ZG3Wkqho
xpv44X4+0Vgh55OVqkrdnhWT5soLcHPEr22bNjV0JmHlXDoQvL/x7xbht2IJUC1FsPJwKFqd35Rk
BXeg1t1eZQvSXyio0pBQyXIeHbN5ThKl+1IEwp1IYSlJWPDcB4Hr9oiJrv2FAHBmZ4TYvKCciYvY
Yn2Hqz9FKdUvufI560DG6iBo/J4iByQa7LbS/eFDMbtU70w7Wd38oeI4azjWLtpnGFeSWQqZipAB
pl6LQuMi4meoHer8cUJGEsACD4hg9qeuk+aae41gGOebfLaUyyqZ7N1qmnOhaoakpAxDu7veFUUe
u4n8oyET9FEOd2muuNweBcR2GidjjJDrcLVO8vF4N5uyALSOxETCpyvxvMUD56bsj4hlgZGPE/hH
XAorj1+fk6mlvGIvlAoYJ5/9Wu4I+rJoqBlQiU+1ekyWt+oWiswoefjv86E1S7KHVmk5h07pPtkq
c+GrEKmZpFVhJgY2CsLWRHqTvzGzDfvUpcGkmLbRFhuaUMj1El6dvBWRiwUSY+4WkbGKivo1Wvcw
t221ncrWd0TQ+yBJ2jJ94Ypsk+cz3nNdu+vaQjn7DV2Cr57wgpLjq9vRHtgBUOawVrWhDGTlTE0p
DToS/AuOPeXFgXu+PNjojonrYUq0VXxz0V969IIteBe0DMyVgOBMusqART4T3gf+85nm6p3IKJ2I
x+u4my7/P8303MHfEJy64avxYgD5Ctq7FXuRukkYJnLjaeBbel0fISr8KjDb4vQl4KPLeffjMGKM
USrk40Lkp7pj9OlkFKbRLkRIBUecV8nl+I1ZHN1kPs74kbtUxZ47+dEXtSQ40MyWPfbp45AQEuj8
IGq8lUZW21g93ZkDUR7Oae+lAt+/MwCFyP+IH6Drbt11PYZ+AnrzZBbcO0HtjTfCdBybdefwQMSS
96w/BR3Ptyj9S4zqtr3HDbd6FVbCQK8pk6Ldy8FfCi+cXjiVlX6TjnoIhYXBJL9JpRL6372xUnLq
3/IdekFboPsEKQYLUNhOMQ+5LFwFChlvklAPsnllL1Ls378sGV86tGm9x9lnt6CHUIHXbB/Mn89N
ZItMa7U/Yusd/W9kDLhnaO+5eq8U3pxmntG/zir2cz1unzF4w9hkdvRQixlSG0h9TiSoQmVHI1DS
saFtWr3+I+q6p1+QXyEc6Ekt027jbMWdXbtBuvGRPybx6CFae9ipcPpn3P/4EOjb6oXkhbh8PAiy
t5cSECEeGZmHFSkhZaCriRhfM7iqveK5bTjwp2R2M5we3vneOAEtVMWxqxgc4OZW92trOuC437iW
Zf37NY8rqZBBwcgM43W9tBmmgeBtDCGhOL1HM7N1MAQHcm97S33w0qbT/drBSSHsyY0ZvPwy3136
0nl6S6EYqgPynISMC95SXYo32O+HJi85FEV3ioZYH7RVKf41Ir/kk9tq0vCjty7CkM0EvrwIX2++
xSVp3U7TUBuJ+wKyF749kn/lVwZ1MXTvH2HK+WX42REe+44kveQJPwWOInKDdUUi4kzC7RiHkipl
MPu3XbiPBnCqWjSIREQ4icfGqJPEJJQElSdTO9tn0GR7OV7GarvyIVmmayfrlI7bB1co/gWd+Pf/
qYDenU4up8EaZpZATfpw2O4udjk9LpX4E9kMGqAMthU90TzvrBP307aEjESxHrehpbm7ZEsi25J0
f6D60YBQ3Neut6DdGdi6vqgxLuqjttiMyDUZY2SjgIx9gfT3krjIPELM97sCTCgq6NT7JcNK/Kis
T8TlzShrTMXWv2GP4Kj0MnXiC+E8lGDb09Fs3VUoXp3/70DdGMoYQqA3fr6cQthUWMLE2XIG7Emg
viC7pYaDuW+QWAgVH5NHUgwhvfo0MD9tumqMireCCBaI9qTZC6GoH+S8zAnrjImp9eaN8gy4ibiV
p+86Y8IHMa0Egbbq8AP3Tm2PR9xKuQwSCjqYBrZKQLgOV1fiMpAAZguTJMYJ06KX+/S9mSt+Z04F
dR+1ebLNMZLboYGq1PyVvsCAd9jPAg9h5xXKQM+9pGTlKXwr2ePhdwC+vh5IiQ6FVu7Tb8H7cYD9
BdtBL9+WRS/NPW8/NJhS3Gv2y/jFwr/DXWMuAD0MkYkvqRjBMkGqadcFdTwbn5cd8U+W3mXxKt1/
N+mv2qKQx5XjUEhQmQxS4bflTGUE1Xw8+iplDCcAkHx1wmlb5p09CZMDA/IXnU2T+yB0U8nuOPh4
41M7zbNc2J11qspe/5HzpY23VrybH9fARPH2wSD+jG/0mZB7n0NJ6MhKUXNS5cEg/fgFhx9Ydj3d
4SIKgKKCSliKcoz1F3f+QpT99UTwcKpoK+bke9l4oI2bQG7kPFdNAqTdrBck4lwckZuNUnxeVTi2
TvUtbsSKPYhd436Pn9foICRfGyIr68CH3DO8fzXqnguXLdWFEyyQGHil8MJ05a7+jhUBRUUQkDdc
Ysm9965UzeAvRZA3ls3NLnqMi5gtmdK4auTDFAWaOfZLgbXdH0K34IUeExNPRdVqt1tfmV8wejZU
dZLlVMob650RIh8G94L30nKWKiUzMQ0CA4wuWyCaCGj+CxUNmF9+nFy/TAK0qQy6nzoVqMsFniru
Q5TIFPdlZ3c7JcmqAPpf6tcUfjoWtYmKz6W99PJTBFME2LMyiQBA8NERtzjNRiOiiGCLqEIOZ3nr
997iEKXavmn4lxeLnmDtEOyxcUjb8TorXFZZL6PoJHMB684XZm/+s8cSpvoP+vBoNLKEkxuJHrAc
2WbC/rs90z4plkL2z34wTCJ+q7Oh4NsRybb/am4Vfscb9eOkcdr2VFOU/iQLtm8Sd6FIlCrJUqac
cjwM+4ISwM0Fp8E6jgzqrwaBPCKgdwICHiSzxJc002k+HH25+caQzv05ATFmIi4hFXAC03hInuKe
MJeCSaoEJtp26Da3krwQ2YnH9peOxKYDloCdnD4KWseQlM3hFLTwmWAIow2Pe//7b0ak2nkKLQVJ
DagZw2r41nS3ioqa/0WK/u/rJ316Fvu6EJT24hWles5cdY9Gv7SgJTRHJynHttLbsQSPShuXntGZ
EFrVk7C8f3FHmw51FQtM7s7OvTaxa1FiPrEH9Y9+s9VAbOtrolWaL7m4J7mYkdoeGrKiZdmSAyfA
lMWh/RAl9HvxdIFnVdIjwm25zBAHIHP7I/F118dm9Fh0hom5p/2pSD4LlEbg68ryNwEEjjTKbfGy
4RJhSy+RpH0LzdOUGtieQ0Iintxstf/AUCYcHH9TS5YrTlu1iowxzSfdrrLOsmEb7iXa3jpFzz+7
ZmCa5oTqrqwrKfiHE7O5egn0StozpGxwsXas35FJ5Dm4uK6qAHcJQf+0MYm7wajm6df5RHx+KenM
GTA7Q0hr3lO6vL/EEf7gyNPgiBK49SaERz6QhCrWBIWPA+OpHPbcWulfn3Zy2jIlnPleKCclRXHY
MdcOtU34fjiGgDHTEBdwBMKljcoOB9pvKKB8IqjVRBmiTvN3jXEUh+UhJi/rFHuc70iJ45RChZMy
F7KvqtUvEu8lQnCMPXVcALWO6au0E1/dw0OxwaEQL6Qs4XAT9KZj0Qr7AKrP/g8uI4IQJhmYzxPi
c5C6cXk1ffTXreoCGNM6gPpYel2sXca/J/jk4ISakKorntr/UxO78OInRxhIF2kgx3bVqIHXpusn
m4o92n0gsdlYPsXsheyzTgXMyFAPAmASdM1lbXdsVaUUg/L15GU2+EZZ7MKHLZbohyQvZoYvkAdh
jA2+7RyDDn16muiIk8aTRY6SI5QXWm9CTDMJktGcX5R9HehTuktMEjYbk3EwOuW7fcKeXfjykncF
Swm2i1zEE/2Uto7KzPHYdNpNowqMa1lYmr5V1V6TP56KrF5ESu6h1Og9Cv5BliiAjn+BdjivJ92U
xD3GLXG7nfNZCeqaTnP+h5YGQDdXqXXhQf5JYBKucJzSIWR7w0dgJlR4gImVPGKfBS4ElzKhe5Ci
QD0oeM2eooUKZK3Wxu0tynNEF10HUhzUnWWPq7cOMZzW08GudYW/bAjjl7avdTuNXHOh1fKmy4PX
2Z5kaZLcQqq8ai5OS53aQVV/xsxE+6Gswe1AVi9D5+9CzS3f/751MzOlOeN+6rwpmYFtXADyvJTN
N0Qa6e669zUvO4+kgDVeJjqCMaWt8YOUzfE84I356EG6Ha4L8B+0gqVvM8SkDZhXF33Qs1DQCsJq
n7HBhLq2SUPswkW12o1YWDea8KnucPU05fFWmH+wdBW9Vy6y+J75is55T7GQZZi15X/ZtzgQvxK3
HNIRdO1C2CmpW6Npg4eN/g7uwu+Gcu3CyxfvZhhBtV+EL3HVX1H3iNCQRLr+lYLAyWXbcoIWwI9l
J8xKZNQja/uB4gCgOGhv1Ht9/FY0lVPuzTA8FpDbHhrAZyxS4kim6YOf9+YZnhY0py2hL5VqSQKK
gtus9fY0OR2LuqGfRvh6XOaN/XegQvR84KdDVe1/UKyUDThmFb8HvXjpwZM/Y3JjuhRJCJepyQrc
IJjRBiVOoeg5iVXBZBrT1eT5z+dCSbCGUx64FOiBrQcXa9RwzRmNRv4Qfi/ud3r12my6lYvgyOg7
9BUfvARXXkhKkUzWENsAfuZFv7QKRZjSw28V3hw6OQsLA8SmfF8RNQw5ogHD6IaSXEDBg91fHU6K
XZykrzoVl4MOBqUYT+Vy4jV1Ew6XXGQE+RdbVLtZTlaY25ONxaxPIsPOLp0mJ4zv8r4mghhNuGjV
vDY73qzjL27d98rblNQaCmt0Z6SDkBn0PJnrenN82Eo9eg6HdF+ymYg0GqOmvBRHl2RFvVV6mx/P
u1bolCh2pRmVqkYQs9abYPDCLtXFR4DP4eK+W0YeFnDkBogiSjpIa55MFZvyE+H306YZEe2UW6Lc
ky3EcCb26bXpEUng+Rm6q9XVaoys+dVdkuhO9Kgd3u500HPsDEl2ShbDb4KeBzNyA3DJEGWicNbf
haICYyUa6L4M+CRHVETjYHU0x4T1/E7mEzCKkK4EtzAcFxMn3ro7XXa6imzAn/Fl3YEJg/n0u6wm
OBcDYo6kI/PfJoTNTQnoU2Rl1j1S/A+EUXfvRpdfD0DdJqpm0vjcgBaXcTQeSoCOXDApN0FIjC6/
cXj1AEB2NCvGpE6MLxyUPT0c162jSFfCqmBipBo80J0PMj3L67oIITJ6myOHmjV++9ab9B9y/yWV
OSCNSxgmdFC5bDGca+xDFWAU9Ysp96gJMwpNAVLCoZ6M2E+XX+O9Tfz5KQj7CfTfgKsG9dYm0a80
RWApBK6tTJyBiNbbHyPyOEAsprq5hHkytAn4Go4pWy9bvK0285ywRJPwLByHNv6zO715eW9U3jBG
ME/9UI5tCqfB3H7AZNsUo2zYWyCM41QMRSCCOjT6g7tog430USaxL5CxZFbuiIo2TT1hCWwwurFy
ZSY/cMlp+7Dgq/vopkiQEazpiwJ2WozExbUQGkFpLwVuX39Db+zRtlS4h3T8vsTfSheWizabtXkg
XmY7zID6Igilo3ufmKOZRlb078sawL7nYuPUFNXUUWLpkuEYV7PmkL9h5vxPQhLQcur6kRqdDqqA
VDAVJvXymQEaSMUke3u4Iv7tr689Pl7Wl5tZXOkpIRMV3jiXXIzyET7ekZ89AJuzrAJVT/OYFakF
HgRdEruZyyh7UupdPwRkGeWG+iGTmNfuSQnwzqSZV4bIeu9Xxp9HShuVyY+IGRwgL6RuMU1ZNC5a
kg8uJcpkNhNiuUfAEFCqIVVtWbNoAHHcowtnWXFxMGn7i6htpzcV4cyVG2MKgWrwXygftYYzwZ0c
0Eakoy8Bsb2DuY5pTbtlfLUMYE9XrcEozDHR4B2LxnSmoXQ6MlDKO9KuDdKrj4R5bt/GlmHr+LrO
gyFnCT5hHEbwiV17wxcIGoVn3qOy+EaKtjSeFphHlXAkilUEJ4mhRaZwluHe0QF+7yIsW82vXAu9
Ta3bEn9B7xS7wzsstJDR+fFeyRntabaMA24BWkiZ/BLUJsv/xd70CVMaXI2L6Ogz7dOanCJ8Kuy5
ZfPt4f6mapQz8xE7uRHl+GPrA6U5h2TufeDbDXdsMid7/rnjp9Y3TZL4z///Qz2D95TyuxnnIexu
7x4xu+cqgPBNXE+knHSbnq5iSQaqD+SaODzbNYPYmLHkgxKyy8xgv5SssrJ1V3I7FWucdgyeO2jV
pMedVESRMighPWMtlPvYpu+9G1Pp5Ru2a8GR9mvYkrT0ZR1vZfzK1QFmbH2Jb1u/tZJGZKm4v4HD
VQ+DSFL7pSpan3t9rlXUyAsdcZek1kWVBa25c3TJb5y6eeUbbFbgt0rl2Od9U1fIgxreLsbmidKf
EUsqgCMx38UC5Is4ahnR+lO5YUQDNtFvaXXS4h0aBTLOQ7JOI7aHlQ39BkW+BAhzeTe5wq8uNq0G
SAs29rE/UM4QLosjbJ4Gz7wGW1Nt4p7acfLJieDiOypgb3oAN6WYc8eY4q2oRKF8H0cwpVQPwzQq
VEX5M88ovROaLHeHW1AMGMsDg9oZ6V6+aeKVQNujcr3rKoECiy1uYlzFFLhnq+xrFkKgfpiMiv1F
MR9FRjumh4LVL4zSKly7kwawb31Z3pFGCDvDE7GuZE20A0FelRa6UniP5/2Od1mLL0PWg2Zqj0Du
gcv9kC260NjnCZNt5WotzyKs8iXRsQbmfJ/+7eUhAXTSOjoNM/9yVAkunHUKigrWo74U72NutfEK
HztXTC/VXLFCp63Zm000ddbiS487MraSBCjL8rx7RtFfq5lNDelyD++pvGZE7ygT3cCJ5AueoEPG
gbFHQxtt9YYWGnvfP9d1t6cVyBTLCPHjRjLuR5y7t1Ty8KK44j1esiqoHGKMWLrp12ciEFyv5Tlq
CtQXil+dAu3pTh9jT5EXR+Hu2++R4DT+6MzPTORvdMUh7v4+sdwYCC5xgAvTkotalVE+LMCgJsNd
+DgjXFkHoLeBZZyrhvX6debAYF/s687gbbO6TnMoyXJ6oKjhuGb6fTKE8fZvhz8Km+tw9D4RkJTj
l5hK/C4dEsbKFbPK685x6GbNL5tr3/8tsi07yceHAeax9xFNDGW2HSCVdiISvWjqujEhx/1S+9hI
OhR8koDiJ4k9PyhE86dBeLxQGMXeFFIG5ZTJQni9Au8jlKy2oZicaj1r8s03uedJqlsQ1fLGmz9z
+LHGvm+14bGZaS6h+UKk0WmgnRWyO4SguCtb+bu4li9FC45ZFpdQVN0IYIdYezA4AFkuYVjnyXfs
6aotJVwusFoOQfG/E/bnLHBXv3eaSEuiDp0lkuP1D95NkopzB9zAm9V0lXHnxlv9GgJnWS4rbkjl
h7duTup6br4c3s6TRB+QlZ6LTXd3qhnMwilE9WLjcTBu+4NHnVMnvGWamNtu5Scxou+6Dra1ESoC
YQWlceFqSdoA8Ai/DwYAHC6KwZF6B4LB96fG9MrANMKrpS8Af7v7WbNpCsGJR56OtG57aEEQReMm
197WwuMKdQgXss+o+CKd+Pc+Az7R/+W43BHUmkz5lKd131kjvBYvC1+/M1+kk6xXpJUbazt/UcpD
HuGUmyfX3MRYjw1BuHEl8NrnqsfBA6R8F/65lKtbVOOVX7O2oO6zLSTytScmgI4hYH1NcXf2n80M
HrVHZ1pFN7hAimDsJ/NKvfdpj3G5HGe9J057p/K/t0K4QuUHdsFVu7tSZwZal5TURokApHXljQd8
lja/8kqTg4hhMf+IHMKp+RJssJzfNLiYwszwqlwTp8M88CbXFjMH+0Y50/CytX6VMTVtuUMmov8w
mSw5DJPLjmFneQAXPxoK2BilR+6SBIwwnG1AQh1IJVsTrU1fwyOI/h354J6PZBRbAkP0v0tfQtVo
l/K4VGlmty5k8ydeFjvon0/2Nfwa3idqN7RYyX9ZOMOEd9H8yO9i3ED9PHzOy24bin1911WvsOhy
Vf3RNi2iP1ZLBK2J7ZUcoEqsxV+KnSVLzS4FbqtRPwIz5Km33TWvApUylrrJNS1PO9LjM2KXlBhs
BzOCrvpbRY3pjLgFxnN77hiqfVxHO5LDTyhymIa4B3CAHTAJkSjZI8kdoR9uOn881W1hhy1M5sGf
r7ZEB5XpcCmn1mr5iK6lM5zCuS9HekClytu2vqktxBmrNtuJ5fcDhAwYObiJFHdH7g6B2rjJZWjJ
1bWpwUszm8dvUiJJ02MAAo3nT/qCoCg5VL+ctPqmmo2nioM2YsA6xHlB77vgFBlp3HMZStiAK6/+
9PtWPFfdkwaNmbUg3GCHqQGJYqj2GA0tFQcH4gg5yfVkmj7N+t4jjOJXrix0y6a7xlQof49ZQiM6
+lV+wTk6nlXWI9nhSijyzbvTRPcMlWHiyhvVr7Ag0tTP/E/Qjj4XC2rwIzXHgb9IP30QprvpNVqe
Gc3M8q6LqKBCU4TgVIUSivmZrviqHoVbL42p7PkQKUgEftleMHfR9k3sEgqjyQVXOqfueTj255aM
CHQyqf6Tycvh99eigEdhiELrGgF/x3IZs5O6k0OdgvGCxHN0Bq9osxf4xw5OjLBOd4sKAUUaox08
Wat+krm2RBfw4zTuV/ukfqC+tXB6mwlwoe21xYff7n6dNVMwKF6a3QfU5O/r3gq98c+6rVsMzMYs
M3mvLT+yOu2Ldn4E+dqiS2YCDB7I/p6iuKRywXWXZbfw8goMTiYmnWpeMB8x7DEBkmiDf3zFKp9I
GL+q/nVWQoi8eUpmF+GB/Ulx9XCljATIVtDG28myySy7xQLqWwNMDtU/oq5Xseox59hIuxWRBaD0
F3VLFUul6MF2lcXAA2qZIarCOggDoTo0PRnbFo1+b2DHnn9KVQBxPUzzzw4E7HyjXZM3djJZVWQM
BYLCwubyxsEKbkdpn5jY14WXkNP7uhVtsmH+NVjcCvaow0MEg6ckXsXWOfuhhiFi2aMLWbrIftdN
RXiI3tg4l476Aya8HmGgq82y5xgyjBbO5gONb/VzdZG08rNrZQx4F1xeA8CKBnJjVNgmFOW6VrsG
gwzrfVdBcNlKW6jwtMWy5YuOAMttdROLw3gDeiyQulTBDIMw4SJrUx0UuCtiQHvsUovvPJ27sqII
mtp+a6N0nQ+WtdCyy1NKjbJMQn5b0HWE/bngUP9XfUHL+WIWAmRDcOQq+sejC4L9vHSzkg2tQcyR
tlMT6DJvwo0UDvNjNVjZ8xGHKuYPew1t8UtQULsfkzRetxY1S34B9vR1ls48DulT2Mfklz9OXDk0
lnzX1K0moZPJJfFCUexzczxFUvFxoJO9+ObAUadfeXXzW3007zvMQ8Lc7ZmYY54IHahOK5KkjBKV
3QBX97VPat7zjbrfzsmxwlypRZT8nqzrb9/VC+d/OSM/muXL6ouYnadVVyxZYXOGQv3dqPuEioCM
A99Xwj7OX7YqmZqSIm30AXJ74KNa839uFPRte6za/4Nm+fqGVweMD2QeXcQzX3goz4jWj5g7hvNu
8cj+apOp5EKgnwshaXrGoKWToSRfHcf4e7GvKo1vEFtVuTdG81C8PP15UyZBALKNVZGthvrqY0JK
ze1bjZk6oTv2l/nWcD3F+x/Dg/H06B8GtM5n95s5ZNB/PE11yaJ50DMLKX212EviptWnBs/f10kC
wV6ZomJCW4FrlSZ9Gvbs10jQBUa2XKvIf+5+4USwGJmkQuExkC7fCVE52FAvRQ3yJx6tupc4uNse
PPG6l88xTqwlEvRMt/aL3yZmKY3sYA9+NFh7AGcjQ1WpW5iTkXJXcgn1K9KYGgZAli+/lpslhP65
BInszdzhSSxYaMXHNzpNDMVZ6VA8F4ZXYijDBOLGeBlI8RK4nDw8b0UseRMk+Y2GGQQ9eJ3oU8mA
mKOqRrn6x+guaQ4N1ogcI23zZhKWIvju0O/g4H9oiwjGuhwjB2mfbsiCBpdcGnwOp+1+Du9hYZq4
BfjAjdlOHZJJm2V0HoBoWu6AAYTdMCRknNRyqt4doJRbXZb6B8mN2U4s8Qs9wCdyqTpAHPApPAgG
7ZUheMIqiAj5Iqj+cuQ5XMAFMUOaxKWP4981M0i5W8/1c34ounXEcr83Ma6pN+iTc0+dTDbp8nmt
l639mP+jZ2JnQv6Hje/ZLE/DVfXLFHSsDpLlqvg6/8dWEzPAdoC+gJKQgoBy0nM3FO0A6GyruBBX
2IBwlRamzYgebpZYfBkna671BQhKIYCi+LUht3TMMzHuG1FEyY4PUQGsI+gDwqpm07q38Cd7ERGm
uXWcMsSv4rHdwVPt9uyxsFP+D0Inrn5urfqcSBEh7Wh1cUUUOYmuU8q9HIvIO7kSO2rgMQWxs0mC
myZEziJAPZJCBBka8S3QhoMVqx+VrWbNMyJQ7uiz/5AZQQWksSyZ4+LW4CH13t6FX8cWUR6NOjUn
jHluUWHIygjcrOJd3xzfm2CBc2EbOCZbukQUG2ft+/Ep5nxS9u7IPABzDUZbf3qwKalRX2ARSHvU
Y5E2bzuyeZpXm7IjcU8bUHPRQGdfyddz3MZXgJ7tdXHflXeScqHC/3JtHzirtBTLme4nghekALUX
jbNqlcylKxyi7psQg3UBCDq+JK0vZPzWUYhuANjfIbsMg8hgXW74B2aNiLtZmz2tuG6iTMAdPAW/
l1mpLum7RLHS3BDJoIekxPd9H73fVq/fOUHh+xoqpKVkbsvhhFqBk1KX4sGKTye3C9vv19DccjP7
HKb7bh+DNZ6uuiUygKo5WuFpkPfivVOraQMwhsiJY4T0cFINtXR1J/UrIR60MTzpDu6cGtM+Ua2s
fcIVfbBN/u6l0TUkXHngBoFZGhZQYtZF/qrEnG/MO19s8sDffsf0wtHnOuO6m4tZgIv6MxwYOPOB
udtyo5xmSGVUBFNlqwamDs9i/0f5+NWCBZqVLJeGmGRv6ou4/Ms2C8UareSOZOs5HZ3lC1W/sFcj
gV55eqNnSK+ckttvNkQbdOq+Ln9ZFAwRXAdxNNadxID+tNjFyws/8QsXPb+JxdXUX6wpi8BlTlYD
026IFp2RZHbrvBt/xQfEee5/o3q85r4XEg988D3yELjmaL89ak8wXyFTOWrCwCVDGzlEjovm5NYJ
/6LxanSR6B4j7HyQ3Z7SUHycFOQF1B7Bah5pY3n9YECkoqbBsvndUbQFYarFCXDkhpy7GSeLDo62
1xwZvQRbfrBxQKKnx/sZmj1gF9rDahf7RUbU1wQrDO1ky6j1S6FkzzxSyH+dhKmQUR4yXd18AdX4
xnzswXPDnB8dTeNxEWeFGJYin2EO5VP6SPaGfWfgacXslHH35CHPjJbOnCh+tmPojTklPq2rInQU
RT7060WEBCPNuvOx1DeDyCFBxVRG4+TLpIhOOa5nUym75V9/HGZP6q5B/KWie1nstVv7jxPp5ex1
f7jHyiJ+IxI0TdnbF3O6a7y+LWcsN2llPJinxORsfqad4wYQT/duxpcyLAmj0h/GzJJqcmrAEWpi
xoOtX8xdf3Q4wajFl4TvHFscmrK3o85U4JoPMj5vfFL/pYFRAPnzmaBFqfSyCfwFdWrzG9fO9EyS
lkzuo78yjLr0zbnTPIrv6OPS2I90BAJjPcqChsBOuwPFGiD5bqAwGXbQmVpW57prMSDeMWZRbgyq
wcHrFv9HNA381D1wL3bIK+pBDQ1rAiOzEtpmBzJdO8BTFOMEoMPAuCVVfs91pDNbWdSE+Fl/D1+8
NpGLoEIAYyUhClIEHB5i+6IfkFPxqSMHD84QqcVSV29ce6v4zAoAeB+IkB4edS4oUlnEKkQqXplu
MxuVAD4+tRnU5hYgbyVVjyP9i2sIrWLtg1n4i0IU8CEn7Kp/sxubJCQHqCxfRv0Mjo8OASOnjexO
FjdV1uPqHa1F4DOUNsKbBTuqR4URoscUxVy5I5ze/kpzPvFVyKFEE81Wezk6SJPUNKa21OaSbbVZ
+rCyGxKAYKt35PBsi9iFPxpy79vtUrYbWJT4wdGkUcRYdILUbmKybHu8uATuczK6gm2kwB7iD6ty
KoNo4zK4c/3hdNgtQVWqOxg8l/T+Kqew9dfrGZZteCya+1ypW2AXIMFd2jcSKgWZkrN34z0U9bj9
+ySD4cfIWDDdqEto7D+RQrFaHZksQDSUVKOhK7DECCGzChzlKhhTqdHLUkzWHopOVulUy+SwRtUh
e9Uo7FFyaH8oJGQaKCeIKxXc9x3YXq5nP3ArKehgzLCJhv8kB8o1/NH1w+9kyzwCRsMEW1AUiSLc
CaKQZil2vY3ztFAWNvZaxPnuTV6gJv5CJrduIk/k8ILW4jPnQWBGXnmMfGvH1lDvRZ/9v5jG3WsA
tlWPO//ctYx2ImekAdzXAgjLRwLiYvD3at3FlDauUrTTaQTWT7SP6raARwXnA5rx6j7w35xEKT7x
VoxQsUNICkA3t7iV1ltQ9ikmzie4Xqo1SQDQx7XHJ96iNRWL2t9cHPNB66+JipXPUc7cYv3GGVJo
DPxg+1rvwq3lgd9Sh1LTNCAqgZr3INjCc3RzkosBz54HsL49F1WFUHuhMVJqsZRzOvpxNNWkawNB
Ew4DA5Ifla8f8wzmi2eo+ngTPHORNz7Xu4hSbvblElCaxn4eDEhmPoClGSefsTZE6Guhyq8mKwp7
cmWlvv1YDpz2+aRapBq/m8Y2UF30luoLJrOpSkHzUv+zxYrbJzwbS2TUUOAuQxckuKeLFXB0Y8Tq
yUsbfTS/o1AVomtm+aR4R8iJy/mzfMDKTeaoAna6/KmIfEn60+GY0i5QKAXOyf0sHo1K7Y0d7vSV
PQtts9xQyaYNQyIa5u5ShvkCH2hi69GZ6/GTXad4YWvw2curnvlvT7UovLt0kS3Gt4HoxcmLFgtg
Cu2vDV8T/9Nth1HvZnudhHnYYXSnCeZo5xPcNAdcBnfAk5kgUOQNw4UxdmFlOIS9wXBTMDUarFj7
2AVHH9hWu4piK4BEpg2xNFVYyc8L+xMuAMeqyMWk+RX/Czk/zJv1bvkiLeJE4WJMlaxdCkVhHEvN
BsEaOmrs0diQ+hFijLou1Fw+17nAjbZr1GO/KU6/TMRu1GcJ3X2EKeKrTGTuxO/Y9Dy5p7w3xQO0
lp2OUSCXYPeWuRj8pNnSE/BcKIvyeO2M/JWjDmcXGltaDCVKbaIHuEB3yrpY0MVPIh7dECbbWKAL
Ev7M7TRh7jFTgEA/7ibNTHb8+kk4bxv+edflD19EQC0WaTeO4fQIRV7wDrclLqSQsjke87STpWmt
TQtzSUlSZNYYirYPjXbpO5FaCWY10aL5B7un8JDde300XVivF81cyo4tQgDIhH5tj5EEwPbCj3L4
y2ucEQgOOPoB/6GMK9XVmEhGAd3WgIACBM17gFjJvoleDR1zyW1P15Rrot5+xz/CpPUONl8pA/UZ
OjoI/A8DysjGVS/33ujqKfwGaKHRE+FKvFdpZYNqqA4ZMXrwVtJQ2F7cECRbDHtjvnLYKg5LWgB9
7h4R0yzTI08TATC1SP0TkfdyGWE/0P2JdSGbV2eblwDuNQX2p/BZCeap+r9TNXIYKkxLZFY/nAUV
itpBnLpNInU1KvSl8hBeR+SWRGkQUrN1V13QbhnypS8S8zOkbpjoifO41bdRanhCcy1Vqy+7Nc00
6jVv3oE6MDc1rzXrWiquePOXZ3RyfnfPaf1wnT3+mLO8+iwwA6CL5IokKSsaQrM82EVe6RJv+pdH
Jmc5090ZJeGRlT/SCgmxrg51beNxxR9R/8YaJNNXQ+O83dVcHujkj3MpYHz1UQpN3HMkMP/EZKi0
L+RtZpgLFgFexYPyoNk6Bm8QSDJ2dk72MeMfp6mbdh7UlZ42z40toVbjsoXNAjXDzoZtl7r3isP8
FHixhfAWNCg6wIdRmGb2O06A69rv2slzL39KNjr3eGNd1+yz6P+6fTtNnGUf9B9mHPhr01GRK4lK
QeqYe2yYVNAK9grHAwnGdrfdgBs8NotDOvkW7LVEdr1iYch2KSY+gQcEzW97waL/1+4ke+PUzL6f
s3eB0CuOOdnJhkNQBYHLagmXgWArJz91E4d0ZpCE/OY8zAoEmt5L0d44Zs8Hgv3fs1ns9LQnNN7M
80XAVUwHmkv6C2TO+bNB8RRGMzUytArUW86L075CVgSCbBNmsvsZsQMjx3tiZAvAwajRYRZ5wmUL
LkxEFuQI4AsuY/OuE1WywYDAuTME0huJjJEAL2vKr0a3iwt9q8y4N2V/WE1NLrEzl+AQMQuAsu31
zyxeaWCLWy0dhVcpcZFKi5PxciYqY3oaOneyFMHnU7JOD5lWtNacpgZGOnK4t7OWPBqO56wciLig
F1U0jsKnPwS/3uojgx6/AMa2+IESh/rLQhuznKhOnQPz6NPIR36v5dei2QBWbs2HktTMuZOlA76A
T4pWk+2zJcO64X2p6USjbYSpzGDJpXLQbwRQH3KjL2Btvi9/XBLRc5CcEL4tJb3jCsJ3RIdFRh+Q
74P5Trm1HqWiL/knIdaC/n5dDtbfYmI6PcgQ9OjOzaJddQs7BYjpig/H20wm60AzdCi1FqB+3/SZ
n5OFCTrBT3kenvOdiv9ITzNLjiVe34V1rxcgSnsuoMssoKKlOXbtJO3uUfLDwt9C8pMn7LAA5fUw
2j03m1eE6eGHT5VbfdjH96QtrmflHD94dNqzAY0Bmcuqsxv7gp7SC11gyn2B4cxjqMytLEsp9VY4
/MUiYw/Or0VRv58QWPZU9i6jceFCVitxgAiByoVQ0jqsYYs47L/0RfgtDWaj0MPyDP+7g4uezSev
sPJ83K66VqpwzMthPep2RkmCqdoLqPq+uXB+gIZnqGn+BSbFH4id+yblNyWgzj0+KyXrqRP3DLtE
Jyx6fauJHtkObMnNjuipKNPLEuypFLfM0u7/SYw6UumKvzAM40TqTt4nSyL5jryLUPtQpFmA64rz
DVUYsHojvR+9gqFv2FvwkrJ5LDBz3zd6c9ouYp6HzV2xHQbtp2q8zdHuhzFjX1UweizTxRrCMSsc
qywVAfQAEYTqs8vwP0NLDi85PX9nsmlNrEl4TJdfwlPk9aJqIkHO0MRfxpmUGMM+LUOnVoiDJg+e
EwKn6z9NqBzyb9f4buCgfloqzyVfsuX6Ff5Ncu3CUC52as/SaDrDjFBeBd2yGcrhKfbDCJyzdutL
d8VYfajuZMWzDcKpQoYotelfk5SRXu96vEqyaAno7P0vLplX5jd1AqIE0uIQ7yMnFsfjDYiutXIB
VDMwzwsGQIRXbcqIyt5conFF3WlXNHvNikU8vn0LUdqtK92kF0Aho48+F8kQhSeGfPD6XoBTH3uH
UcnCkPH7BjaylgYjjoVayv8fiDg39RlZ1k6D8gz6r5xnXS0SMo+Luo6aoo4lcpNZTS8Mg4b6TSeq
MRtyzEzY/sZq7RGl2tE3eiGwQQ6hNmSt4AdwDLMyjYJ8JsIF/S9YC0AqXcoReUP/eGpswRsI4bt3
9q41ZSIjZqq48FA6e10/Chn1R1I8LVtrqGzZeGgY+VTmZnk6miwVRR4uTg7D6UweKePmQtkcqFad
ZtZdd8WaSA8kPZIw0L3Nhri8uB7ZxZ/mszMWf7YHZnhE8q44htyffO0Mfue1f16Soq+YP9OetRDM
59pONmhK3BdV5cn3GV9ug/m72fd8CKZeFvfMtShC+8wFU+dc5CG2A7lvO2QUzyh1UqDjnt75759N
qmsztsJTnKkfxlySykCupZPOeu6SLsrgjQtxo20FFv6I+zt9IIMZ2ZG+E5to4EjbL8RAcNvlJwGp
S8yXBnqYxqLaYnjt2GqUskUogBQWGSJ0tSPMCxLaZdF7pDD+glyPKp3sxNyeVDS+/U8grziTX6Jb
mKFt9LdU34QCBeSOpjcOB/9CeMe/mP4XwT1v3RMBDmW2kLl9f+QCYWh7wrw25hJiPQnB4dU/qx7u
/pp2ioideO+f57DIBktyBSN2RdjYaPvjTuZCn/OPnFzKW0qDb59Z/kburrh/mpfjaj46/r0YI0O3
5MYGHh86FAj7hupym+dZkOs+JnT96+gWcSmWrwekdQuUz0eKj/TOOpT4R8kEDrnByWOiBkN5klaQ
JU7t2L8QIjdf3WwDOXQUOLyhEuVzsovVuwFi+8rlg4lUDzO1x64C9iYyB3wg0AR63cEYasCXLFIO
BNl4Jn8qS2Nk3bBGe7v3oafzWNxvSovxtdvxpi2ewsX/r5oEFPToyi8TOdyK1QMBuenbw0r3y4f+
cGYAPgIzS3VTk81KJGkNbse/OlgqF+OJPF4cDQCuP5EvMwp22WG7GZLpKc0N9TcCuTMXL8vNtoLY
Pzk0bXQfhBMuYJkpqDGAtMfHFZO3MQrbcjxWUINcq0aTXSyzLJJMM8kojiFccBDtQO5osD98un4p
XMUD5FFZwXkAIVjp9ol8ILb0LDacmg4zs+fXqFd/ShurQJK5ktv1eTBhYJjORb3Edti526MEJcZb
QQoQhk6rES1esAvGeGKNIbs2ZeDIGflZIxsGcLMbY+uTkKk17ZDhmwQxeWgSriWvpLNPeCUA5/m2
caE05tEAQ1p3i0A6nwJgQoBq1VKVlvfgF+AwQI0e4Yan5P+aLiXyqMVsZdKtlfX+m3S6dEkklfXC
Pbjx0u15/5ToMZl3DnUz+/vmrGEt2gsSyvbF1+wPtfmArjrbh2b/U67RYwyfbrCjDBcp9XN1FotE
IWgLOUTZ+01RQuGvtZCGcImYRsUodBq+HPN628EmoFKov0mKXfTZShTq2J6SX8x9f0YK2ZXMC1ux
HKmG7y8ucXxKdM/oT3u1yqXN2suOzQgCAJbq75riUXO6Hydfe8p0h5WZAPLOJ2FXrMJhqY6Toc2o
LgFnm/42BOQsg4dhYYEwMagw7kpEhjLP/OcsJFs6xZNnBKtCr4EDsZZjp7fB8LV2JCoeeRdRFjwD
csXC4P39noXi+rASxLHAZSx0sGmU5e41L3ATID90+7snj3yHMifwR//f8H+xieT5dm4zVXgd6Se6
JXDIcgPChMuoznNcZ7hMXGQt/7tfXU4CZUFUONMINt+oj28a77hAqhGfx9nf+zU8hLmWnh/Ywj+D
rwEk6YYsejRqqFAs3mgnHQjWqcs45jduyuTYdsohEAf2FflG8NMhSoh9YNaw7INVKHMRndUwO2Q3
duxWjlbHY3K2arWw9yneqGfw36G7CpVmOtCYm4GulmZlFkz7F17KamuHFB/yItbneFAxLx5+OG8u
qj0ikBGkavhimp7IopOjwzBTnlJMffh8xTNetitowQhps2juqSG66sZ+m2EVtTWVs9qgK1I9FNfE
5ccnzqCXfFqq3m88xQZEP0Oq8oT/aKbT9K20yl2r+rpLDH1YqjQ9qiuiD+xUimLBS1RuhGwIjC03
wDTPeoV+Px4MqMRzCHinY8mG6MZdNDOTgOlZw8CdGfH2EduGGU62TIxTx6YpN2K9UkqpAMG3sCDy
pcMw40w1+DYDwP1MJG6i/JlFmq+PbUgNPw4NWW/5KnH1sf9FnIII/686gwiSw/LShbzSXDZMXNh9
8Ipib0wgAebiAauTWpBfvl0GQkQf+DSRerdNXlsSyMN3v+7C2ZGokLXPbQbaR5mDx70hV7jLxl4I
gkH05En68xq7ZhZhQmhYgfY2a17zAijAQ3gkL+fYHdf+K00EdhBYW5iWM7BuxAnrnIkMETjIuQm/
H3hTfR9/Xojmnm+P5tuCK4UPNJLmjBiD2JmPTNuWRgXasqzwwLi8uk692IMdF/F3d51W7HG5qKo+
HiRRQMbk5YO4xFdNp5GCpmeIyjf0rEGVFO0S2NwAWI+I88ww/w5evZkpyY8MNZuNQmYVyvRqQuml
ZS62p1mdowLZHY0nHe2vYbB3778Pl4T3mplfAs75rX06fd+Z1CPhE6xPSlmtnnACWw8w2ywlnxFS
wWr5yUKStFyW6F3szlHx9EJsjWJHoAdO5Hoki5NPp4aG1vsdgcEqnUpyxgbdvNi27LpUfJIvkxCY
NQF1WtcZzFQ6Fe0/9+todKnZ/LhmuTkASL3Od7iBxaBBb8H+r+TNl0Fy4Ys96+LsAXDBwB/w98bf
Jqw/VBGhWncaPdGj9BR4MsqKt0zaX3sKdAniM7YleyV3EHz2L/sGL87ySx4YnXq3wgHnxYj8GKqL
n9cSg6KlOQmMCAvUI2IRvUow8NP8Vontznh6Rf7QrkGMytAVOuQ49vDjNtvGxza4MTY96bEuD002
mcYRjDYB1ItrApe4cEK9IYwuRcRC6UFJd52lC6kc1SIj2pj+wTERUnzdZ3Y3YRFfGb3TM2AsUGTo
t3SWRqyZVAQEbjXbHHsU8ntVWXzUoM9gg3AMaQRCbiwsWlOvjlrJ7nqhsMc9J0ddsf1DH38UOlUE
MD+2eOlwGFHDiL/tDHlCwCVB6aBW9+qYTO1vlFq1gWUahsStUxIPu0DQzmmrdHx0GXMaSQOQGRom
t72vjvxCZXSzBfD4vciyR2md+UyQ8RFy8EHd4dj55JwW1uM1pcUSSk6Qf4asyRRU2KFUWRK/hx2F
2TBC7+izVJu1cYVCUtyXMxD8to9jwPi4N9yf2rWqKHKNy1ousMNcsETRjAhBDetdsHFF8dDghd42
4sdJ0pGJKa9dGVPa8nfS+GifP1fvJOevOj3I3OW5f4Sxqm02v9w0t6Hvlf3ssId4bXDQzQUT0qnG
qP0x8F+QF7uNn4/rhUdBhndBxUWg32+DMwbv2Z/+n3tv8c5Fzka1YsuuFKUYN3CU2tsxq1TaWbCC
Cp/C5udzoqgup1eSnUV0dGjP9vTeLkwEsreGL2TfS1XhTJfJPBrLRi80RdEyOQPwMPpkPGJPX2ui
7gPemjWBF97/CEh+R6Y1AunOuaqQDsWH8HsdmMRJi5On9jjDdZMYxErohmNZqsVYmSvha44S+k0U
bpaKtvhQ8kMmBIfhLyLPjWFQTnhIVcl6HoV3JagR2Rr1bgn3/0JlssyWmI1SmABFX6uubukTtEhH
1ngWcPXFUM3QeRqOMwV/D//oHDAeKGhntYTSVZ01YkdD1ZUq/6H6ehmUCyDxJvbhj5MvRDFDP2NB
kg+bJnPW3htf72IHdMQNW0XBY1j+RiuSU4FCzXbPLwXbaNkDSjyKfI9P0TF4rClq9L8/UKKfqLNa
zikcenF/Hkkj6oJbGmxmyDUANnhV59kN1LTRcmKVcrEdxOKD95C8fpQUscJd7fTHa9DsUB7dOQG+
Dlx4yZ+bd+bb5w6NNpkZjFqgaNehAn5FZ1d3anL12R7euLnT4gFyyPsoMKe7EF/GCtYmJb6JAmzp
+ZKfey4KhvSFp6lKSPSoKC4yiHd+O+CJC4GRkFVaWB3pML1kGjhzyoWy2RMAsMNrPhDshzf5QM69
CcF1yUQuWvvdxXtzMa0ia5ucRb8axR9A//vTOpwWEXCopRtGBf4+HSn2cF4TXNgG4/CsDuvxvYig
n0h3E8EKbldJeoS5EN0Exc444uBMDioIrTEd6EIjaTIkeX21fQzCN59Jj/cOXHLz/kjK92nnW7Yj
oHMXIlK+R1Fj0omBlq65Ge95Qrsneveg82OqjEnEVe14G+aNM3z4VVF/aXLMAG3uiUObzSv+gw2n
7HXJsJHEP+RXVwe0En24gUFm+lUIynghIO1Wcsa2HbigzilBUNK9HwXhBYIUQDtS7jDAZ6xx625/
eVQB8v2ZtxQ1isjbaLgGSIBeXNFk1QFb6SUw4k199+tADaJYAJbQ82z0OFDt5lLIPfPbtiIOXASf
ypuDskbkR+wrMnjzkxDmuEVQd0gX/VAIAZdoMhEMksgCDlDqOyxk1DPeYix6Fya2UgdDAz0Y0bVO
tRPAkpoJrcdYVvD2A77cxhpBY8l2lhasv90kukX9itLxb7U1P3WDuCWuBX/utRCCZG3zRA/5J4QD
Mg2pp50S+w+bLGfgvZCcG0rjJTrNNOJ1pdpOZMyGB3bYVgh+suXkRzumFFA7NGIsagdTrnBTGYcC
Mk+ocP2tfW+fuyxb9sq9GqJ7vsjQj3CMPQ32y6xKsybdH/KuNu+zZsqONXDmMmR5QAy+3ryaqJ1e
AdyN4rExXFx/WEUd71s5oIW8MKPKjrIifLrHRhGIAH3RcbDO3gc3NWxyTtuDvpr4Umy8K/ygdd8o
mPoGUsaYfmrZlDSEfpr08Fep5NhnhTAE31DMeofUi+QqxZDIBAX1E9fLgiGaBESM8AwtpUAGLxZH
7sT4BR80+Fri+yR3Ovp/YEr5BqDnhuQP91gElucFSsucTOJVvxjAfyedQPupjWMvjJdKmJh+zTsz
+Wc5OTImEFrvT/V3cFzH2OG8hMv7WR5HXjEs7GQtjcaky1tSdfi2gCoc6VJqRhl7SYBLes+ukOE9
Al4OO9VdwzQVW6afrgOXjnC5fMCnNGl6NwrN276vWN5aLonAbjuKVmCVkNQBe1iKBOnVfHSEJR1U
//ss3gLLzjUyYAXIiQFpynivBCA+C/kbyGXOJXDgQif+l3GUzcKHKGw7WJhqwB1v340+feZZsVSY
Wjk0XVjENbTJMY1KuoOxwJr21lV72DaKdWFfNOQeqGQlrBUP/wUUc9uIp+CFuOzy2SziyHzCNI3C
H2dFQqoTMd1GAilJkTqo8mK9VAMBo2DC4w9YEdJETLF6ymwdhqBrt57e32S/bOxxWSb7ob8phOQK
s+rfSfVJ8Ki2lMPIvyuG1qfKfgNFoheootNyYgY8hybBOBOhdvAgoFp1f+0wYWg8AkfSBBiTJDJg
4KxQuxTZ6KlQgFHtb01SNSHWwCMzNnninO6zHzHaMqb5uMG1CzRdMrL5gFoVnVFE4w/PA7g5Iq83
XsFKDN/7ghjAEN+yZk/cptx2e3Qs4E1NAE1sCIrgZckuEGRXfw5JRxJSr3JfXWwUnAXUnSOFD95y
76QkhYz/jKtzwmcyN0xITvUdM8rF/r3/b5PNQb/cEhPeGBdm+DlfEJkIFUkxhPhYsmFDgGmuUVeI
uhXIqvjHB7I8QjLmbuNUX1/+RPtYuiGe0n3eBVYjeDTZ2v6L3V4B+kpEVRZ8Tr50wQPMUVSfnSGv
iOYh3JB9YrXvgqXBWY2wBkkqJsSpG3xKcwg6xKPGxYrUqnjklNH+7EJNxPG1xzPxDbJZBgSgxkXo
XWCXjl+vsFcZTL2h14O0TE1dHIHjs2PWLTvsc8gPtuhJWYNiu7AjIP1wS0x0+y9uTfDFtyULZUim
+VgMpqg5B4DjEERU5qDpu9r/wsUMidboMoZcwFdDRX2uMgmWPHlkDDGfz/llPPEpCvTO/z+8d2rE
uCld/BhoQcyf6Qu+ibBtGfhRnMW/5gBfNXS/lCgpjwd6JgRAchJFTN/YEnI4QbUOlLWvsbre6kiR
euPAjD/VK0eMjVjcFIBR1WgtMDqrNdquJNUHri8xyBoO0j7e603m0VaSC8vgthPNo/4wZGjRo1NT
T/z0ZAmFsQt1epipP//k+NDQ1Gf2nvYlw8wWzJs5O99fFHMezLsAu5pampT30dnARiqTIjRevomT
qFwS2FGbnuS9yPobIlTtPnb2J1IuxwECg97juph+FFeF5k4w1Q9N9uFxy1QeKum9fQ6jfpcLzd36
oSNe+20jKvveuFbodpwGyBY3jrCFSKreSGYTKp2jx2duTDs8B3yFjaAqojUwKsZYQi6JCJ/00IoO
Cd69Pg1AmevEA+19aIAm12+L+XM5iHj/sGT+1nZSpssUMCIZjKeHU1imj5rm5QGENcNcGj0apjqt
mfRoXAeFBKjR+utiKqTPIwWm9/4iTddKi4CeI+QoHG2UkFoF1nLopu5tWC0+0aCNtFSpIfzNp8il
Yv+ObvK55IVrrqLL4M5xKNgvSwMn42kt0tVJcHgqIIROpULoQTAuI9jkk95WvyInSK+fh+orthi5
0kdsoeTlT/cvb9FEeRK1UiQzYkTIVYQw7Ot0kVAdsqOuc5uGQqYbCy1EUxvGp0mKzYo7eKKhBNMw
9GudJ6erFKCQ5dQdWbXtauG3a2RTNO9uQkOI+lHFnKXFKMW5r1wJUVryT1vrtv1jrDAc5C6sqn3T
yWmLZl7nfsfMrf1Ck4VzWagcG9OLMKDJfz6SEiSzLDv/Lo/q1f419G3mt4v24+99id+oVPs1yN3i
MYzaoevYrvqja+9mRYfqSeY77JXcPw9x9/q12Eevh21k/vinzI6wisW56fWT1GgyGMII3tHpch4x
umoVAvUWommaGXC4bN5Bm2WprzmJ++JYsqzR1iO2KoWElCXmnP9f1Im/OoRyyMcwMvYhSMx4oWEM
dcU75aCpkuRhyX/dJkt4SEXaQmUUjhXXiJyYojDBA6Z6aoZYmzypfCwIODImafrSTbnRz67U435u
bKcRzpqYLIkGxr/MWkQeah7PJ8TF5gL7KZGew7SzFBxbZv+dCFeGYJXw6Hb+k4Y/H8TR8UxGakqf
NA9gO3wcuh/2m5s/WnNWL2ntcUuNJXKga58yoYPXxP/ARt4HrBD0nu5Ox+PjmbpbQYF8iTcqQoKm
ohTN7kgTJA16A9iFgEIvqgeOC1SJarVHoUkz14pEfgjVUIuifGYJWRoQ/+pnJPtErXda+hSslmhU
NZJJ1ENp3Q/fz3St0Smfi1b5Ys/sA7X2g3t0BNFfLPCrkITRNjx7J+NqAvFkxK/YdndFbtdZd56L
fhe20TkHk8h/k8CIBatnqsgXr2GQvxZsP616T6DVgjwx6VacIQaHUoK2nhxmskXykPbgTqmYyHul
eBx7s6jV3fHV4WQnQpO+Z4JB6WgRdGAtVMdF6sC67zfR0mcuhgzkHvDO2DUXcZVjiwwgCm5p3Kjy
g4gh/3KcOORrlkqQoyQV/Z2HNt/3nIuC4kAwI6clihD5aYYv0HBuRpkef/2keWZlK3Hw9tqXaz8V
C6HM5EeKyfn4F9cbFXbih9ei+/zVHUrkw4Div/35cCYpk8lFcU0X+7hr2NIfEBHv1lqFnWoCEq4h
n8Xt7pu6NbqkofRZWxFYaPEYw8IHPbjTT2Pjo0EfimdgMvcPzvmbKk5lJdQx3Jz/vL7+69d9ZN7+
S5iwdSwX70PfRNMrXwZsEMFtTBvZbKiATlrDTmhqDGFpqug77/4TVverwhzTbaq3Mm6J3XA4gNKb
NMQpKT4COVh9kI3kAs4uWcxlObjT6MiYqxFZSmUHxElT05VMoitf+tml2I/gA59auqaBZxx73AcM
gVeHv519e4Z+IU5g322Hlyv61+vLxJjS8Ynrr++1b3Z6ryx1K0BhD0z99wlf/2Oj4QsinBOjYGpa
/Qvh5aneQ7iKtbau5K/kFvZPFq98Y+wdq+NUoD9MPWyBbtAbAAtExE+nSK134PkqfbfI/r2Hq1vk
3EIn5CZnTqQacvX7gMcebQGXLEqPTv+1jdgfuzzaZX2Kwn1CukYEfexh9R6CmtYcDrL/9ARZRVxZ
HcXoqrl98fB/9rPglBwRZSelE899VmE9uambDq28LkFqBwJRYYU2B5B7KCds/8wRgyQCfJuxziMN
+jfyAUdHG+iJeFuzV9OySqDRS1CkciqOYEQ1In3BYCbi2NTGioyUVPHGLun+ge4qAwWgovpFeaHL
5eMt1bbbrwX0HxRbgy+4yQKRXrfcxyEzlU6TYw8/jFYMujEG3OdBB6Xaqn7LeynMoV/lc8pqYMGN
nmACF1oxETs77wICrJ0gL5kpLzVkTSRZXF3oMNDmr/Jukr/5dPMtQztXEgeHl9hVDM8p3RAjta2v
evjW8rfgcg5xGDucQad4HbtsTjpEBe0S4ll+IOtMeXozjL5TTFHBe6XZ8v7XNsS3Hbe5+3XGQCbZ
Ex/Hjvelx4bYRIDWf3x/DlhAeLKqLOA+GiZJgbbj769GQXBeDRpOhpHYcyPG+psL0fHjcRyzhIDg
wftLChV53KpkgP6d/Y8eDasTDvVcsS/WGZ7Kj9nL6fVzyaqDut66A8w3B2S5P+db+96MOLd6Z/E+
HqsKg5rpvyinpu4zxNXsQNr4Zfn1tYQeVjr0fSk5EKYYMaiKqzCiBMDMZQ7S9J22NVwWpe/JNLXX
5PzAiKTh/5X49FyMqQyQ9ynDmJmx8TxGcd7lMe5G/7Qnnf3se0IzYCLHb8WEz/dnbyoEqxNAB45d
oqfp5ZzsfhPjKjJLs4uVkxrOrhyorQ44Z3ELWOje1yW1c0/plsNIQPFGM5AyD/byNx1qcK3CEoSD
jroiWlBs1TK1zBZlHv+TMGFxOPKuQeglmtuR5vScdOuwxKR8fUpimbpjw+ZdrhzGI8MIOEwW/2uG
tnFm2ku5SA7/dAGkKKlLtJvaFtOBk40Fc27rCKhFnw7+7mQMt5nT1dG1MnSdOc3iTOrO6rqMjsYL
+kNIzCukFzj07DcrgoQk2Q9qzIpzb251chidcvDWUSc+n/S30ZN7T12yEa2qPf+wlpnsnV1GR4Tm
ymTJWOP/d2TV3VHPatVPsdubvOy898Vqe1xKBi0n+FGdycBcI9k16A0zZVrmTeJKuBFjuiy5rNd8
fRHMfGecFmgOmN4MnI/DJg6Sx+1T7mMvOoxdBUVRH4uE3c0fNQg3mPwNILUpqA51UZfE5CvPq1N4
Jo0xEpD5s0dV+heraa7jV5tRzVrudgcVpUl+yMVTD2NDdzJ0EdTzm6MJ/DvvKIzQx/fGdojuP9RO
Vdhqy8FYWhjf35KiUNtGhItl3dmSGtPi5Z7ivCsbk68OHfsNiPIV7KUmYRYAPG+TtHdBsGL/Mgp9
rEDvFu4Ybu32BxsUTaQ5ocSTOmD6Ls3lZZrU181G+dGOZTIYN82ULaKIhIAktQFeE+1Yb+5J9IdR
KhoJVuTcSQY2jUewN5sBvqfeKD7DegxHz0WFeRV7lPg667+vprNbha67qGKfDwIS3SAwKFHNhOVg
8wTpk8tQKuFkUZ7rRcCNwKYr+oGSoDJjWpJzHshmSaXEFbxYQjXKzu+lYyBddlO9ZFuCndHU8zFr
F6U0PAgi3XpPi/brwZY88ucDaxG0JOHowUVjpqRFh56ygPfvYnoIVZeyOKFc2YLRGok1j0Pm7nLa
IjPTW4l5pSkmopIB1t6IPpyyB2r6OOCJcGo8y9qBvQtkgDeqA4bNDUxsV0zmZqyqbZTkCpz5fiBj
I7p3R/nMA52zAVJHyA7UKYDqluh//BhOdV5aa2TJX5ks8xrbWVAzxABVo5Hdpo1gtAuq+6ObWvIU
gC6PeFZbbfWUG1EMUcyT0so9g7fZss22bKiBYNXgBSgZ+PWS/83JWiUxVSbZbqq63E4nscPyniHM
EI6N8KHX1cJESDg4gPba78HmavPPqVye7XYBCB3Oz/vf8jcgypXy8umf45DMi4aI4BmVQwRhxTM1
Y+7KJCBl053vqM6VOPQ/EWsKKTV7ERYSIF5sPKxyUR1Y0ypNC+GoK9Dl/0IZ2glJ3Ejf6CKhsWeU
SKFFWKhHyiYtAgTQNNJKm10qtV8Zkv165DKtbzMg/7wcUP4oiCywK00EsK6dC7Lq+OF+vg6ASY2Y
5SyVOKR/C/tT/Ra6VGLBW+PCMWZIb9ag2CKhTWuJHHE4Q3BBdxudaDZIbfKzB8hbQXcT7se9KnKp
mTUxce6zfp2dV1TnZoyaY8mzIyOqqhqYpdPMrqCNBj95uoBuVzgiNKIct4x78AaXr8ngSqbRjswm
vHK1RlgYuuRulLEBbZsufinQAj7aUy8HUeZIsOVc8q+ZjgL2sxvuJxnMQbThMI2+1NrMwDImIDVw
Gh8nj8/WvagCD8+eAGwjht8Bu7UMay5Ay1rl59rI+p8gYh0TeKb0LybTXWMAhz5fY7BmT/ysyI0m
s037Pu22OrodCSiNTe/6saqxERi0GpgF0IAO/02JuL6Knw1hMWidq5hGFvaTBG5VkaOL9bywlIPx
kQy0imK63K2cRwM7Hkf6TyLgLuXgtb0EAkwbN/pHSbYbuSH8ER+aGMDHsPqrwZGIg5fU2q7o8IDb
2MfW6GZ5/sLR2osQ/N1Ap8pTLKWCOhivY8R0QP36VTcQsRTavU5O7H70oy6CK9zanxlTn3we40I1
ZTjfINYl62wQWniTW/DVOLVL0I+l7poAUktYiriNj1ly4fXfxLhr7xKHRJv1zcJ6qV3sbc9BUqHg
tMlnBqt1eRh4ImuLP33/kzHOl8W4rZG6J/tELCF071134ftgFCn08VmhaglEuPRjiN9U0T4pDQsB
FwC6jB7O2z6o2pt4qzPoshuhNtTxPH/ms3Pt9KqlcBhb7BBzNxOHxJQpChRSTZ3d48rK7e5qoln/
mOV2rqTOTzDNYftmKY/lt9BmN3pZ3ybfK8HQ68qfZS7eZTXOrQ6XZWRUaaSHJSdgJ5kewgv+H4iA
uoEE6s9ddI4R8ruZ0JimoBumxlEJ+L40cwQYamxcnRY5y3kBRystLQAhrFVxCpORxtFeCE2naSGB
8Rte1YFSTQ7aBl5I6dKtx8WOVYFE8hju1wWlIVvf8XI4l8wmuoUz6fiCBgxZyshzXMDXoaJ1r+Bo
y2mQCYA1Qi3SFYseDQ1XYxmFag9GMUWuYI4knwabSBLxoxEzmaIESGoPD6zeGdQjn1QDSXGZ1LmC
FZ85QOUh3FiviVmpgHjwm9m3hd9aUaGYAtkNyFXZiq3Kr3qzVjllCdXcm0midVFyQBJZcYipTqFY
sNyhbl3QEdeyA3zan1FBKtX6sSpv0djotzY1SwYjJI1I93KgD3LA67KvTeSGGYept1EhaL4lkOF1
7sHufT+nDIH7qRtoB6BNaO+F6NjLda9xsQx4ecSynJrMsy2eqxj1zM+JDIY6q5PoEheNahuC2Wqb
DQrrJ4Z/J4lmwBDqH5DMaXvce0POg1/9vapg+OcGHnYj75slMdo0TIKDT+wzUVBWt/V0i0hTbFVQ
GyULV80RFQ2/4sZ4vuhvB7yXwguE8xqABtpfMkgfYKs9UnIXdC0FndZqvvXL0BNLKgxsHePjglZl
rQAEQQRfrsG+8QtNHb/kcedrhkjmzWyIn0sEpy0598N4lfQWK36eprrseeJBM0R04qpz5Yn6O/Pz
ipHLD42CuQPsXCyP4ULkGlESEPdjQ5zdXxBBbwdEv/GW4jPOb2y5ogkKcOBGekPpCcdEJTNCzt7P
RRmvMTO8gbAYwSkES+E5kLxT8JJzgaVyQLAZEteIr97+ATvKHU73/sr2G/CbG22R7ic184HspMdu
yutNrEDOR+zvdIygfXOVXLVHKyrJton/nadNwnLTCq/SskV22NuaZeDtFhofAwrk3Xhrw3GhvWwl
tjPRwdfpFxitkbNnu5MY8rhXmUw041rUmbdhbJZzBwkkyZHRtOVhHLK1X9rYdBPjSvUMGQYkei5v
ZJsqF5SlthQ/Kr1k+D74I4Be20sUXFnolYpblPOAFQPKN2cvWW7n5O/Jtn1FiRJTQeicDX8joWx6
YLXkJ3At/btx9MNO+cRmk6Xq7XkxaKJpRbw96CfiNd0qjn4nfdp1Ue7R/n8FD/DC9HwVHPABoDTY
Xfr72GVQyfxcyGjIPw6fi7PYJMwUVk1PhwFnVUxN5PJdtG+thmQqxAqNFqp1Nkb+h17cY1h2QsEg
Tjos9fwelLTG0CH8AFflwJB1AzZgF8neAh+26/jojS/4Xs3ir86ZOMqdIO2Qhk9xYNwuWskm18Ht
NG5fLD5lOg4I4XC0WmrpZ9W8UvYqv8NY74Up33Uinpug8FYcOlDQyeeFs7GfKj3d58Xt9ivkAgXx
c8YR76hooycIG2lMdZcnC/NXfhxBKlVKZYNkkCq+t2YT9Go7MWz82atY1NzgcmhgjdOcFx9+mWZv
cIaViSgFM+WB9OJQc5wc0CSpubETcBq+MlA7XhbHAe6WsYMbvVHkjHHa5/SopTqeJfHxCK1XWqrD
J3acmTCAqziqW7fYx75yKVUQ8Dj/H6oWQZ0kS8KRGJJJgWWQlft67PnSb4w53ohUT8nr8AlTQhEx
TXSkfUIvAska/2kNWdLKsV0h9j26MyT1qXCm6ymEu6SvWQVC1+WlqcEVtoIZwWh68stBbvhWdmat
ibO8WoqiAWdQRqH+c4DnmcEpoEJBgLOktAbKpc/ujh/AR11Q4XEVlSLa1JrL+VbKUSvgv/oQhWnV
IAoXyuDOWNPpLpJ35PW9tmUx5lxngCDnObbXw2WfzLKEJRCxZPfOluQYicSZ0E3UxW5Z/XYhAMxF
oLvOLIyJBiMxVJ89RgEkqxNQWyfu659P76qAjnHfhdiJtLC7CnPHe8yL5OTJtnFlZ4BcuEU3Caqo
hrJWPja6WG36lIbaFPN8jpg3x0eHBa78W7P2K/QGOAIph6A9stCRDjCKw/TWq6+zrNbjMCFQ6AYD
SIUJlrF40zfDN8ImI3sqYJsVUcE5w+cAeJnwpFBPs2MdVCxK9hILOM1c1Nb8Ue8Ws9AcwDKgodmz
HW3QmPnyVIi82dxD8B0lD3r5RuPrCD8YHyGTzjl/VnGjHvx4mJ50RKhMnsWzwz7hOHk2FjFDYLsp
K+IMPye50hHsAfKzYFHigtqmIO7uLJ6wouBLMOSX9UERcTBMwUxzyDNSFX70ttDR1hntah/X2FJv
GTbvhhA/2JnE27LzVttIQm4KhYM3ThdsW0gZkJbpLtce3ZXrDScmCoWCuT3OZfd5qeMRzLIGWRpb
WlV7JcfGrJWiPv9qcPuI7GbtD4zy20zPiqlp8WgabzR+CkSIwStRwJfS5gV+RltgtMWbPU0CjAoN
FylHmB0A/0zTenqdb33OKP2Dls/GSlwLsXRxSvBTGQtomKp4iQXdHD9bTxZMmaXSUoNkJPgDiYx+
cok+RTgBEmFXTDFGyk/a3PBUEbscQQKUb97AppIp8DP1MngPTh6CAT1H6cZcF7D2sVoSddD3gBus
5a8b3Cdx9QjT8k4YuwL397f0+aYAASM8cJmniZ9df/V9LkKM4MySll2teZYvQMm2R4Q33qB1VVYm
zq2gcLL+zcxfLl65bahqg8p5iED1nNddrdP4H5XGTR3WgApDXaYS24qy5p01uuKy+BMKB/I6Aa3K
GbLLaLiSc+Dk6zxh3WpEZ4SIlRvIGJLMPE9rZoLPrVoVWpoy/SxAEEM+r5TNFr0ViSGmYls33bRS
w9Zeglz1KrMF3PC+H06Pm2S9sPoyXhRUCLIGdGaD4BMP8utr3zJFQVuKAGbl2E7CJxNp53D8m6PT
ZhEjxAS9sd0iElMFFqHfB5z3r25uXmKItVjeZYO1FD5HlV5YdYGuhh5jwx6ta0yloiesRxQcPqsH
k5CDVGcek3+s6POAEYmDXZi/mMjgLpcoPUzmr6sViZDhIo07LaRhvAv218610s0W6029rrJAa65/
wMAIPcmU2ErSdy3Swbv+DXOHvYouThBtiaCnQ3O6qRSsSKODR6EsoOf4K1LtoloQhvuSJU9rAu1o
udj8PJ78y6dOyQ944mJC7TXiZnY6+K618dBv87boD0dTv3UcVMuEUl8ZyiQxBtG00mpqvO4V9AvO
rOTltAvzQSwmP/wBhHBHf0nai+X2auAw51W7CKvTAlMORZ17itTJmlLJT/VcnjUIHTF77MyhFil2
hJHYWV3/wG5tcGra85vQ4OuFtkHql0NuvEZq49dHrkeXzJbw8KKzYQSVyooZdh+UIWDk6WMtnd9e
gnCVCzFo+wPpiqV2EW2Rfss9LTCSNwrRFPjAqwxK4swaNJBVeVtXcnkrnMoBpga9XAP6FApq4iA7
X54hw0QHHUyZJxKTFci5eFL5qBw52IP8U8M2jXYB2mk20sY3Jd/B/RXt9PjyDZ68N6n6G95bZA0h
E3J1ARB2IaK4Ik/S8IVQPC9xlWrTFBW+l6DgzVKN6AmdUPQqDIIiqG0Gv/lrxeIKGu/TuoXut17m
lKqV12uABo4T0q9xqK2YiYhD/Jspqh7ZtCU7wJA4fzw6g9eW2nqrA+rNebkywvSgc+O6ikjC4u0L
WRjIBJjHjweR7EfbqzugZpRtVvfFYbMsLo1ORj4n0A70db3FZwywM+21dROL0PzVcALC9RW86D14
r90zNp+9eaGVwyIIwk/AxL8VUBSW5U6Lb/zLq/6Km/1+ZE2nCtp6QXS7WaDJ4/kERJocMk4gtM51
W+Kb3TYYNKsUZx8SqbmxXyIEd1pjLToIIBjLqwtk7M1hYosVdWvgtr2KYyX4nKWUQgv4iKdV4fz3
NX/O+IqmwkpQbAPSjH/Pm03xtZ+F0LnVHQN1W7t5WzdT/gNo8PmMaPb2cFCoSoo3JGlObBXOFx/1
04UAuFb8hdaKgeu5i79nhu6qkZwHqTF/BncoeF604Ybwp/bYFwad35+kVGnnOH3SKhSQAyA70bDl
tSTpmen5K4IAOGKrHRSeBgd8btRT5/bL/kdcJ3HgQ29PUQPa4Spmc0361Wz4niz+UBprZh7sHXXQ
2DJxqBkmIht6ZMBGYqW8IHtWX/WDI/GsWHn4clPO9TOuoDP2zT/6/DLnjXRa7Hh7N2s9HMEGMPs8
hH9TbyokDhZX4LcfXpNIcUoigMByq0cJHHXtUhWbB/ta6lkCysWzBDsinzqB7aGPUYYERkAbp7/8
GeEtGt4DwZRqU451756HyQSgECnDEifs4Xz2vFRIxg42fTOAvBbfeSS8gtTXo1qw2L3LzokuWAKG
aenGegCT63ZFoSj9wioZ27mzMboRAUCI696cMLHZwAV2fQeoF5rDmwOhYGqnFuHxvbKYFmbbY+1F
1TTffCK46LirGGpDkxtvYqQ7SacPl9aro+zl47pypVerrjm+2XT/HFQA/4sFadMlEpHXGQqhBKzl
EFMHnvosLJSDR7VuAxpY3d00FDOwhVar7hOBf3d48SDV/Sqp9WF2vPYLd2QSnouqxR9WZZH9IogG
vTqi2tJz3dkgD5IH3LeCOf7q4/CgppPDqV+i0yUumY9ZN5+9GUXSiDJomb/xf9M3lHzpXztR775d
LZOrspxp7nhmjeK6SVaqONlNNFinZoaazT8cp6YuWq+sDXQtJMz3eqoNk0BcXfKc4sR7gAn5QWNC
IOg13rUWKqLqkNoC49DFun5zzT+jdYINOO1xkylAF7VKkexdbjNxrf2GaQU7QBoaYzkrUKnYXrxo
lweveUU/vPStWMaJ2oAlXXhTFSfPiKXCmc7/l6DX8TclbsJ+oWbEqMYLuWLTGccvw5Qwv8QYJslo
UVya+VbMl6X+86N4YGDR8RWKZQeoGhBXwEyer9osjo8aO5W5MUCtAInyIcqTnpnLI4ZcOnNb4uDG
32zeh1Fyas8kp/s0rVkB/H8LlxG3N/H7DdPr8Q9Qpl3p6FG3MdEVzVby0qRs9v237LOgXkulFQCE
OtoTmGIL7O7MFUflKp4FqUS0EnWyrrQql1yhavE9zZ36BMmjVqUfy/MqJnRnnMJJjnD6QljIencx
7avtfzQ+HVUMN6MQk6xM9+Jg430WGfHEWpaYroSjnwyKJLLl9m41dyhsLhXudR+ets8CLqLaNa+3
Mkks5Wd2Q4MRtCf09wg9wnEnrXgy/9w4wXRWv+S1wcwEOtrVada7+s6dJToj3gVsjPRM7t+gXsVV
J1F41pEgvsVKoREwudptxFr9flh9myg05tX/9xM7UpfpNEoDZSSUPULPXpDJakosnJLaK3T0NefL
FmNZtXRv+86ASgdJnSNxxFZT4rHM8n5SvhfcOFCGlvP/dya23X87YabbED+uZsYqVmKXwixKS5Jm
m8rDpkQF458ESXf/1vjQLbPBpXh3ruKbFmSoms0LwqaDS45ea0OogtJqokHM7iaE9BdyAZd42Ba7
N5aaeizWhAKcSkCi/7KnsW/W9w58un3OIejKtCLjQSKjUOQ+meWO9Mt7SiocX+/7MzTkglxejdeS
e1aQNEMz/+mByrdEowY9bzWMhl9P1TF4tVlaEYFiCCZcAako2U8UlKRTQcfW+8wDplGTmsPCOUrc
1HmYqhTX6CW5k4bdwA4pitEY3ueLQf7UC3AyfJQcFBUUfcvFmuescUuwVVeyl+PR2irixxiqxxT7
5ruJYSlWRYIS7p4HstTvgzacyseCfdcZxQb3LE8MJDwmRpJsJE9+LLcxpaFyGOVX17YhRr6qAlcK
ZccALcVTfepVrnzU58osx6JRDzZNjKFKaWHJTtp0j/U60bVlmMY5mS6olFpyaL2s8XzmstxUi4ir
E+56QpDshowSvYq2MLpxlLLbHhsQt8wk5ABc95w9efcFVktH2q/dlR1qUKGBCtr4f7ZJIs8bmxUK
FKaVoftvwVE3B8kwa+qwNTkgRuS0K19VKZxSsztrBAk/5gS9yn8YYc5Bq/hXJa3gqRPO3hbuTY7F
/D4gXn57AQcT043HaFDju1e1p8ioI0XdXTk80H6CQ9IM/2de+dKOPPEVBzJDURkRf/q7QXQVNdVm
K5tCiUuURWs+UUnEpuUb6Xo10kmse2zNjvi8oUDJb9SzFaBBqXLnC1PGDOSeCkZ93+Pab74omFAJ
02JevPxu/C99UuS5kkq7mx8ZPsDUhcCHyrBlGTYUYOri1rLJWKWJe+gnoIJbn63HRQNrAuaSq8LW
K58wWjJDDpvEzighk5GkOIMMskxzDxjDVcJ67juD++sTnzFiU8Z8+yREXffcIXjsCiaDclCUnVVA
y+r2/u4SLLyrmIHJx8L7uG0mNUmfQzhCectmZrY2DWLXW7AbvSKx2kB24yozmdjzbX19ACSPYgDY
y4is7WQdyi2bPS/UKHUFLDmSpb6MHIcFGSPiEZS6hDV2cV7dOE7Z/Dg9xvTQsfXStBGlzGXodX0H
1hzLfcfWSzBU3X2epwfELfpYlHXC39imYiskDL7THxBcaVbF/WXjHEgWpdDbxDxRvH3MsliszMU6
bSdWNXpjtSbWUWHm/sTbwdQwZF/+Zx07qDoRsW2wJkJwKL0FV8padVnjuRJQMPVI80m4r4noxxPn
mf/8My9O4rjkPSmov828roWlEsSxOHR3XMANFcM6IlowF0Xq8vPyD3gF7rTyH1GV0vVqPHOF3qCO
DvHOF7LzCe/P+X/bhsnw3aUgYya6h8H8pCrCRSFNC5KXXnmViRk36Xs2bArkg+PnjV18Tn3dhLm7
xUAxfzg25mkgg15AXSdQL4j9w9jzynvUQj1+8/HTN2Ft8MkPjv7M/YSlVqTa6FxuuFGEK42LCpV3
P2v5pz6XKA9mKUrc23iM4K7tAn5L7Pfqr2tNkTMB9X1nWUC/SczREqAIjKwuX+HelxRHycQj3RTb
2Z8RqMdiRu6mesHa671PCipIFZgMoGUtwMp2tdcFUf+1PllDdWHHNW0Q5wLGhVPpXtRg+JqNQfhR
tvPL4z4H+plzgPzPptYxIP3BsMHbirZDzVfrC/kZhXdkCik5GbR4moTpRzvlujHsshgxbwvZfJCa
rN3i1FudadCZZkHDOSGo7hMcoXj8wrKLOgLeRmBNmFlCYZJda50m4Y8jk5HlfyPonxBG0oilY/kF
jn5GuBq5EIAEavEC359zANDOdN+bQJebgORguNmMlrB4C3oB94RGfw20FF3X1qUy/eZCM3faiPrp
oyRaW6NwlxOJmIQNwjue7RVyN4a1G7Hfxx5Hy8nX5nZ7qV+zHuBZQZVV4SP6rRsJkl/tF6GqBVpD
53nZlCfqeeZwa9EXu1I4am0rGVHSbNyczcr100bASfC7fw4ETKP0JRziErNFKcsGEuoZlZv92fbl
Gc9IJsp2Dz0JUSQwlQCxwdQYFUVzqd2Hs3BSfjHGgLmwm6qc7y11jflZCgCIujZYmCwk1gFSBCsY
gwS51kFzxQ1b4fmzfRRRKTSmjoB/7xkKG1Sfq5dMTwDt37o9TBh+IweGfQ/nO0wjMDdiaoLNv00f
SYQ9CooamP8CHN6R0KwmG2X82trYuVqH6AjSUjD+6djDAPSv84uUzdIPUkDkbR4y2O/CU6UAutyM
iyg9Y60cx+E68vWOOfFSDPTKgQ7GmdMUITHteTaVBo+g5SLn58+i327J6QBRz4p6qJ32W4nf2Ko6
kJNHSXCgtj6BfCxnTSf38uMqNj0BUHfIRuW3+Kh2Fr2NOZD1eX6vR/UBrC0sSYthJy9BV5Tg5PlM
8E1E3a0BGXSy0i3x9dMyMg/s9V9G4cL3Cl8+BMr2DsOgKBv+pFfC/FGKVTpnEyebNmyt1heouNcF
JeEaH34YzxPwbcMWbWqk0lt5ZuIXAn3YqR4J4Oyd2m5Untq1n3/t+089z7EdfOBkXKzH3zArIy5G
Jtl2NxcpfUlUFPY6Eb1CcXLJHNhBfdeAxfUQIzGRNa60gzWxWD/koUSVX5rQPyMtJ7E0dC3f7mda
B9qpcEeTuInblS4p90xv6DX15m/nR/CyKXTVtFCr4v2VemapsFxS3BZg8foB7OkAxZyregedZBXm
FlCmCUKkH5uxWJSglUnLs6MYhPOruruAxxrTYocmlYzG0ayX8s4sxmVYY9pC5082Iow7ulxsdVmE
N+nINv0SWt0m0TWIcJOb5FXmT/Dp7N+WD4ISZXWrp53DLeJ5zgrKDm1ofYUltUDWyL3NMvhSVZSX
1MtxV9514+sDo7BfIv3meKVyB0+05NDjiRsLpAncBqB5CklF/uRnyxNVE5r1mlKuS9JPCoftEkJi
5hGSQjDuzJfYWoXgvydrEH5qJV7mxxDmIUMPrMSmtfNU1bS5AB+/0u1Q2EK6OOBFgTV43nomVzKd
oHAUZAn8qJ3sNUKjlzeAQDwHNFE8e7rf+TfOFY/WkOTJBFqeNgWLzhYZ9exvpi/IAXKR1XBosvOy
VERTORsA5NxU3VaagQN9n4XuRAYvwQt69Bkyw7HyLyudMqDIjbB8ug/l4cUmaHA7a4F0PDLJSK/c
JQtG2Qs3E8+sj2Lnrkw3iUwuw5pMJOVYvldA+Co8er8LReNhOGR8xuOPOILpV4zVGSwPmEsFXTZ5
yUppym3sXKd7pgqDAeXkZpnai9uTUsfK0Fpo/dJswbXwXqVmr5Pmua7aihnLRRNagc8bX+lavSky
FfN/WLosYS/BlSdsNu1rannITBbsiiE7X12k9WCRg9xmmgVirlfcDv9CduJZmDKyoa039JaLTmBH
Fup+bx1CKQm6Jk45f/PYQDgYQxwg0wvFzvVnqNeAUtKQAP28nre4JjnKfRUlWIVKHscyqpE3KaE4
f/jdodA3IkNN8oyRhGXFgIAiVEzf3pocVxlxQ4ZWD6QjyLdh5+dJRvVHvZLuFLqolAsD5jqyd+kC
TnD8UWNIpppFz2Im6NyMauTIjjFhsdxj/oy1dwfh2Ud/LcW6iKUJR/GhvFNdFn+SqthsFXxsTS4s
6lYfmLtk7vdJ7rtRN+pfJN8TFSSBHYxO6prBY0UCOqzIUz49Y+owqfS2bpkXGwy6wnb2cOD3MOsi
5r5qTB9mtHANiVbbDvqzBuhOl5Fd4RGIAJ9oBUBxAQLzh4ZacbSbLOmzhsR3MjUXG5kE+06i2N95
IWtJUtsY0v1J9Uwxrf1PV1sb2I493RODT8wpJaFjQZeC17r2TSZqZIhwcppCILvO3r+4Xar/IZvE
niq0jAtMJ4FeH9jOLz7sNF2jEZ+/hvyP2ldpRt+54uNtBMY43+AlwDJ0tLS0xJg6seVivuWMjHlI
x7J2r/ZIAV5l+DxMhGCUVljKVH4eFrBndGxXNSJgLkfQiXou2I8LRCZqF8RfyeettC5lgKF5nOd3
edZfPo4C48M8RxmCaWxwteqQ4hEGAL+m2KynMrWimZz39wgpGerrp498Ys+w5KpXRJa1o9ADmJJ1
lp+Hs/j7qyZ2W5Mc+JP5fXNXhkzzVRiPhMx3NQiBNSgqk/3AcBWuSOFzxo5KRz3LAgpR4B6HZNx/
1uZhngYUqIRwcwFn8ti/IanMPwu/EdoXJKL9vF3WZjREwzHgxXqxrUluZG3su1GaGuLRy0H9mmeJ
/Vns8uPSsaeP/0LFrTbQu8wJalEE1+d7Oy9RTHk/kSjxRaOoEsXszb5RBQYw5T+pQd58lF4ATBGU
/y79igJmFpN44f4Q7H4R9GyI1ebh3rH8FOvJGS+rcv2HLmLn038RgWcyxxwXp3DKlQI1EA7hfvXl
px1+wtt4I37UUT7WAVMu7uV9jtboYiW7HVLP/iD2YdwXXm8PYvBoHSYLWLejVUvOxMZyHid3Wk2U
jnFCa/7wLVQALfTP0CEh3qg4ntwY8m2HzyBbGILrS6+bSJuFvPe6Soyb7OkQjytS1rOTXYAZ+Dd9
2tRrRMnZhVrfrA53rG8/k/9LYBUR4IUhXbd+bHLwBXrTUChbDzxYlgUofgBqS6Wd0jI/41bimAD2
xnnqIhtBvbsypYNAoGWsdy2uGW/7ZFT9EniUcRB7j5Kz8G8MXrdLRI1hw7lza5ONB1BMaU8IvgrA
9UY4lU6rEg7StlTLZe3d0//KfXw8GMXjBwy2Bs7WLwPtRKQqKfeCCkmmUHxygOQGfP8R09WlbbRj
znIEfDDF8x7O+oaUTTAijm3tX2xXU1VaiqE/wYWNrXPWJyew35/MwqV9DK4chq5SaY7PAk/JYgqp
K9ilncbbZ68upz3aDBKymetOaOGVjJ5sIoyVPc+Y2CBMD4udzhQFSaDbBKEHbq0MAe5ErnKsfYN4
fjZxGOb68I2jW3oMx9XCOJs8a+YOKXK+QLHS/PdUWVRLr/JrHPqft8a9wh4SQmozx6JHZexfNPPl
EQqhaDglpa0v8a598ZLhV/Me7uyXaf9GvtIid/Ttdf2zFi0hNqWMpPIrXg9cBMB28IDmGETubOhe
pp1ctckHM8i4/mRGODj/IPQvw34hvsL0PN2vZ9D0jMRFSNY92DMW+NTbRKQ09LAk/tsVAFS5MUpJ
wf8ZaWfxi8ZBf7ytbQx74XC3JJaj0DwLKvH4Bb1KBrVZa4MtKm96wXNqz3i5Txw5vhtG07NWvR3E
tjE3qDO7xNKZ9+SVIwAz1sdJVg/KDmcnmSuM9nATsnMLivuAyHMjvMyOFfx8LEsfgEVuc+tlQrSZ
UxdMOoB6uEwJ5pdSqyuPrdmNAFZidI55B9x/4Xp7aZo/m6WNFa9NpVQOv0033pWLm/ImFGQR51/H
wlGvfUZDSavGPaLKer7c8E06ibSxAjZaJ9LrMI60mS1EooS8rP5VpE0pDQ9DkN42KXzcUv3YVJ9E
zFV7fsS0eI0bhS0czIuj1rEHdwiqIuyxdnaZKiVk8PhJw2E/3llx5WgAfJiOioZLEwn0lh/m7Xlk
3IPgb7Na+q/HpxHrbEoF371D6u7CgBE8aXYYjtpLCgZKtftHymtepIeqINKZPFjtlofcbK+SH6Da
jPgQe9e3wWmPLsQOQGIXC3hfIHqY0z13RN9KQYQqWjU4fTC3oMUty+imyXwYrn27sPsvsrSk7qMw
N0ahUGZavivZXOHaXRzlRlOdjUKBRVwHd6VjEUR4G6fojsetUic4d1mpF4IIwc7XaqC7RjGIlStZ
O9FsjkQkk0BHCitrt3uyyG3bUGDqldH01FoOW1cID5RpBgV6O+tGrrheWW6kDNWhdsKntZgLjaTF
1imyTyDiVHopRBnSpEgnAxVSAF3Yr+knFKTrVD0V6P0S0YwuZE4H42+yZBg3STrzwf/yywGALkx+
KMOvF0GLre9adextFHa/peqQJQIU3JMf8ny5ejsxe6BPpr3E9YToUHG7h64CtKGw6YiPCxOjwRxm
fZB4qIAscDdFfTo0FXlzUfS2/Zi9WlhGYL4FApNJEYPwDXq3KJFmheIFpzEcGNQmYBMW4ccsagxN
HcpBykbB7IGxXNzoLMfeAUkogoUL9U+Riomgem8i+YFajIGgMZH0huONsns4JKSzXMfga4OssC9a
o61dUYnnmHOI9R04oU9yvSboXAo8EpWnQkK/H1hbCWphlvBa5d+GJm1wak42zP3a5nYC8hsRHTUK
V9ksQO4G79jI3ZQxU0A9FOR833+M4jkRqTtSNDu1rD4rGrGkJEbpu3KCZmOBhll8tL2GFJ7cUe0t
67QStNNaZPQ29rq0/bO6rfy2TP5KWK9adjctEUiadEDAsmNyp8ULHoDRAh33lBOxa0JDYQAKjGCn
Vffbl7WPsvfpnr7FaL/9PEy+1p0U0e1ASnfBF2JCLOS9pUW8v0qa3a4rvH4i17809ukuy4Wn0Tih
1Dfs2GSAV3RsI3cOyEMmDqaVIX+fGQxm3wU+674zBbaIIKVFGfZSbZm7shcbUEIpMnVliblCzmNX
nZ3Agmk/AI0rX+wK+a8CVbLi2N9Eb3fmNHDMeWC+ZnA7q4F0tHmHYMhLp7ghcK1pyv4w0yZ6reMi
45ifqbwBx0whErrzgn5jMvJ8kIFcih2F6Z4AnwmtOJB8tm5cxjuXRrWSMwvo1xIu02LyUnHE0Hs+
T8qSenSaA2OVdrCHK4RpqMckxBxrsuAksk6oKpO+7ojY7H/G8vZlxXG+1Vp8VVJblA1RscoXr12K
DSVX6RrmBN28+0C9Vlt8G8p8CXGCcCD8cMCmsvV7b2gbdBr9mVLpzxPxQFNeevKE8V4gPG+yrfPi
4A8MZA3eQcjk1ruMK+vI80bXjfMgME42fI/2kRoJsbijymV4+TjdZfvR13RfWnpyZZkyD2zgByqw
WpVucxfWT0RpVKD99umq9acb747P6YrKvUHpUfySxawSG9bJ3MnNj1ZkN+enGYERWNpg2eHAkP5q
L/dhgv1BydrarABWqKcqJs8VCOndjjnnhrLZyQUBxa1vyMR6+fPAzaVCqYixO9l/3T64ixEqFGda
zGBOdzJNGcoxEzM6bGgDVL+7ghFoyGw6VCfJFuOsyNEEDzeTZPcqtGgRKPQSviITrCp++CAnZL9L
ET3LLb4Od2Wji3jCcmAY24sEx9kqIVCCHztAWoC/TZKjR3geoHv7F+orIegTnRAbRixmnvDGU3X5
uXj6t5AoDvf2FM98rshlxBo3I0Woe2PISatCR4/3isvVWPoal2zaaoA3nJ+LSM2EQ1GqfqQtr94f
/BJ5oaeF43qNctaxfSzDkki1BwEDFKopV7OnMQy0tw3eTjUOSwCDtQ1p2iKYPikQDdBqCJhFsXBU
UENl49QKU06Rd09IBdgVpUOxqlqrIImj3AvrnnfO0n1nlKmdckuy6nMzHGUbZUP67qvVgvnPXk4+
Pljn+qez53jVajH/3tNp1gyhEjMnng3rhdgZSpxf/Xiv7I9Fb2PyxLENTxY2Oa9mXEt3gevuS0t8
yNIsBKw+73Etm9BAwq33fbG/vz9eGH1Ri7tCkIJUt2f2ZFCE+g7I2pn3mcWm2ECI54XY+5NXXW2K
NgwiZD3EuVHfEUo4jC8T6UPswMBMlxOQ6WcGIoW5BJc/z7Rq/HUDMKUm0ilMjqzFCyvtlCOjliEy
rf8wvEgCwnUQlwK1XXhOQeZymmgALOX+gOEQg0c98K2pz3ks9x8nPec/S6r++auhK8tjk+tFTXuB
vnYrGcERccfn+V9Mf8C7EkIi6eJf4bq3hPzTGJjXduz7wi6QS4L78FCJFCRN8OtkuOL9ltG1P5C5
0bUsOuCOxa/wib1pBGmttPJcs7Bnv9H3JZ8Cx5c48BhaW0ZPlivBnK1M4tUq2TnwSl4ZwrHMw6Pn
f/sjdZWFja5LXz9VUxSQO1ryGZThyLDmQDG3AKoI1xFNKx6RpZuZDjZ9EAw/RwjG74KP/pzDchf7
icUxSofz39eNXN79kaOqAApMSvbMWgtGtuWxyDtcRcdDcOHNY68RfEH3ISW3Tc66olrjF29++Q7B
J6NKdm1peKpd4TuVaZAW8AhwxPhJ/LmbsuM1jWq12v3pWJxP2A2oh04K2BoTBO/5LmgMQiEEP991
1auLax+TpQwrIJGgI2pcw6gfL11Y2pQTzByQO5r7UnnzvOhRl5QQNaVjlLU783r75u8A62sfbd7R
pXcsb0BmMpOeX6RZ8a9hDRnX/5DyuuniGKUzbDyMb3OrgE2eBCDR/Nv2ZXLT/UQ8aXlx/97ntGiJ
mTxzvzBgA7ZnWWRyZsdaIR/XOSo2UZqaeYCVj5tEdfg9kceXfQdQbsXVAOjHpsolw+qIBH3Co1ij
Rn2jYWQSKfMFujMleWzsWsXxdF1luoz9BRPuYaxRIFXTwty5wUASYWDBHGXIZsQI+lVDsgaqSPO7
XhyS/GwuPmLvTW6uVWtIWaCUK9aQK3mXzJLTNDOLYiXtzYpvgfIKkewaFYddTwuMRlaVL+kzUZcF
aQhyJ2BY+5YrCdk+rISTiZaOEw3w1DTcaJpN4gjpeXvFRlC7OUAXfAeEh/+FZyTceOW8jHqfN5yv
hmWWy/qWhIXkbC4YHsz+Pmjm6QORobBHUqAM1+Pf8zgkOqCNDo/5cha53SF3nirCt1dY1y55iAW+
22HV01IYDGWC4brZzbH6eM5vuZsJDctPwhW3GPFXm4Ada3dQnRa4Ey6OoNOiivW/76LNvIkFI9kd
zBoSkACoHg9Y9/TcUAgs9h1QsTYlCYloCSd13PLd/xAKShi8uwFLBLlOsAtk6bNTuzCyfWuc9bL6
R2gJR4Bxvfr2yPJXE4LOmpC9e0Npf0SJvv50qz6iHCgi4jXr5jiV0Yf6hkZoHlWGv5upbyFKDmyL
tpu5xekbAmwlDzxtMiz5eZiNZ5DifxXOPdLXK888EZN11ev49aW6vlPWvpygxhq3wcGCq5zCjawD
rzeCGv0MqVNe/XRnI8kw4PY/jaCUL68WLqjDLwbkb5guuBYf6dd+Dv5kqXhTt+H2moPXxoUXb9B2
1MwIMPkdRYzkOmutpEndQxPb22CH8OcFRXwyoTUyI+X5sLdIThtaxc/e78HgAGN3A6SJh3cymSgJ
pEOerbJl6g+l1SfI997U36UojU8QQwrdZw2Ks02WKF8qroliMjmW2gHfnsFl/lFaL52jf+SwxSLj
qvTC4u3dJRaC/UBg0LCPWz+Q/diLLL+RTtxe3bVunl7pGTuUWxD1PZkxvvACMr4IJlW4bLcStB7o
fuf+PytnJ5Ql3kcdwPqUkRENBN00RexLtymBdGMLLl1zmR5Us9K9LUgApib5YEa9E/OVjpodbIvd
hKD+OzRO0Ts/1oSrIO4W3RF30kyFNJyK4q5QQYFuakTnrWPvvQgBZlMwABC5ix4c9R+Z8CSDE/mz
WPtGLFYowVEeXFGh+eHAkqEIJKxNF5EryzK/U/HM6Bhrji+2rEIFw5OzJRtt0c8T+HcQPXuXSVuI
20COWo1h5UBYU9DOLCTw1WxjXLSosdsEO78C7vX2zSiM5y2qrE6ObG7SARv605215aUFNO4bHefm
bLxqcMdJ8gb14baypczEq4GaK0jwIc8zh8mZkrg+9LJyHDyhjxDlycwgBe15bYEasnHfYiNn60vD
LdhoBL9yiZd2nGC+ranKbP2P8L8rVOB2a6OZnFnu+x5JhZ1fb8PlmXK3H8N370q4RIWOS8+BpW38
XEK8gkqdF8Y4kJs/RsgDQTe3RhOqm6859ACTjuav1U/liEDyuz+njIVq3VjcQKdpclHJt0PuER6I
BkfxDYimz71FmYMfCHyb7HdRt8LW6niXnMCia7l32qO3cCDFRH2mqrQTi9XXN3+Qc2wpzGOQ0prF
n/7whEiddwvkIFqgX4I9SfmMbcyWcOI+znHabIlXgYSM8Bol2J2FYiWhoASnVrz1N/GysqBqXru+
Ac6bjJ7HA07HeRQ72xN6TI5i+tldRS2DIRfvTG5/2DDgzvWsoKtT8Z2V5DgY9YFH2aqOh1s26xgD
TEPo4TtKI1SemNPLB3TSxAP2R/K4H4LpK/uuI17X77kE1Xrjtyd12S0vgbAvCndN5V5y8GxIZkDl
19BXi1u0rov0HFfLVDwMmd5UdMiyvgKHvQuDkJEqnu4pC1+MrGg+knasgnU4wKyjLVSpDOn9l/vO
nJkNYlyk+wZdKyCZHyrcdZQ0i6eWpC93GI5uDEPhKfhTv59d8h60cXaVj74o6+ECnYINE3Y60LY0
ASfvi1WjvQw6xopQewuOqyQC4dHvheLlQkLML0v49EOlaXN/+BGuZ0uGaUTMx9SfMhS6QKcocoIj
qilSKsV/KzpK46+WqbjxX9vFLFLdvOy0E+QWwAEOOGg+Ws72VKz/yg5oHD0cZENN9tSt0bOjUvaL
iC67hhXq9iUaL3MqUeK1TEp9GUDxaPSLn0HF/QRGZdGvnHU8lImMHZicrQeJw2wCYIPd8bqAg3eu
FC8I99jYtN6Mh0GmVwZCwJqiHhODYm47PVFomV2qZ/+QeATGb1RjDwTCrkFmzS93SyU3HVAEMgTL
et0yor9o6+46l3hhxH+BTIlPu+TzWeXutq+WBqoLKaNDkYKE58qYlytktlrWxmR6hzn7ib2yFr2J
U06csVFuUBSbT0HUmTw1JoChM+rAWlNUCKB9EOLI0Tvqm6o7EXoerNcS/vyz/o+lI3pcbLdOO2ij
ihums0zte2rsVgBCI1CsizTP4FufPmgKNlg1zHIyZa2QkOOtzXv54kmY5+d92z/WbpMaohSk22TG
8tLbjK0d/o7cnOoBC20Qxo64nq8ZQ+f4l5NSLJ4HJHjz6/b6B4FXtRnGY0gwlN6oFirynPK59qjW
1taK4u70IvzSWgLW847qhS0KclHNw66aY9bC7Tq5e4/Hb0ONULltRW4FNaBZ+sOGEEa9FNeE9fTZ
v+I/ZnjNi9kzUq/EdXpgtC5wZazYn4ITVfoQ4Y9afaiFA12spFRcnzOb6Y0+bpfxaCi23jw3BLBH
HRy5lnogXrKxrn7SEhTGd5MrUVRoaOIfjCHwy9ApcF1afzPpmwTAUZpS9MHKhm3eBeq02XfCzA1k
/o+M0ixapTxfvDy4ZYz8iUXXhuyGL7zZ/Lt6LvbKTbZDiOTBdFZUiOEhnXdFvB2P5wklRzQ5ZH/N
HSnBs6SYFOcUIGDCX2ThH3QkPBYfAV52ttlSFqFlRZSxT2FH4GuF0pQxE/YQ/Oa134nkz3nB5AwN
Xet47I/hZKW2NuY0bJxTHECaHCc7C2drw8+Xd8Vg9xqGNAreR8CN6euW5vUvvc1eG2pSLdDmAZc3
uPyiGyLd1QiMEj0DUVq1Hhf8yb3eo+RPWL0jPrkIHwMyq5dhZlPHaIMPzka4VAkBXqcCDxMLApOa
MQpvmgRnr8rX7jqo992DYZ4KOqTx3Z0U3mbMuCXtYThLxm8ykiLtYj7bkzA6C0GWAhM6PENfTnzi
QzJgfcB/vzWgZhpPXUhyImUzUUZpHVOLpYleAVq7NXogo6OjBXRdDy4RHa07su97ofr3O6klajoc
/tavS9AViMwJapSgJ7G9XL9b8hOHKUrOy5NS93LmIJvvpC1cKemE8oL9Bx65PttWyJzoVzHDqHFl
saxoe/m5n4YW88h7X7SDalHa9P2zbAA6xsp8d4+nDWkjVPlC8GJXbo8DuSS/T/phc3l25VFLtgsN
EVjRF/1Mytg5cKTVnoVEJQ7H7CKg+XaWpddl2Y6JOmSaYTWWBsxKL4HawDdIUEvSMYpjpOQtol3t
2ngbwGt4jsJe11d7z+rzBdzQ8FMqh0F3Y9sN4/6CB8hEanIuv3ouu2WHCRP1J2hB4hh0hVcTO6wa
OtapUkxRn3ygF6ogaAHXCi7oTe4bRYpUAEFc5RU+jfFxCZDmaEeUKBqCQ23dcMSZ2xQoaPG4J4sG
YiaHCJYA9GxdNaPcZfcnOiYgncKJs6Cvit3e/XnWMjOCJKMoHV/Kwyd/SmHDApb1y6rjn2X6aTVz
GHXLQDf+vJvPOYwaNyO3lW/UKWl6lqgOHw4iVeVHl/fuvFdNkaI6LIOd5fsIskOlSvbnc9xGFZGt
sZOue2cUUBnMKQY864vJ7iWgZFHXZpZWtqLmsOgurk6OlWu3mPJwUDOvNOPx07ezakBHoLMjpvre
7Tna0Fxg4swSli8XMtfzJahbVrZSY5/CVx79SuiLVd97apyXVrXTU7lwSJEF7i6teuLYTEX547bn
HCighJsMxNQfTG0Fvvy7o3eOQ5slakxf6ILSaV1er/pWdTtFIvnOp/m4yuNiwB4xiBC9lFvuZ37N
836N2peKnRCnnSp6J5Zw4Lqg2JSRbR9n6CozhP/ujPV1okZ+K0yY9lvP9Vczamr9Yijp64N02kw7
Zsb+6abiF0eAU67UGs+MdE8veBUKlzme93rDr/M7G5Y93IhnfvRvbZzhaTkEccyow3ywwLW5iYZN
Cyj2QIWQeqrYvSUcvptXSsIUpoMXePZ/NBt5y8481i95kQJ9BOSlmD2QK754Sxsq6eEnnVRsingR
0lL3FYSr9n4eEnFRon9iJNvovIhCiemxAWdzVHLvobroQxEzRDFY06gIUUfOlsVqjrWeULlNb6hp
kn96e8XWZ+LDq3yAmhHvQLHi8Si2YC9T5hE+j9hMDcFh8Dg9F6kSTmCzNvt718yuhDkfxHJw0Y2l
2jjqwehzHpapUOEZi0QLSqknWBO+zux+x/P4O1KTuPUhsL5tXjsAHR+bVPoIUDBk0BHOl0szuwT6
Sqr27wIAwYySX4C4+yafAyIQX9qId6bJ1ozTCJkHIafslVzZmtnFjtt5vOlx82SsasmzllE3llW+
oduPHtDYBZ3FH4jOJVt0nvpMGgYY7sfCFsj0qt2QxB5IH34O8/MaZrfn7mEbJZ9ugyc/N+UdsM4l
f6UrLdXSQoOa2wFLtIZlI9lDaokgGZa4Uws2ci4Bpt8zcbEuKqJ0eB+hrodZt4VmSkOFjZ7fFELE
yVmlUY25Azh7q3Ol2tPefirb61JKccGIkedg5YO9vBa1Gx5ai2WKJDyo5yqK2/3q9YYYX4DOx4zf
YFide7Wi7hmL4k/UCitzQ2suwPFInAAKjk5hpmVPXqBFtlWYAPoJeZ2rtRlSMMf98MZdDBS7XKPw
UpOXUP7Q0yKvce3fDauN6z69CXsX85PuXagkLGRG/wLv+n+nO9eIBqmwS/3ivXPo9ClXfRVrGGuF
Vr3rybZZV5gfSabn7B6jcFJCAZB8LMs1/femq+dYSKiDgJHToORzp9pn0ITNRXK+XqX6bhXZvTh+
X9LpncxGo1+JZ6DWblH8rmCsqfWv/vUx9vymZYxoMVcNVrlin9DNItpbUcKT5c4nSK1fFQUJE0F6
8vqYLlfdCLguBagNJzMwPu220OJnskG+/oJPMb9BAca9S+3UfJgTqhb0RXllGqV8GKsoJwDLsJ2g
CzD8k60085k8QeUbQSLeLv9WcEVIDVqE6qugPOR2+2OODV7sZD4l0wxedQ0mQiYTXYkmAU6ekv+K
AFB381WpSdoWXiCS8+8xKvIcLhezwlHOeB9G68zKzuE8YpVzU08nSqCMkgg9G9KS/PQKewTxRRAc
HkxQ4HuN0mJb0IUOKOWcl600Nj5RuxHC4UmH8eLh7x7IWNqkVBusHD7gE67wrc6YAqBu2v+1y+Od
h+01Ra8tGKrYdnvEcc8RRZN8ziFSKbsRmx6h2Gzq3BbWvTRtPrB0XMzVSzLFpa+Zgj6bXKZYVGVa
+DQIkd+x/3VbSRSQNkCC5J4RGLn9qYeocjjnnC4Qu3t+Xrr1qHLla9AmBeMFmamI7o0NiaLinCVD
6UlQ5sB0Sj9kLkG3rQ09tAMHSoq/HLrc0SneSniSTGgh9oeZUGYWVS3ImjTvsCVk7oked8bJ2mme
a9JKiKk6x5rR73VOIVLGifs6WuOvDFumMrD+KA2tBmAw2eVuqe0WpP2TPUHFP0OT3ssR84+8y5EP
tEjouvFj5n9DrAntCLdNn2Eay9aaA3I6N0DVtobZeyGWbg5nXJlEuSmzxfwnqr5tWJ40AStnLovI
roTKFKnswyYeWvVXvolowCUOgdKfFSXGTo4H69cJ3b2OiPNp/13IpU9vXnrUIsC0LrpE5j82a8Jd
rd5VKAoOFlzClsKiA/LykXEE2a3o0OvjL9cOpeeY9HpmvnHZdqfMz1qnuaqA+nShmiBTBvDpy1MO
TngHW7hbj7YogMn/YtazKjon0cwTYandRBQlalb59UQM164ICdKykFVHhRLVlYjE226zv0jhJ1MV
v0/xklByBmTXWEwU7QJvrvcrjJ/U0Jt4I6M/zDBsvKUq5C7SdPa9oFwoAq+CQlY302MRo6eO9Y1X
bE3nBCygVsqrEiO+ZHoxw+ovcgBKJdCkfUVeUxYPZnPdIr2ihcz8f99bhebZGf/WQnb4I3sb7NuT
VJ78F9+PPRw/A2EkAS2aaMJRwjX4Y0gsXx1COFtNCj8V1AwnOdUyAX0t5RC3jkGtcNX+NDLGvVvc
x/PnX0vbSNBpKQ1StDqmpeB6HpHcgAfngEkPJYxdcWzEAEN8x/jaqaIAiPxCbZyvMpiWYdM0HHGP
ji77PGwvdVkDVpNitl3eCZ8wFESnVk3Bm0u7VtsoNJafRpl4Ni096DRjTgh02/aNYgIar4SgouCo
idroWG3wqdeTgjYlrnrLIAxt/Li4iwsxawYTvdbH28QNRlfzsEjkIA0VElkNGAKF/2UJs2cQy0BL
CiOwSmdYRSGgwbA/hTAFz/TvMAsecaT1T9udEgXJb8yGILvWl0TZuSnFFa9jHzHrxdfmuyPrTbOf
ezdHGdMWlbGeV/1QVSd1yTPkm5lCMzOpz7dwq1QSBIB4UqOZIQOjSm6Hdbq1C3ryNkUX7rU+Gl6R
5ftaMBCrpYYAxrcTNjXsJxdyQ4BX4UMMBXcAUZUKTc3f8cZF3iIqLB/dRrkeT+hqLtlKuYrwZo4h
pY+IQ42SfRdp2tuIUof9KUIt08EhhqWPkqJvDzKEIiZKf6Fb1VwdQXQBeBa0gm75TAr98PvUFj8Y
3QAsO5RCb2S9hdwCQJ6luE9VaGd+KqU8YUQZf9wiY2R+1K8vBuFwXAQMrCKesr95JxJ6/fXzj6qQ
815p8ylcsJKOSnLO+P4DGRb+kZS6wtLR/WyBzatA9nyY1DmaR9/9iDvEOdkIpRWYgTphrC5hckKg
lZiYh6WKkf0VxbrlBthbAqmxheR/QHb0C1BDZHEwIK43TiX+UVXq09MgnDl4iHPvG+Dxuon6ORyA
YV1/SU5e5apw355Wc1g88IrVwrom/hf1mu79Gra7iku5/+XRfKtnQbN3d5D4J/QE+Txxu6ZjI0Im
pehR5Np/VRnMT/sWEJh2GwQilQ5juFxO4GE14RIGm3/vnU/vrcDoQdtM1GvYAg4ZT8uHwFxBa3eW
C6rSDkw/xz9SxPgpcDbvHfgWl/olO0nC7yd8HjIRZAGUPFG0P7qm7m8CMKIHilnRzrAENTQNUZ8g
Q39GTRY38maOfJDn3jhjYTSVFSmyeOq1VehwbaINDU09eG/I3bm0TKKdpNMQJa/J8nKHubjjQTFq
cdmCQA/ALwomA8jGXskWSds29K1WJTuBo6rtULfpU5VldtgVpucg2p6IFHsjcm2HRX2ELzjI40wy
k6F1kddmNI6Drq5zIUhV+K1AJ/hgXz3swLjSVqC7uPpiV9KLTqslnyXbMje5eKNYfbSbU6HiMzcu
aDO32KFzUQ82qGeNLPN2mmlk/Op79rK2JjAcJvewvCRi/3VIjoc1Wi6lL5zIacWBG+zyX513M62B
j0O0R3NZqZhb7lGJ9ztLAS6xJCs/vMpQo1ySE+D08wPH8oajIxu/zMPbzBeuVcSIavfnoloOwBSJ
8W4S3ADPtQC09lWmlXqLewKMuE4C/ob/foN6usW54/TaBNKrJmQ4ZE6CCnJiJpEeAqF9ZNGbqJWj
YFoU4lalOVUlbiJ2Mz4+1GwA/5X6G9MeA8pkBA7dvG+nzAuwlLk/mfu4yXXo+bWX87c0gftbjWje
uQZy2EtvhKtzT/vkPi7zN8xZNlazNy9gB7XGZj9kyjwGnnAbBhiSd449z12+OWcmKBvbtLzFMYj1
oLooXQk8OzQS4ccEIfoD14UcuWZeA/9i/Zzd6jKK3d0Tk8Lwcc318ntTzJ49mUHeSA0WLqs3E2w/
A3kybAjuy2YFzfYKlEyurG2pdZwEMOqKCPLJ5amqIVEZ+3yTOa7Rz7eNlARrLCiTeQ03+aUzic/7
sCcGImK4BGNdEmO/8hBj+qHH3JYyq/SLrlOHvT2Zrka/vpSdWinmk8rvTv4mkQujJ5Etd3XW3AHk
cdvG/yQyz3xwELU9ox/BCO/hNH0XbwY22dp6Mhm9PEfc6gGFNw/TLHtgb//zRGjor+QaYs9jqxE1
KMqW7rIj8r259k00a1qU2xPm6lR+pQ4fSv6xRh3Q/ETYJLz9mjRLWN8IMGQnwnEQmImlBriStOrv
W8TlSrxMVOLzu5cq8r6UYvBYZYUvNpj5xiQ12ytlajtLkNMjURWiUSv2sEF0i/OHJR2wBfkV63Ec
XBze/ltSol/58r9wJNxweESLf45rqtMCX68xqBuLyk5DTE730Rfqw4EnhyAEyDZk9bsd9VQ5CFUg
o4nLBN3s0rmUQXTA+wKyKVR82fKTiL3q6icVSZWWF7kEFTNZznZ6ygXQ3EzMxDaftvD4teOv/q7u
GBW4pgp40p4qg2Irb5c7T19gc2DaUmaANkQJ0s+fMjUFNBD6FkcQ/+eu6W6X6cOYpTnpgs5y/B1c
qPPdECvU283/DN9oW4H5Wfo5xdH8EM004NJlVcadjbP/Q/LpOmpG5YF7kBY+fz83VUIAEETUBcDo
IEKOMoyaMakGF3SiLG/o0lWeuwztkWmgRlEmugbmdcmUvcw/2Epj/IBKj5iVaCPiwVfAb8Op2zlw
vRZYvabKv1toWIb9DHjU9TkWLWOIDknBSmmnC2dHClf2U+WzQyaeOPL8pKta91aGEvfNrCoydFOf
JMvIM8laYiqzpcK8E/4s+J5qgoXyY/2NuwVsMccu/waad8u1zaatua2OJ3H+1fUvHZawYoK7M8B5
OFdPnvI+udwXH0LifTP4zdnoTgI0//Mb07syIrNezsvCjSN254WvDCeMduAtAhSM3W78EKBvKEVX
slxuBxTDCHp3kkiBNJiSc7ch0/wcF2St2kvqggAIxW3slmm7cd/oT/b0lgFdqunDD0cPxN4BgWHs
JjuU5MSRgUqn7ow28oOaaEkU1lTDlXO0ojPsFPjoHhqetgh4K1BjP61BpNl72BZdpx0+FTiG3srY
hqwnIV2v92b9JpGu9FK4Ecx7GDjXUeT6tE2QFp13lWEHVc5N56LSqGSeJjV/XBiV+wmYqn//e+I0
C4jUjg/ohavxK2qaqrSXvcTaOBbYmMblZajOytL3aRAF8qgPipbw3wQgHKtNPQVHVE/M2I7kQWqP
GbH3XIBUml4UGa5ApSS/dXTm5X19hYHPk8zGG5sB0R5ezNBpX8FNDJkdw5EjiqTmRK2x0oC290v0
fUoinOMSeUy+4AkryFgJ77FxPf/N1NklQqw9jMvFwi1hhF/NyjpIUlxpMMqpAS1U0oaZtyIGywMA
5ZlEWfpFIE8TeoA4eNrnGYZ0G9x4bkiYXgQm+D4WCmWygrlmuNhokfRuXHAx4DfB0pUAhs7oPtH9
xjWjN5B273KDBxVCg5T83AcJiKZuDqexzQ+iQEHLY0/GHP8TRLdoxmTbjXBC5EcPdNm58SJpNIYr
TN1nSN+AYAG2k/nBouy57o0X7rkTAp1vx8W2g+FgY073DOW9ryJXFgB46o7sNmWiynJzs8ViGpMS
iNkzwt+bfhNkyKAQhTGDiJKYx8DbxD0mGVKKPgz3fxBYBPVMzTeZSUADcOSNyqVILk4HNBFC/fNv
qy870zlQE7pHOZ07Y363BERAXUd7L89JzeQQMiKPkhmzAr2Ipv1sTmJyEfqG78lsv/3ojPChl6kD
/VC4A1NMCJw/A0rvUBprFJ80plFxdR+Q2bCD+bSL2JdjB8T57948M+DFjmAMpc9FFuYiC66ZoUEb
W7MpSu4D31a3n42WIjwxRGpu6wi5Uk2nyPv9fn1Wr/6xQPIMW5oMowK4J7WlsNgk2IHUCQ+HzCnw
yzOGF66YXyR4xb9Xy5umOiQiJr3SDCWOilmGQUcIltvzQ+xHZmfoe5fj4iKIPETb6zlJtS/tx52Y
DGpjTYvd14R5MCbL22jb0PF5WMYElS4p9VBsPemNMPLpTLuXqodODgIxPXJajFbU3dk2tLOPijUf
cOO2vzdF2u5keGYqs9qMHeAnkOmk2hgFgcoXr2plvUBk8cK4TVzUJadIQkMOekts62M9rLzLP1jd
3W2qZkKS4g7Q1e/9kgstQO7ZQ++Oc/wxVpaHsWXB9F3adFd2l64FtLh2NFzCWbAhKQJc3s+j/9He
7njX25J4aUAe9TdlMmqcrQdkY3WyFSMzRryTwmLsKjeaVxfFLLmuD14rmO1CMWVMmPVPtbjkBbeN
SoGZ+PSIYxowVmdWYH/ewUoJfIVUGXmOvYMWH11Qt2ERRGPsGeLy+8MxWu5YZAug8Vh+e4ULmK0t
00MU8BLbJFKfmhSm4RBKchvOHaat+hQtGZpyPg6J6TY9Svh4aOPQEa4LeVzasgwcT6nhrJ/XLAxj
2QOS2c2GY5SItbclgEtml0mEM6qff/HVqOTwDvAS8hMR8i8UP4MwLWhjtsK0eaX5qctxwZvwz2sE
bEA/dNXt9kkJ8pLjOgHetttTmlT9E+oT7Q/EfWGeJaFrv6cYIHK68reTIkgVV6eKqlEoMAN6/ow4
5i3fftFa2xomrEp5kn221uH4+lFxni1Vpp8MHfmYg+hPMW9D6ai2Dc06ciwIFMtvGmvknxVZ40y6
xE6L52Ij4WLwVhVYKwvoql8zoze9aBfBepGZVY3JL+TARlbOL/bn5DBIBwtGUxa3GNQ8SuVwucoR
P9R3/JczoX5c4q747dmQxorsmpAqZdY7i4/DDldrQIVYOfc/WLzSIIg37Ina2W0E1JnnMoDIUvZP
XwQKQc7tuQfENRFYfHgr7CfWYmw9Uup0sEmDEqzTbiCK9iXLXAkSCOZiqLDKjDTLPI6tPXdLPwlc
VoxbZB1eRrZ2QnXN3xoqr0jyQ8K8c6B7nh7a6MBymzqeunrYYlG71I2UTtX/wS9f5dNs9VvXM7tu
QWNi6ILGxfuXCM5VOWySq53ogeHRbtcvDzjeIJvwwlPSxICBrNYlTo1SAF24/mWkc4oed9Wa+6zA
gOJlfG00IM/Q99uWjCI5sVRXRXmaUb/DIcxjuZa5Ck8MgCv1ImLIM9i2fBwJeLV6R3FMdNzqFXIs
Banl4IPmH7n299T2Vpe1Z64jEbDvPK8zrN2aKgDEMFN5W+RFOgBY5rkrqqAzc65m0TQieuwtW6mq
inCRY7UGu4RyA3ktkfk/sdYatGtbJvh0wwYTBZUpVpxaQsLxzjnpI/Z+PtZCcaRDHac+BI551CCz
n4I6l3Xn0NOIqFd3sEikO3zfSFsHkKNaJICCIyvERWv1YccAFYJhD83C3uILb8k04ed5Fi8q1VKF
d5Nqr4finj6IAOihdklAqQ03rzqqMQ/GKIPXvajqtKcgBpkPfXU0lmhbOzHZdJ1kZ6BKWOZl06FQ
SjMWyrwO71/5B9itMkIoUncu3BeSbNe3eqQ66dtoh2IldyMyCpm0d9qhS1Ajp0q3L/8wDglj4asG
5dmo/hlBEdZPNXzeppQ22+xWlIilqn8SWFTH37mHOxYuGnldryDtHfA/u6UAUSNc5zrSoKWO//q1
cwFHyH9XNCrV7Fata84uUv4ezf69BzyD65DlrfzjfpEnTni6nuoawwYWDiOKBIO6zjpgJMjPenN8
VbEag5XiykieBOwn5pYnSf+RdP/bQeWUQORKNYzxTR9oBSi7CefqFaKLrsmu8QLX0y9VC+S3BUoZ
QQIZ8gyt5o+kcYA65hOtuVAXxjgtkneF49MWgNFDE7VFhqEi0yciRNCxpp5KCDYK8rFIsICPEYpf
NRq7fkdvU6vFgV1RsVyMPr4lOQoIBlcorv9ZcqfnFd62lImT/SrmYi5NxdiMuz//YEdUJTGF0uxc
kxX8cLBErmSrJy7x5IKLG3EFp7h+MNf79ZdHdvPbo0O/U+r3i8ig0Sz7Uq6KXjNqJiw4fSActaHv
fxtDQEKZk6NOm2efpxaZfyX7r5mcZdiHBvJsE8WCYAKF2GMp6lNGdtZSYVtHtI7YudhVvSwB7Ggk
XFWGRTcLTNofWF8D7KLgZcaFRyeO8amlWR1iFewevs3Ya2LK6Kp+QP0KzBgi6U+ldgmUq8O+ddsu
3cKTroHu5kAVncpzfEb8fFKxyDiwqn/dLMw+EC0MMtz1+7P7ZKWFZNU8X0yxRXUJ7OZxaWULlddD
4esxSGcjRqY3Rhf1d3nXDXqRhI7wPe+YeESLl4tXzUSI/rVauoK9e3qQzCIDqFwQojxnrhWvRYHe
MdX4MdJZWnoUUQO+8JDgh1aZ1CeanBvLMJRzyLn2X0b0wAMqudj5007kz8FQjx5YC0BiF3RriDnF
LAIktoEP/r80OtxPqwRLQ9j4wBmbG9SHGR1N+A7tQm7GsNfdzWg/hc/dN5Af0bJ3yimfX2IW5rKx
8Q96qnBXYhzfKbb45fPFl81w0usW+V5eFNkk1pOgvQRYEfxcKnFiDlNMNFqA7BbKDuUqGjAAbz8g
L8+BrVPMR77iBL1N1nGbILBCYeNR5pn2YYuXX/Xb9e3vfg1CPjcMGm6864CvkHRED2DS9DS+7hl+
ZJmhfCraa03H0Ua6yJC0JxRzBGUr8i6XhnRrMaGFcAV4laD+ab4wod4b5hrF1QVOkJ8Nyht24W11
OCgyRidv32MMKjPI3hMcFBHXOeFaRGv7EtCgQ66ZJMrEmu4rhgmrtMn6IatQE/73EaWWTcdV8T8+
bjxSuSiatQNIIx+fT4lN6EFHDc6Q0dJdr30HSDkJFcDKxskJs0uzAjq4J9Fhsx97Wy9QHKeAbDiw
VbF8lDyQfi2zfWeBpTjLXz5VBAUL86MnI80OI5AxCHKQvdwaD128pdCwLar3ZX0IPRzyxWj2Wn3p
6n35hk2e1CKl+rQ5J+C5QYCrGQ5O/eCyPKA8Boy+6bKSJzqWlaIX4DC7/oCMby4OeYKUuBVpKo+D
z9ZIfKaXJqCwMSxb2gZy1ka1F3bNCMbJNGYQHLnKrvNxLB9ubeXMy0MqdEIv7tWF172+g00mpF97
esD+H4T1JdMhZhVYrEF7CwnhytyA+bQXqXiQP0/CEp1R7IwDWtnth6ZVsOMyk9qWVXTbnAt1+6XG
hc1+Epf2hOsquwwJxgVqRcStlZV0K5W2AfloFVg5NR8MY3JMGs8nxNBlizHh8+wVmdjiuBi23+XL
/kthDu0yiSdAhCdPKXJGXxSUgD3TKQuAMQWkYa6pwhagJz6bEXC9inUKzndYG2SFRywLui3HqjsP
u3plbgKQrTC0JUsQEsBASYm9yUR6JS19tqif94VmeFx1XUQEoAsy1MFE8hMZQ2ZLkRu+Wu3xFPXM
Oz2Vrc2Tp/khbxTzJ3UTg02aFRPOAyhYQgrks2DuZRvdbJmEUZIgY2+NZBYIJjYt3pc/f/sPnNuo
OxvXfOzCZS8hvVC659a62+oywIasv3l6MCPf6LDj+MNZKzpwE8yb2kbDhf3yQabeqKVpdXq/gr/G
MTxqvBmGb+ZS01MNq/PzFYCobjOixa1RJbZ5pUsx2YCxw2LSci1sQlWKuTZOrvQZOOcLyZ+8n8x6
QRkD3oGjxWn54sXwlVI4/RtjYwYGMSmyyRucHP0RF0spiQDhV4YY/f+ADQwy5WjKZ9VZQ2DNF3yF
vsytL2GADzaa651sXE7klACB7FIN0rxVINDpOxKo75Zfh9yLAOsPbxRjukIFpCSaNpevaHP1Q5d4
2pXIUpbWvBgf4nlfBieSh2yOHI7u3FZwEuhk9601FK/uxQ4xBeL2uJLMVYN1Ivnv5ltXB8yAwHAl
mxAcCpkoXW9Ni4yCVPu6rFwWww/c4+TTd3KvsKMCFIeQaE7rUegHnKlXMT01y2xJZrrhEYTU4v1W
K493IUBd3E0Ng8jsEKeLniN5QqyEizNhse8LSZcASZDJ4QvAlpfXZwb5CsC0tqYXc1/W7mZQyT1v
hUER42BHtRtLRQluh1R3AKttLaLJxHOZvZF2mVRzyYBEOsTct8ZkeEW1KlzkLrZ3Wm0jnUspPnOT
VIp+owuJ1wPBOjPT3l86uZrzk2/8G6UbuvWkyVnNn4nHebSJEqOcxs2Md9SAAMlJqMrm5jqPsCBG
hdVzUQM6nxitsblVMThW9IcYTi02QM983fYkER1ImY8uIjC59INvPiKKT7cIj1LkvjUZXqjBZqDg
OrJcJwzREiAp57zGY7Qvj8kZwEjAHLWUP8OJVmAf4yv48MBatwYIUhuxYDDTArVsb0hRWg06GmlX
GiAU5TY1bzkue/ZYbs0Rzg/EskOtTk4UixjpUSeuCFDy31dZ8wGOJmTkHuhQsIqBfxgbSNIn03oc
DMs4vCPM50e+8rIG6sBYlx80f7qSHVNJKbKN9PtcYOZr/vhvjhME8lo7rQLk0tG1lyEtlRe+gdnF
DeNDrniERL1IZlmFNdDaZYouaYcP1fV1Ff/IUO3tbSlhzhaQOR53kHlEb+DFvq4TCe5vniEDBa1N
uBD+HvFVOIKrTocewgqE9+IXjF6etiyFdGgoDT/eT1QOPJRQUr+nlVUXhsQOwFmp9PIgsCKCizrU
39xKvcLuZRNYdDMOpD8T75CDS9bjv1KFzRGLVoN4Bd8rLtg8oiU/M7K1HA02G7xPTZWIjWNTFmny
3ZqoOeb+g3x0i3REKspYLLvIi+WT1TUHueAtY6Zz9y5IiD2H8qiNK06o30Q5o5u+072tGE0Juaf9
0vuN16jH3Ku5/MThOxoVUjcaQWyLjmk9R6IsIizjOATSMmwKFsLETqfk4pJsnXidMAhYPFjW+uBX
Ll7kcgQMI+tqfu9pMKeNeYRqOlHx5bD07468UgKtmPd910IqvBY+TNTRhnMDbrf2rlybBa1M0F4g
/Aoc3/9XTfzQQN0JkU8uziQjtTY7zeBfkBJXlNKabwpRq7z/b66kL1cyYJLgqajD4ayenAWpPuXY
63GbPfsYDxEQ2EyC9E80I9FgpzI2XIulCW28MoruKybgLV9d7PKoa022YwMFQFg9m6WY6gWg45Pb
FJ9s5LbNW2b174/1McV6ooc5LvRt94WDrdmldy4C5mc1hD8/pNWD0Mea1wt4MntfpOlWzYBT1E5n
M7k4c/d5TLLeptN+Nk8g3V/bIiZnxaPE0ABi3BxozaveAK+jcu2YDaTEHD0uGgvaOz86GHKOwMZU
iqzhfLNfEZ2WzqRcynO+MbyEbffcbmZPeHbnhL3wpoHJ6stZBvu/sPMXX2vqeHY1gSXeCwjWc8CJ
bzGTzzk17chKVvuDUXkLz1zOdumatWXh4okkAYwd2tm+xWrvIY0Jf7UgBj1yvyH7LDJ+WA2wQ0I5
HVn5i9fSaJwAOIUfXBENdXbeFYF8uWCiEoOXPrLqqKhw2o323Ldj9m0/HJ+iIYnKj1r5LGHNdO+r
3sZY2SnhgSLwcVcrQWcJuMp7dhB4/Un1YRTZQ5UQ7OVtTvCGrnfRL8OzuuXk9czJ2VuYj3OprUre
VQnIBg2MaPWq8vHpT4gzYefGNqOMVYZfQQ1lkIG0iyQFg2iPFvTzlu4paX1El/m9P/hegxxfmpG5
Z6uLb56YhEFD2claq86WSYelmdQWKLUWJKacPkP/0iBOPMz3SeZCRvRdPSEOm2tbeFLPSZkll7ei
tEKJe8Kn2kt4YB2QcjbPwSbf14hR3bZqRKTCVVCN4ym8MswJ01opYye8OqoIvyB2vZzce8USPWmB
U9iE7KYybteFzv3260Mz8wqBAXDLCB3MpTsvqsdnK3l3Xi4Yb1imvIfPrb41nmTUknUQv0+RO05j
UFoEVQTz1dCVK0y4y2RlidXB5YDLsyLrxD9hDM2GrPVrc4tSCdroqDwq0dIAZ8aHxglk3kRO+nfx
C+yEzTjQCqDzmqJQAphvi96DxM0UzfbpVYbIJHVwP9ICrUSPebaUQ50Egw8ZcrXY7UWMl0DxYQjR
UZd1mWv7NsW1qqCdhhQc1VJ6exWEA7Oy5KcUYP9pwf/ru/S9hOR+ss4gYS3imqNqJrOqZDZpW6u1
h2ebWUGLgS7/ea264P/2sMrAYIfXKo0Ma2n1KTYlJnvkydB7mlGnmWMldHrzD/sJlF2rPtda+kLI
chvH03YE43TFAm/HgDQNCC2cf5tM2CMoyspLO6PG/UNACdCoDh+9mKHK8PDhNrVcNYSERUSnU2gN
pvkVoYK5Fz5F28kONWmrvprAsEObe4uNRhIDzUsBHhne9muBm/5jgKRdj8Nvaoe10aE81bJgg7v9
jChdIJPIUd8EORPZf62LXIAdimYN7a65WxtdQ/Rrj/ylD7oUrW1fX+4oJvWmpsUVO9uHjs3NMo6L
zFpD1s0PwRhT2fT4AlC1hcksEiU/cEo+DZw+Btd9JC0862Y1vcEaydQrPKn2VYotsxKqNYdGhQJz
yiJhOusMXXOlwwcsHaEw85HERvqFwON+vjqtAgLlC16QDlhE8PjBrHZLMxgpgdJXTA6isKt7OuWo
B0KEbE9z7V4R43HbLa0R9+So1cCJK09biqMJG4RYS3zck52C/zLJdgR14UTFdO2Nfs/QNkJN2lkH
MtPzNDz5yEb5xCW3qUUu3+buCjw3rhC+U/p1VrhVd6LUzByomMu8mYMWmUrdtf1hEURBPdcVNqMn
WLUvO3tAwl2Z9JCpl9B6mii3Xl+6ALHwvkBNEuF7hScaeH31+uC/jxdLxXbJdzbPVFBRiwf7PR27
G4deyLG6K2T5z3TCfbjBH1ul2uErVa8DRRolmipbPZ/sMlOQievXviVFnBV33dMzo1ChPiJqERIc
Cf6lV1n2gvH6yBVC51/2N0HVXkz91L2mcY+rPaezFroMnnhwelpwoPK1cl2b9JaSuSrDba3MHkcy
7BtG1aLk27NfljLP8jWx8VK+9o6foSRKL6NCO2ut60gF2qZAvBXjKqQqUi9klO0mCdIaozytMDEs
JUOnJSzdq8pH0o0UDzfZHKvL0urVABrkdH8lA4dhsZYCQa3R5P2DSpcJT0IhNE9I2PLhhcbAz2zz
KClrWU4xmC5i672eLhie1lC1dKH7Jept8AeDxL6alFkkBe8HDX7XKkOCeR9WFKmwPtuWBtzeDovO
vjox+dC759m3r8F5u/662AE1xWgR5xNa5aj4B5k07alciVcCmb0xH4pSrYZ8cE/g6o51T0xphCEz
S73lcKwUuQHvrwDpzSh/xQjKTf6vmv4V02M6TLTMDA0M7HO2SqJMZxlC2TtFmO6/fuYfMGkh3W8k
wTCMVA8tQKmmqyQs9CV+4FkAD9b0MPP9WM2IE/4TfTeZmreADr07GMpHHXYQBKgvofQ5EhsEediJ
438EVt6+gQykFk9slWSo+XGM6ImiE7ml0Ndk5icwoCZa+2m/i0kVUkKtj8pAAjCfBmUkevOA0Psi
DL40hyIv4A7IE4ltJldn+eKwjBdq1UMXgCK5BafMI4Vm8xw+f+3WATvli8YbLMHiguZJntIuZmgA
av63df3BqtPneT+ugeqtTMOHY/jR+9CtwrksgglqfUbRW1kJ0xp7zmlf+Tlno2OtctivLX3BN4+9
UG5k5xs9erTt7vOSdBjKxqAfYL0QpoTSXBQq8GDEeBkHCO2QYcrT2QUH+aGkU5OlMZCjueedbeRg
dIvdv9BsV4CnrbO6ZALCSyu5R+rdEd1k1p1uNKE9ENB3lIWg7i6Y3J7B9tFlS/7FGhR8+iWupjw0
uN/Sz7JNvQJ/5UbzI5wQL++vShjyQR6DcbTzRAb+Ldqsp4hQwcpBct/iYTe6ayexz+Bd3HP0jUDG
LtuiDfb0qdibXAa3x5JoODSrn0NIGa76B6c2z1bhTJxVBkA0J2n69a2nSQxXBErzXbQf8zCo2p0x
arZqrdeiIWUAgM/ONM5qcjEck/QCf3w/9eeBgCZmWhed5088aN9yn0W98u5IXcuqklwx+WsoGwA5
tWL2Md//uxF/H0PCHxhIaHlwmRSz9jB3FzlmxzyUOlbmIlE5ej4KPNVeVC6Qn9JxA3/RSNbUeNmX
lvwf5j3QfqNSoljhFZSD6Yflh5Rm5FdH6ENCgMnTm/ZblDAN9+pJv8OOQuR4F9HdmzglXdba3+ep
kjB7JsRwTCkQ+n/5ru7zgvo/ggUMJEqi0H6h8lvjbN60tUHZfeIHRdCo2x2k//RHRB3oz99RmUsl
ohyqZDPwxKWFnlr6Cxd6wJ45kwHbAcX6zIjI/Ff+9YP6xTa6htwxRF5i4HHPelLME7sy8RlEXIrp
Qmnj+7F2khh9odn3zKfopEg9pmGuYACBmi5eSpVAVsXSYjyryQrdSK+Dxwgpr0bosdyiI9xQ+xXa
M1yZGiJwYvr2akkkLomaGE8Dr/u10t4DlzNH6IEcecLv10U/Z2VS2BrqhOtpctYMS9NkGSIYCLze
6Fqa0KeowYXKBEmD3jlaIQms5hLgKHnkI09F2hmil83lmpBp8DZBnkq1lDWu7VNVtq2bPTxnetdG
1vUUI4lieQW3ITA/fsl672fLfSQsyDNgxKGxUCCI8oasrtCijsVWcyIPqcjxmrXVfAFmeZpfr+ag
oZPapG0eMvxHUidE/QqR6uNAi97URFoHVys/K5OSW5njYzRwd7f8RDT4bnjT7vDNYnn+KiDzsoeG
qYpeo2lyP00mcBGdseIUuQa80IlCQjiaOxThmZnC+FTehQx9KCaISwf8mgn7wyc32kx+NgwkDamj
kSzoEBlVMtoF8bNGuzeGgKAjfLfVn1WEjAsvI0UWJvsOkNoXJVbKn8NHa3G0uto7M7qJhSYQpv+N
FCkmnnLBuJ0CO8RNqAap2Yu5mxHk+6xWeg4ZotWEoRbsbjB0EheL72yxbUr4r2/2wTaONLn07QTI
DcFkkFDpkXt5ye/cfadkX2I5ZZgqxKbFBn6QcM4hNOVUu45Di+hgEli22Pb3JnhAklWj4sgES1vz
yqPUU5ao+OddOw358l2kSZQtVokQVUviO0iI6cms1Ncq7ULO/IIl85ctPIDcfe7WH12AQu2ApW68
bF4mRouB8/a8+bl6ZXB507b2ldzL503w89aXslQ/l1tp07HpFijAX2edipqTjaKqI3uTcQr48YsO
1Vguuhkqs+sQOuByCKZRhCiORK8bVs2R83I0GJckia/TQqpqjznSPPh6xHjLcF1+L4Mtna9VUi0r
nZT5WS9X2X4qcHVZSKfAv11wzG1hNsQXDihRhjeGLPpBtZSr5OG9/iUV2LNVkQhJaP7/JaBL7QCK
xaDKjeWoHNAPZgyTBZR+cHPHz9SUpjvmNldOuJEJ+MIMTWtp3DrFDWZ0Qmv0IrpBxPbkECH+5dFW
DmS5l2qknyRMqaptcA7auS5Zdes/D09aXGkIicorsiMHKjViof1LjFit0ssUFDaPjNRUVNE+dd1t
KHs5lIedBh44O5xfGlnEbKDLmzvkoSNiSuBGyz+05MgjLRCjOcJHee0HYT900h5wCWF6SXWmK07C
qwhFeAJJgNlIpXbHeT7Szrhm56gNwrt5aHUI31tjQvIOGgRlXTbQQO7lKmEDN+8hXpy/BS4jjcox
kCVBkuiVUjtrHMEFMZIAwc5oF3X+OGBoeKCyO0tra/wT+yckSN0ALuPnxQzB7x8MAgQrP4BXwRcD
uWbdrKckoKtLofvFKUxOFPxeRAVIjq1nZaYuaHQ2x4kmoXiqCKh4pjM9DWX0mfheQSZDzoit/IqN
a8G50yh+POrAUBABJhsxCj4+Uqrxbgpk1Db6svudvmZO9wG9IxnZkV4wVjFlXgujgShwxFjHHP+o
GtJskocZwfODpGSgdaFGyORg1PBhAHj2CsC4UUUltA3vBnwhNAqWWUAjEIOaaq/Y9BzR34qX/jDK
jfMVZT/HPZ/mdDCnAzlmdZbg6fsq2COIfmZ04faEKYWAXvgdWa/lEmt9UMuLDdOzXhkngkm/2H2w
6xsaTv25Wdjk2XqhU7TpRRC4h9XQUQZbzupX64RyX49pbZpqlOERCfo/LuADWhoOo3rCVh5vmlet
447mDDeRKpyuqihZ1oHReVXoIZc9ZOSGZWXAYQqk1GX4GbPG/4bNCulpKLGSBU8PSM7XOZ+EwEup
bG8i8RSOZlkII+JaqTBzDCHFhN6VZPmkdUu6oZI0CyJWGnBJNqjNNAAbDEWSmbzAt0dMbiRxqk17
l+Ekumig2VBf0wgZGWgPJ1UE1UsYnt5TIJMjXFA5TV/wG25jUTJNJkwrGstRlXN7t5XNJCwwy1oZ
nOHHh0TE33TccPsie/0Mt+bjNSEBc/LVaap1ZvCiWCzzzZH8l/f3QbudEdrOP1ND1Wl0Q6gSsY9Q
y9O81C7nXmOE78mf0YQfjYEyc5AAjHS+PXv4hZxy+RzMaLkyi1N86Btva+/6DWz7WcyOYo6IsY7W
p2L0naS6R21hFo741wS6GFg/Riuw6w7iIUYXJE05CScOIj4IlZc72jwpVIa6e4IXbbj3OW56vfB5
DlPHzNkOaAaGvNlfGNx8zZTv942ugadZmul2GeZGuJY3teG8Y6QWeCXWcNUenZ9nNgd8CD+F9z2N
aXbzhEu1hYfQHjC7nlrr20cBWvuy4PIGA7mzCal5dpIpfi2SDWAN5QUNTw79bFG5SX3VCCCGhuTz
2x9+TuauSfS/dGeCcPlAwjMRoeku2d380F2Qbzs7wB6hbouKrOQo3m04dUq/1dToNl4eP/BZCZ9O
/+2UAKpL8O2N6oYDaxZX+stgn40tcpdEVNmNoLAY1OygnpafqlzeBBNNgkWDlU//CA5lgSI++tem
cY55wRYQt7oZb5IYbPHf8sKAgmQt1UT3Qx1KpM3ToVLSCblZ9BP0XTsPHNJ9WhGMflFNG3cqmsRY
XjYvKqHycoC/a7elAZYtFljZbeXGiGwQviPJ8ysLSOj90MUmJgx7OSJ1OoOhXJxOGzv/hIPXJquX
mSBpiHiMb1X+BmFNDw5neYGMMcB/eQKcanaZsLZe5Q7SqMIKXUTPqTahLVBFSf4VHSeYincjYca1
KRDRGivSXfS7XuiKi0a+AmN1P9nLEtyVnBpZlzytknOpFztjlqxUFH182bKBiIEwIdcVIS+xDwDD
hw4ji3366ZDtsC5TzirVgTJva844ReKILBiGg5vdKK107t7QRWgzO0cmbVblHsqpOmDSswHIJ6K1
KT9gpGpcYtWn5YtMalUCfvFM593pcbIOppQmvKr5OU1uJ8Hce+cHUVXac1KqlKcwOnGDk6lckH3w
nhiiBhqVl2KA7T7bYhOlXcxLuLFEWGKx3u12pE1WSSXIoXDJa5oTh+Ca5rfZlMAiWkIWHyhsQQzV
R8ZE8asv3ueGS/V2rmoIWicC6QgKAEqPWZuqDuSIFVckFIrGUpz9+rWnISM5SFDcep13hxjKglie
tWeFQnVaxIPa7rBEbzv3RPzZN2nW0o0KiFAoSt2dqA3S58UYXG2CpKwe3XyvKSZrM9A3+mThUvQX
hxEK/NDmMPQ1b9md7RKCne9JRV9BwziOBNJiwjFa3euM0+ZlipC75p6STxSd4ZqNq9XcPSr6RXkH
crnBBnoNasx1+i6hFAFBvnPh2CQ6+Gp0/e/SBM8BhCwkNQidASSLId/PdDQAsNOfq5RTe/gED+bQ
l3wYJrCR2izG5CUFtS1OGmpT8+o3BVhzzPk9CbirBBaGJPirgbsbsf/TjWJXVPl5zvTuEK9lztMa
G/DFcHbREqTcZj3pM9O9z1poP9GI5n35nacYnm4OeALNnriYbq6xAt1aouMmGiA++PG8nIUbmWQw
ENQr+nNQ1Sex/v1vOms5diI1gxkO+P6unmV30xXKcFLWzm5FRUoHSd87anN9Zucpy4Ed4P0EH/15
dOVvPpmULxUkpG3wMwe23sKJgP05pWrYDsrt5g33js60n6Gh1fzgHMBfkX/zo0NAqMD2brn0ZAqM
r41V/ffUvNVthJTFESRtXIfOvzybMFLxgpdUa35K7RppyvcORepYVjeHu36uDuTGowxM8bcTkI0D
8n9gB1s4Xe+bgVG6BzQRxlBjwiCspre6uHOqOMOgkLWaCogIW5F2UxRr/2hJ05X492WOM5xgABkv
Hxhi8UtCbxgI0f36go29SeFirpfpcw/yP+khkaqT58HpeiODxMqRwJ+swz2wnIT0dCw6tqF8TxxJ
hO354YtdHMZA97lXu12vF+o4fh7JviVk06YJ1bs0b8apDnyhsMDSFF2mrQvDsXAKEOPToORBdJ4S
ydPUe5ZHpX9xNNQQ7WipU59ZUOf/aTsYBro3hDUzU7vpw2/xMkdth9NMesIDmP9qecz4FkLm1SFs
kE3Ni3jdlcOOG4pkhGPQyKX5QxTl6QqhOVMhX346g8WK+LXJCaI9hCxYabgM0GJQbibJsstW7yXy
B+4/X30+hKaHHkDivuB3mYqZOXc4n299OG4OWdUP7GtW/8C1ve/4H+15SRPLcxX7t4BjHCTjdjIQ
HzvVbjD9zdD139h7Qgqg1F/4EQE65RTQ5kvYlLnleKdxxWcsj6z8wn7LKMloVpUkRE/Nob/C0zeo
E0jt+w//PWUXJ4Lms3MW/sW8sL5tqr36WqJZGeQ1/axFQQiXb/AJvapFZ3qcfZK5Zbs+LMHgtGeE
Br7lf1ZbDHhsRM6VkZCSoero1eg0CrbmB3MBoShxuvX/4gODe2Aa9yXm175ShBq/roQnukcesQ7/
hVzsyeodqp7Y7ibEL7/xnRjr7BA1TrAekAJD90fEHtfA2hC7fAdEO4CjsUojEiVTDdwmcAyVPT6S
f5rfK9/fA+62gyl/5DnblgxRhKsat29qzpBtzd04ojwsQWD8v9rchMzDYdr+BqDKUTlMJ+axAY5Z
rDmTJXb7GWvmbJtxKkk74nCfRfUZ56i6eaUZQIf7W4460dGlb02dJPLsrcZKw7u133IIIivi6hKX
NJ5rLwQ+Liz2jRUfU0fFBVPpJ9m0o8MpoFbPAlQfPG4o7SD4xX+goqONqPbOgO0yyBpZzdtCxBtW
QOivm/KLqh7JMxOcFsKZCfyKH9mJchZS26Nvnpf+NOwdEIHbTk2lR8pJtSF21nRqjvTTl75ZSf7E
W5Vsj6mNB2khyGrQdq7Ck1T0h/V2pzK1hBfexpyoilySezEBE8tNTZDBSCmPYM0f46uLTN0mqn68
de6FMqGBME2HXHQzaRz5wVyCC2zY3PfyTedLDgHywRJ8tFy3GanH1LIda6KajpEpjDmCgjHm6FAI
fsWIzGWx2ZXemg2WAp0KQFVUAVBYPqUJQFxNXVt5NAKd0eTwqBciSMED+8scxOzBKQ0O89HqMhWK
pXRqQizvcBPCMeIi+VY8PGFIfdHRav0ACnOOOcOr8dcxJoNJcvryD+SdEu8T8k4qcNl6HSYM8xIo
HvWfN+mXMKP8e9cpiQqS3AKSNwptfHCAPK5ce24Oj88rCCsOI6ZSu3oySV8ypF0OIFg1z/jvkyAW
tzI961MPLiwgGTql0WvVRNNN8QVJHOj/uxl+j7LezM+4l2srCjd3dFrefEtBLrp7w56eRFHHRcog
68Xbj6xEVR72QarQAwSSTDp29V7gfutDjlkvBLZnU94xuoUe6s2W8IfiIz5oa5YD5BntqNVKUK2Q
fHkbfnuI2pwyjItR+vpcZni++smoN0XaWAOhaxTqLvoDFx29/GPDGDRXmHn83dDIa82a033S5mSz
fBiMq/0ak6KGy5DxLb3oysh5WH6rtRbCvSqVzW5iXUmOfJxnGgWdoZaS+aWFL4rcufI1V3HYweqA
2AMLwFz0XRe0qpRc7WXKOttZ1aLI04AxEJcirp7x+1xYhcFEYba762mdOS8WG3OxRowJRMO5PV7x
O9fK+rY5xUMi6RzYBT4D14/WcjkcKapa9a5aa/LnRdoHY+1iQNPWKt2LzFxlm/Bs3Ng98CDpn8zY
Fmi1mlMkR4ldYaJC1awvpJw4wcdkgykOczvQdacNVWPosv1n45/L9ABErxWe7D3nnctJQKO3gCCT
9B3jdgL/nb8KRQMj7fVXnHWdNmEJCkP3uq7DBeqUHK02xZCtvTzB6xg9/k+jGE3su8216hacM39n
5l555B6aBYx/AEQp8i5SWgePXM36yUNOo3Aqe71UcfnXWmDehsE3//yhxyji3LuLPPHOAV+yVKcG
KOPQTgclc1cKnbsf9oo6sk+RwaAaklAWUqX4LEABP9UBM7dR4szoeKUkDmYxa8O9KbmAQrXBDBxl
9U+qXPZjNMZ6CpVIGjUWL3F/XKUYW3br3nCC7Rt3yh5ZDBxaUT8/LJPeJCaBjOscY/BHDZjEmd1J
ECB7s+IwN7L5XWhYDl3lsjqWy5KCpWywaq3f8xEVHsZGoSmrNHfk43R2YSStT/vScYx1J7XJBCbV
ImV3mZSJOBlEd1G3+d++iJd+sjBJMgbMc+zbYuI6frDbXvHSYolO7p+Kea5IfH+3J0gS8ypP1Pl6
AuQkcMe3YM07hkSpa+ZDCDqvExB5CNh3WYLvOnasdcRutaQbvPPjW7qal1Oe2iDbejkaGnA82a1o
izVOVaBGq2EKtNFcAyLoAnMA2I9vCEt1aaWmoecNziTf7s4BRj3mrk/lqPhJuVjIJOVzyrWRXFZW
8/c5z6KJWpyXZjhaJCt8spL7eu0sTFqisHsUjGtop1Fmf/S17WbgUgn7l/E6u/KJ1vCFrN2WijDr
tMm1jypC0tz8z7qP4A4PhcWGGKpInnzKIP/tfVfJ0ApX0HioqFWvZnuJ8nzxmdt5AoJlqyfLolvZ
QM4dAOYlvoiOhtDsp5COr8zLqihInVd8y501jl6F2gQ1D5MsH4MrbYISl4QfFVa2bMhHIIq6+ng4
cmzvNmQcWIJGiKzeNEhXRZ5Vhv5BD7eAAsZGs8UlQejqdy5KORYVkIKvsvt3Eq9uD7EVeP56qRXk
ZZwRscOz6OVnGpRtUC1uzMBgdhZWMnfM+o6/1ZOQOtD6n2sBzF/pAq5FoNxAbjMybN7jSh9Nvc91
AAFgi1dlSKG4tYKqCv3qBP2UctY5AClHo0fmFzzyzCrvyEkOw0YvaF8SRRAjCSDPvNhmxIJF4CPt
nFnTGc9X2pQ0EL0irjS+A7idZEw2BjKl+JRMCUUMbNCNCE3n63NWVl6uLfY9/TAwVGHT7Dg7ZN1F
GviiqpNcQZH4RSW74ipkOGOdU4HB1vA/UXoaQva0ItJbBbaXzhDYz6EtUtnhtUR7yHJkh/9iLTI2
/VTMQlqjNuSnOWpWqMktO83xX1VqF/bRP0rSDb0oVHpACPNl0EA7OyYFhvAM5TncUtLYkofVDuJH
8chPzYO64Bc0XgsyI1poMg0Wa8K7UUxgqDcBTatq9evj3Z4HZB3T/MulfmGBG/8KKSbmeyhuYLTJ
lNmKGCS+RFdxux10SHy8QW3p2xmFo0yI67YYz8IcxdBMXX9+G//IwZxdHtc8eIWBw5+KaKWgr46X
uOz+V9O7WLHz1xBgYqMOJhx0mDTldMheQ0zapvs/X+5oBD0Qsi6cqo01InTTCSrvgN0KKVUyy65Y
2Fw/lOhMWZVfx39Hq02TrXNVPfyqFfWPgUhGMY+r+fT+fQJMTwE8Ss/2Djrxz3HiJg1fyqqOz6CY
AB6BeIe9neJTcmU2JeiPh5ZauCeZHaVhEXx2ei/olks3ifPnue74fa2QHHz6aEvYbIF0KoXXmObh
zTNHAO4eKBC3TggE+5bGa3ApGJ94VEOBeNDbbBJaDLNjvV1IpS6OJrrQFhqV02E1K7lv1DYinGam
ySjXKrfU6vIOnHHaWOot7YpzDyzm2MG/i/gNnVzIalggofN1CGAbl3Py3CP9LQzj/d1zu8KdvexW
gSSXZ8l2Y2cGFQ4pZwR6raAXPGz6J2hwx9EL1ZG1qWFPINL4cT7jlylzPTtgTR02/pumYJN5swl4
9LaKd1NZ4A0xPNv+IWN1D/4nMYpLTWnS+FldRUSO4XbVAroWqrfrP1SOIDd4D/x/bUi+tcxdHCKF
Gz8ZJI8Dwbux4SvMoA+Yt7tfHprqPrVRUpboR1S0RBiINLHY5R0aDdh4gDYKW8r8EekbnBKIHY2i
yOrH+FA6buDyMviU39b+e1FaNiQvXzVV8KrjnI++vE9pBJkXClLXB8ZUp5SiDNPIWEAq6XfgjepT
GyExp1ESQ8AIcg4b6+dntjJqdQvJ/V5+GaaTgBnM3aNBYXOjLWTnJqWYNK7pILsQerNbZkMespWB
6aqlA8BUDhVeNAdpV2MPZ+7wLMYSylrXjbuQvMgoDcc91udayzBWalFsuv7IKA2ldrTZ/r+4jMC7
+02c+Trf9ffV0uqNQ8oISAPCOunHc1hB85p4fDrprzhXHBHbp05FJnzPpXBhzaCaGyrT1r8/Nxi2
GCgibKe26JLALTpdy6lwFXMQbhwF5QZ2KzWwOFZ6E0L1LTeV9sywNdNmhoQurH3qNNe3vCkBV0tK
OcLk72LOGzflnGZxJzmivLjrrwo58quia4XoPgAnIs1Biu1vQ+QOiMbHN0R2w04HbhepRf7W/wmK
kH0gWnp394NDZ60ffCr/BsOvqSnruilYtULBe9OLa4w45O07SEFj5C+b/bPYW9YQzx9sWj9E636m
kBJY0vlz50qRq/5uxSUCtXdehabVOY+XIicnUhqP5bAuqwI3fu6r8wY2WI0tXpbYG6FshMsVi1up
FrMh9r0RTmzo9Z3Yli2YGLDLvX5XPctx14zLOzY7qCBYR39DeAyP7y699OspXpJxrPGkbExu13WN
C5Aw5m0+rPoq2nNzKafN+VePom5Ae/9pYuzYzUXzgtymviPMwJ6t+9vRkUlEeKtKA12aketd5wr+
svinBYReHaZlIo3ruPc1OMVQnE+EfOd4YnoiWHTXo5lC89r0vjKEQKpd9QpCdPfYxv7/uZhnFDIf
EggvCweaPle/+EUN9jPRW0Ls2mBs6pkRlQ3Dmah1qSHBeGE8pZuAJvhdBxNBFvvFJRDeA+WO98+3
GCKyeWAtbwzU2bcKN+tIK312dcTcQu1qvQKBAqnb1/qc7XTstCoYWpKebw1QjWq5KQN/fupUX72H
uzAV4EIFGe7NdFdtMxuvqiKAD8KUtdX+btapXdPM/O05dWi/LqqxPpS6DmLkPDejmSqenX7UOsea
ewBk3HvVSNyx6wuI50mhHdcNYtvDuKdECo2mISPxEs7lKQWUdZAAiE9Hhi7KdfYhnvfE79eURAdC
7MFDoALxaEpgJcMPzhSomb9FSB2OmelShH8F9fwdCi7MC4hut6dmb5oSqFmR39WZ7ROA1ZfwURmq
JjBr8bGG5+lg8KmUfAMouWYyyMs4+RT/oxk6VTDlpQvSXNyi4qD2xyukbAhJpXUrbU3iEob+dQr0
uLwXA4PxZNyrVXkjn0oeRv0r/Mu914+2FmkYE5dJn0LFFj9ts8SAdLt+7EoUXVmRp4QVvHttlJSm
gWJk0vonZD0NTDndFz9TuPiUriSqM3rC80rnMq7TbNGtoBgWfazVznObJ4QEz2vsWEl0VehbW5/x
lt0Vxgia4VCB13UFla+GJaGdxO+Z7/B1z2dCf43hr6o547P4NwTaZuLKa7ffXVZmonFMl1xEvuyD
NaEftfK7OXc4Zw4R/SPcP4djDFicrjkUYs504VnxwEpjvGWyuKwCoPGQ7Yoggl/0NeLNb7FP7tLd
8JKPgBec5nAfyst11gq0e3ytL9uZn4n0Cgv0dax6sMrnQVnMiJmOcOTkIEp4xGz11ZvQbKwcX/sB
OjBQJh6dwMvVrqoHAaE0wAr5Vmmea7J/wZ4EhBnmVU4MEnyFtbkk1PRbgMfe2piTm03qETc5X93O
GmrVn51ijMrLSDx3KTXOME5/NP1k0g1D/KZVQxF+PM7j7zkbOi02giAi2Ab6qqp9TlJ5zuhloB3T
tmwZodakfomvuhxtS/hddu6LwkzpLZpajFedmtQe4VbXA+sk1Mfg4KO66SdTiMV9sLwEtqk27pQR
h5bhV4KWpxg+J0ghwI6MQZC3lS3L92VbKBrE9aX24hsS9bahYHhemiyTpoLhgWRQUvTeRl1HLSUq
CZ+wUIxLYX6i1iK50VJoemlcShudR75RoB0ZOR22a/NbNQK0Bby8vqXNVHUtaXgahK0tYm6zhXXB
Xs3xGdVmuBEP9OqZ+niryBzMRKm4DzsT0euAAVq4Zdl1kApCEiTRfCMHT27f10kK4S9Teciz4lA1
9cmgtzgsKGNiERRKCwWVytuLkSqxks/kta6k+Rd5YKUfku/m3GD08SNfF5fqtxsiiDtKkNedCcZK
Tt7Gk0oaTqJ0M3LMbsuV8lS0N8TaZBzp1xTdVKijQfVqQCm8HuhBjsc1HjedK8qGsbZSI0htFAMP
5pzPN73hySEvULZNZxmvU2lONbj9cT+WAMhuPnjlTuuobr/xtRY2YSMzHXuAoXS4102GA+h7HNLD
pRwsrshVQT+6aenLu3hZ57NKTKtiy6iEHuo6YuWEuq7mnP3b+eW9ZTuJXVtuFPU8VLSwQDOd4poE
o9szBj59CN12XLCJJDhzjzj1vMuWQ4ytrdg6wTBcHwipUR9XELytLN79qmNik7VwdouxNNre9k+k
+2Rf6hOzBt2uwlAIfgaTPRX5oYt9mBvjXp0o2Zy9QxbvOq24zCilNzRSlBy0cfrIzEcebuR1XO9e
H5lri3VcEPhGX85lzWdA8AjSuI/xWtclXrMvP1m0B1Y7psbcJc6DwAazjiF6pPsu//OG55p1nJwR
hr4it82xjq5JRwxceyyBxeVvV7V2WwnBInv++udBUN8qgrKeG7Bo7cFcRqr0ae3f/ldJuw9qfmlu
MeSl/8OVx0fBLcnbV3l5HkcsKy/i9KvPszr2PKPWm8vdSNKTalsTtwF+8FfR640smbQ24L56Eb1a
+1GVTNOChr+PE4XZVRPEkz4OIpoZUnlWSOrStcJ5zIS87VOFqvjG8oAdUl7xm8q52OYNI7gHl8+m
4YSkFt2z/y2DaILOw1SwtF/MnHvlFxBVsB8iEMokUmt5LgNKt1J8gTfLMJbbIjqCQguubHhpP1K3
yCF5uvlPnTRsYCX9PDRRR5VMusrfzmdcqXr5aVcFzyUsb8dJN30biDs/l808mnhi0L779oyFuByZ
UBa99y1dBGTdzdObD/+n6gA1WGNpWiKiYftSRQRbHEWWlR35DLgWs35JkE+fZkDq0FOSBqY+njxz
gMbWeBHud1q9LtO0E2gT76y6VA94JNDG/T2kkrE7vG21hyy4wgTPf7TiZ2mQU2kU5yeklPe4liQJ
bpNyObhid6iQzoDB8LD0gLBu9+7JATC+xvRAP6aT1SSz+rry8rrNgbyMaSfZQCrcUupb/s7kkyO+
hrmAMkaDHzosTJgkZua4MBIGZnDyWpkRiAEs5fil9XxAEy0x+OoEYJfc4d1pwB3jfAxkqiDG5yA/
k+JnYUWLLjyFyea1Yc2kv03evhSU6/rCZA9CxzjoE1FoktDEjNDabXj7VM1n8ganh5HFiq4Q67Zl
ACk8Sn6BLQDb+L3qWRPnkiV1Nkl4SB7t+1otlymG7bt69i6Trj92jXVIqww0DrOeyp8YUJ5hhoB6
116+Rxi/JjIoWNQEp/9TLDSx9LcH1jWczOwQ/qYSVbkAOJzPCp/4wOTLK4VKG1R9JAMx8mHEZWdo
7xfyGG+CO9KH6L3jEtz/tYj5GXvMuBuu1ZRZN26osX7+al9eIo2oafYShx6ntg5M3TCk8DFzGdRf
oHvOSnQRZoprbTLc/8erYSDiA8PBJFkPalgp1N5+7NP3dYNLyR99Q2orG516R0Srf4UYZLvnJtce
Yr0OS4QuOS5NIIi8biUYs1xzoaPl+R13agFNpEXfQ0j5a0lsfpUQCBaFaz5a4cnV+R3hs1/xzgWJ
n/j0c6fGZuC0/a4P0MR4k0LrVSaf3r+0Qeg9NWhPk2D8UE89tlv/sOzn2V8ABBQmynhTznpxAp6q
LDhfOjJTGrxFVMyuWWnQYkabqbYaCIkYUSkuZd2zzTKEiA04dXvLSwJcqh3Trnu494dU9SmySGv6
jN8hDmfkFSjTuw9AhUBmtYy0ekKullKruPItZyp/drPteDqv8Yk2VwwzgVHq1O3m2noI/AQM1L0k
OtBUPIa0wcS3rkdG1h0OnTJFhAs63CYdYeZRycYmKax/UCDF3RcuGGPJQie2oNH9+up85WFXAuu5
2LEh/439UFb/MjC6zWE9DE1KaYuAvwTe5YiKUxIk5uoj9UTJ/M+U66GgZlcg+GnISwHdV3w3xic9
UyJ3bCwRJorivPjMBUwDlaFOgtH/b+wy/ZVK6Un8zLUknFcKUGaJkNi5l2HEAuUqGfEVgGAmJfer
JkudhqIj7+n8gDpTF9GCEPAKLpJGI0nDoe1G71gzxu8ftSEz5Favo2lLguHReWxClrPjfDMj1jv4
MUP1Sg4q/BVEYmLZ10IJgf9/YRWTDI7cvLVIKUJaXVz0Wi+WFOSUwl68v+GnnKcB937ztkx2uGe4
06Ex1N5kk4AQiH/eDE0jrk1zbMKpB530447v8Gg0/enISPtoRznkuCcRR9M4vkyUaFam9IKCz/72
RF08XypMQ4UH9jdJq9TqRgvUOfrpidtvEmu+T6mhYijqyl3iXqL/5vfp/ZdgrFTk3RUSNcmQKjpH
V+Si5/MxlamMO1ywtcVqWAAsLkWmuy3btgVpBPnzH74OTtKr+nhZVoOmgoXoQFpGtDbDEKSJMh4m
osmMzsl+d9taoi6Klmum+QjbT8gq43lrgAxmeE3dZ5pqn5eueyCTGAnSHj6M5AVhIbYqM3H7zMdT
3yGkd25apGd9LiMSopjfpM4f5Wj8ioa6Uqt+VGwrzfKwlZq9xkpoWp0HsZya0cLxahrd7Q6eEp18
FxWjLzmZl++zNRZFnBiEoMSzvAzsxhiy8lDWytBhWW9GW5nXg7E51YaTc+f7kLgJtuu8BoJpj3Rs
Y69am47ci5qtJE/OLvL7ypsPXttcF6N4Zj6TllbyiMrUndaS0Aud1TRxs4H2oUQjVaWPKyXESeob
Cf/pqeHMBqxxEZKXNhnU3N7grR1RhaCKSntj5tsW1Vn0ZJi837Gn4L19cKPYUFKT8oVdE6DirJLH
E1xTeGcrQSdQ6ezyEfh1j/Qk483o8RO7hpwKAVIQKrZfEVY1d/0aF/aizWuT8HuYEicNWIdFIRfU
Q6s7DugGvKIWiYVJVrmNyAeaXuKa9O9Qj/YJi9utWfNQ9ovGPrlUkJeccujf1dTWDjLdNSjj192H
1Bl5YUEESI6eKaiyF5yDSbM9JEiCRTYRUbi2zENMS9eUr/+S7Xs9hO7uPnAiI9smrqQG4fLcWllh
bfsXgwcB/wEQrJX7COo/MI+83aduKCvgTghvop+GPu4rfw+RNPXIpSWd1duxWhKqU0Jfb8Bq5nxr
TpbK+Lfzp0tHA9N37iTqcL6ihf+0e8kD/CKF/ToVWb+Pd9VPrSvjKBXD8YuTlDnAJ4ulBbRh+dQG
re/NKCtjWYLRHlXlQ1OHV1MGFNPL1e4vD7NWU7FB0NS4QfEwBwlG2C6/cAi/6mjCvaTTx7MgOgDb
BW6WwRnHwAMKa8TGMZSAlF0ls1G2oZC+z1MC17ZFnUP98Vt8Z82nDpOVbBEjeaHB7RDbnMdTHwCU
FW4lmAmD3L0hyqLqfgiTSoIFSVZzkfb7QHuQR+Twlda2iLqsTkCBp3R/BzhIMvKQ9UHY4hApxByf
ZfUC0VjSAnMVTs00A1eMzns13aPgHumaPu8CD4R242jcl6DryejR6VaNN27+EKEVx0qoz/ymiCtw
1/gExnlwwP1Eyuj/feUXbTy9zZXQeCnxswbSk3AMt7vDMt/9Y//gSudblGlmpUQHRMdYfZpF+R6w
ZWvI7JJx2pvqzggqIap9rNNzIsVi/hnJKZ0hJGdBQV0lEYzH2f27x+cWRZsrmhq+ST0EAxAd9nnS
lipJZyd5UDKmN++5FxmDZpXUvHyQzr6BrNhimWAwClwQsLaW5eEzBqkpvHyAbbr0D5Kx38ArI0c4
ulxtyVHtBeicGMAq4zXuSVl8XAj1LHGyMyi3SZk5dUqM687TqMLTUFna80GuGGRbxRDIZB9+bxEr
pwRqB7CrgMuS2LuCxkWntSFNjgLHC/mg28zVWxpB0+pi59JbhfIRWbw/DpbXdk979tG6ONQbaK88
G4qaFREflk1mpm5jG3qBOUFiERFMmf3pHKhwAkhiCZCzTO8cYLJQ196meJcajoXggkBW7ONfn8bF
F5kDJLeNIDNRWoHZ9Uz5f+aG+/09IrbOHByp4W8EPk2g+0rap/QMNT/oPcUhd1IsREc8TPixjKQV
nIk+sh0nb4gqhk4x5XO/pIU0a+0R4upUwSFfPasKumaiMBCxh3U3/feX4qajpo+eVOjqWKe26WX1
mcH2Tt/yIPs1CWi/Lk4lPGO2GLC6lHKU/HT5+TIgDcZVSPJqeauZcXrxeMaaaF4lyJ/d5e+l2IvE
WG7HYRIkQfKGm0BmDGWULPMz6nYYIo0e2vT/ZbShFlhplAcvpb1gxPKBfg1O2X5nzPDpZ7YPPBJu
r8qhy0kwgRpmQ01buX6Uymbpt0phKY+pjyxvBWRQ4wQrSma7ozIP8iEbvkxU6Vy+j7qxa2ALYjPp
9fC/EbCXqli2D1B5Kxwb3YkLSG1LlLh9OQ1vCOT4Q6HTjJlqW05aCGGeGFG3pViJQ884R4FYcjrd
EQ+TejNwA58jQsZpwgxM1ofzkyNFU29pClm9tNh+lHzbKbSLMO8CedcHeZ4i3//RLJqNqzoq8Jpw
cEeX6Wnrt4LlvHDqTSCXvOXUJ3NUq+d8U39uvk464rcJ7UFwWiLg/6IiPTqb9wuxtqw4PrItu11y
U2Su4kQR8JDPRAh2S9ze72vPqEQvSPEWAOtHwJuvjbPa7diFw9P3QwwjWu2RGrBr6Vyq9mJMgEwr
CkdQAMoY12vA9suJVlfG4FyQPsZPHhWGDqJuBoPBUtpScFshEzS5wEQF1Go2fmituPl1gs1g2tHu
a9ci71Yidb9qNAekMfwuWtNAB+V4IF1QXGxgR63DYV20m2Ii0ZZUXS5k+m6yG4X5T9p/zokqgE3T
oiEbngMDbZ3tzeJnOxW5dcFh0K5e5+eI1oXB60ppEghNkfUaiiD9luDR87DP+zhdnviB8ozdxf5Q
yhEc4v5QuNgy/26T2XRPH/huJN0qfF5O6YZBJAwUWEjeWvKKYj8Oms57yTexMCT3wL8tdlA/9H41
5CU65lzkf9um3Y17ntheShod8OOesD6EmOSg3a8ufxbJjwGZ/Przrrd0d5y7DHQVubB7/A07atWr
e1ETV+AHHANnsxPxcRo/WiEfLyWXc97P/XdXNPGWmevDp3/x5R7gMtZaeEhY+1Gd6IxrgW3ZPoNS
r0OqncwnyM7uckiHbQal94kH8sn1C0mcc9E4ByooDHk4ljUbGxASsm1telaGLUkDF1M1StaXUQ0J
GzmEAFLFpyHz03DE1Xq9BbdoQsEaUvgEKeZUYAeCgf0AzrVXeW9RXr/O9NPGn9fPtlp/t5YxJmn8
mCy9aNQyp6FjbpA4vTrH+/52gCvRlePgwn1yFrATOu443hlVpdvHoQShUXySF8TkFgL8+QpzAEBo
n4m78scJNVQ9a4hPoiZpoktYYNQrINv0qy4807NfXmnJ5/H8j4oIwBpcd/FwtbySAwAV7FrskFJx
MNm+pk13RCIPFpoX20wqAfJ9od3WYVVvvZ+NLTR7r5yxh48uZYS+2wCeHCcrvMmuL/pAZtkNkB2u
Hk+sghsof7SFnJIWXCbcYRR9ITbDvl7YpDXyesHUIaNumXtxJOhqcYqCZPfzSveMwpOY0/ll1IMT
zjInDMIESrl/fioNWuxjUAaUD44/ArGXwGQt0yeEXSDZnzb+L8/Uz/JmKvOkzyS68x9nYhXWNjL+
G8UnxNTKHRPuY3JxgD2Fys86QLoibzRADUjFkNF0Fmz5QiHbaWasFJUjve+98DmHV+fl1B24e31H
w+PX1A+SaeLzzKOPUCGxdSB7p/8+9eZuJRIBD8uMXT0AwKYwtwh68Kj+TA9A0pTfKO0rZzrkJLJw
hJwTZNssCbdHIYs9bvst3qiYEATAbdAs+hdnUm+OFy3gSxVjfp1e6EWi1japjH838ql2NzI2LL3Y
rIGb/GTJKKruUkg2VxPEx+NCuSWEqcUThKrYP9q+k8RH6vfuSYSd0vSNY5CdbRLlD5WBVlZvM6K6
NPEdF9nZ2XhuRx65ymML70xrFaIM36w4djtvok6F4mxMC6de2y7xZfLglU2K5xTblX8AccEllShZ
fSbv24Q6MDF77A0iSm7uBuhbs/EtFtEBObcZkdkUk07DZm3VbedVU93Qd6hIbCIbPCyrpagG2MJH
H3cONcnOBpUhuXyYfSf9vJLM98vPxhZZA8fplXjh+ri1KY9VIHydtfJWtwWhtclhibvU3HlBsc9r
eGswghcqPD7lN0M3pm/DWHsWY+oTVcD+5LP+m7o/ynrFC7xWPBvTWTtcZp0JMSUvzjf5zKG4WapP
m6K5KwWI5X8jU7BdLuOHAXgWWPMxfdSGTYc1l4YPMn+V6/sIavX2WWR4FGCrSxjA7DcbMK9RhG/D
QvGR1cZefI1vd08RP3JCZSv+pXogetVGu0kPrws9vqhJWVIRLqW+DrHd7zjszEa0p+fNi7D7laiI
6eYQz8a6kPWlFv+GlDTt3Y6GZ+ugGfVMZhH9ghXn05vR49dGzrBWrPJodGx4xEARtWYK8TW5VKQS
pi4TwSDB21ZcvOBhe6S2wnqROi0y87m/1a2Lma2zBlyOGKLrHBjG7B1b5DFXKmnW79ZEeMVS9ik9
8HtjKBxH1+EX9NUPzbdaL+2etKgaBVLJsuKtwF/VAHmuXpClZDE+6SxVDE2HwzyVbo8GqawGF+7z
9vSXGTqFfta51c9ZNLCObbPxwmegulalwjSGHikk4OSQ2QfIaS0DyNUH+XpWqRNDSV3kQw0mnr1P
OG7Szy4APLEW0sKS8GhfGBu5R7Mq7HVqRZip9duB1PLykYDv2Zv+wBfMexCoQ62BvC5bbZiUnJbX
dU1kRmObjHyQO8J/67jHORDBsTZfFsgZ1LvdposiYShcQcA0kNm6dg/Higp/eRqaahwnJ9FdCVW8
3LNok9XdFLVj6cv4/ile3yC+jS5uTDlqKILiYX3rtJ/ItBYJQsXsdYuYl6kxBHket8F6iGWggCFc
wn2u8MEIpjo0iQr2WWe90At29TpM0Q+mgVWUH/uyIk2ndMTT3g9JzWl3h9JvnkSAUFcbO+m9lx8Q
SEiPWcZzDPQQFMlIajoMcGZ7TPI1JQKEfc3mSGIysFqPaq618aeGJ0KG2bVeNCzg3VSDK0VlsS7i
K2dfYzpZztKllVxO4mpzTD5pxnvHQCo/kW7LDkyivHlHkjPTAnaEpH1jFUPL6l0Q+mHjrBkUjsaP
YM7Bf7PX/jFBewFbbD6kx7H2p1TryiWqfmJVASwZ22XZ6r2uq46DBaHW37yBcC6oY6C+ufq+BlOJ
R+Vneg01YXOfljxiF7PqWOWxUVGYbR/98quz4VdQzkYOSEx4MXCaDZKj+ZHVf9RwPmqdZYslTWP2
UKAdIlAa9QF7o3K/CAIdWp9NUVSofrZL4SJqc0dZgqC0Zbp8aB9mVObwx0DDQUbJM/4QHf1EjWPC
Y444XcMlWnmtl7zbySzi9qQOfnfHooMa7c2j3U4au5w30aFJtXS6nmh/KOXzu3XDEgT5LdkFKN4U
nQsBvS5MmE52LXsN/JVTtSyVTuJGnYc4ix6nTXI8cuNJEY+cvUkMAdHHllaNA3ENxne9tMn6cRPY
Qg3RoeYosPvxDatQPAulPJnEGZGlU0rA5CDqos5eJHap86uiijLIVDiNV0cPKn5/78aanvU+2MQx
o2mLYWExuRhoIpxNz3lois18hGZwHnI/w9QBRz8Xi1gha+43fR5Q91mI/BUt8Nh2fgypW6Vll7Pt
3uNdcg8TW7Px29maJdPmAnZap99ibMNJZzWcI3wQfNIQ30BMeV+hSAr59RgbAViECBds1pI9oplJ
a7k+7ZQMSHGWWDHmAGp8P0ZhMwqz4mCIw8rUrLacYdCbwp11u/6IXxCmKEs36xJ6TJg0/tXz0glc
Q0xla2ASRm7/xxJP/fhWOGyIa1Ce2VoEGD2DTj9EN5ojJ2c/51uK116Xa57xjXtXNqPKUU/2L//p
VhFV2UdSU/c34+fTH3GD7dxD7UyUNz36EsAZwjsh71N0f49mgNKph6IxdWW16RofZABfuFpHdF3g
QTVdUcCraaXhcr1TuITXrZxbhHffO5rgJVT4qXy31ZgROtwh/U/ysZIR9XuCe9OubFE1b9xKgjop
ETYcbfw6QN1Wk19RAESejA7ILhM9784JxWV3gFS8VwJY7a9W00g8mgfCvs6tPEdPjBSZ65qyuWIQ
VLRHy10cPK3O/5FFRUHPbeKIPW36QP+nSnlGh8p9wP+rQaJjmKwijFgQrFu3sJhFBU7B4m4ctKHQ
I5VO7SCm0X75gVZVboamL6Xt3rk7fmCqINEB9OLsHfQw17An8yXfHk5Yjrsd95tAY6uRCJ41NJ4S
hxxlR5L16N33DY41D+s7vfgi/HMwokf6bMciBVOFZIZ/LRAueAn2lpK6o2/vUBJCHmQlOHQyCMD+
QB59QbcUp7Rj62vuqlAL+VwaQ6Cw9eStdF1HyBBSEAUfxBtDEBPJburec2AzR5HK7uuZkyH10ksG
1UqosqQ6gFN8accMscAktRCjiGrooonEgvBQklHFCXBYu3Sg2GcCgKHlJlo1OdfVV0M6GapaLg5a
6qRLdqk7aYWev3SMnJK05GjwsE49fT+w90H8vBsf7+kDNbHGwDXsRuIZ07nLFR1hzAKtO8iOZ1zF
rA6uk9A6Cw3pHH+pAxqSIKZUMx4ezsaUujVEbo3ae9f7Wir+dcs3vCYWqj962F+0QZDfyCDa9B+Z
4SJc1I+rQOTyYTYKVFJlLaHxC2euP/hWyEkNwRspCXSEgVt9RgYC3Uh9KjKCCKRB44Cg+2f8QMxh
EbUbWtq9ngMzgB/ogY8ayR03qzzf+G4KjFNZJBscrRViacveV7ssHPNOw/uM5ctnfATSyKyz5SGe
uyIMLby9fJFrHT/S7ShY155AD8FtDHMPXPMLMh/yXyqjYfnCcJ+R0SzwDTMr+pBmpLJSwKokSb0P
2hBlPzPT5LEdQNTMAg5coczRElLDt4gaLneEkheJHxDM5TDjgy/lhlCz+9vWpyJHxGJROOx1eyQQ
UsJ/qfJA36FALGeUvCiSYSF68EzReWGRcbfcICcKt1QFTxVJQxAuAjRsMHkWPwuc3mM6RNvp9nPu
9VLP4VH+X4ZMYuDwTHemTLdPwHm/fcvY+DWlGPmFSB59hJ7Mt9MDRAiB8DqMztM5UzsdtIVahooq
R1Y4jXRTpYMemf+MJVB11u9ql15Ar0wwg57dps9wtcbjXW9RhZOKbLsienA//VSsvf3cfwnUyGe6
1lsdwzBdyz0dHCFBgNSoiftiqLx7lQYMhJ0U5hB6P2m8JylrT9pbGbErMWZ8U1SY89r5/JuSq7LG
s6CpvGlmWWa/SnZk/+eSSiGlj9WhMzHS0ZQY7XdvFDUKW5kOA6yGESXjnkp1DxGY7fGb2V/wg5hg
tQaSmftbXWiDHxC8NOcqYxIMaJGWx4eYrZD+iTwpre9+qvyPuBDpITlcCJeRp2PT3yCxIJB+ffis
OUuwzXHf8ozY5AXZ6GF3mWOit4aWfNFcDskIp1q64eQitnorcjDy1uMrTL8tB4aHfSJ6Ny4Ny5Cc
x6VUMr6Q0WAzRfWdj9E8FMo7leWGAMxoAWzjp12Vn0uoTensEsmcJ0CCI2zlpXzBwYafKRb5nd0/
hdyL72dRXLIc2mucaKFQrqAl3f/IniunHgZcVIjO6gDuDE0+SKDhVvNlLOR1jKlod3gprxqqoPOw
DIjcJf4c/pZsvWxOsPT9aA1bexXPT5FH1YJH5U57pkOne9ISX3CfWHlJCEOsGMMKFsjsV6ci+pm5
3ttqdJfIx7AcKSd44t3KIWYDzBjgc8V/SLsapNnKngp0jHAjQ23HthVJW1hKNkV2yRT7GBfg5W2d
w3xVNau6WCrkS76uOVSphEceuvXkWaXnf+CE0SfdfIzej/JTbMJlGf+ptL1FP+aTv7vGtTQyj/a2
S2Sr3/+TZ+Jwt66CGNbqzyj/SvRx97kK6F+rfEfi7y+YnEvXF7RVxR2+F+UCuCxnFRmwysGat1dn
5hFM6bT5M8YjN7ERBmOkd27XJgyDWg+20wUP+Kh9XclLXTEMBtsDYaAdnj9AX5r0iyeHF4yTuWoT
VIeFcltjoLbfmvEVipwR09leSBXJKVZ1NT/dpcsHxxoojLsAcgEqL1G9UqkoUsV/1nS4AT5NR1rM
OXCEe4VEh/iZE+3owAeXZgMcvA7Dd8s2DGsHo/3McqepPqIVGLKzMWGDxxCICbbEhCOPyVV7m09Q
FvD/IyAAPjJd3fUb6gkRwgQRrwtYeHQfk9JURrK5TkKiqa2Kos/uKJiQen2pa+CyaI+Q3oH5Ia7m
X9o3xHmqt0z2tn7lV4CGup0dqAfbtlAzCPvlEnoiYA2gFs+5gVQyZu8/aJFVMDUJEzL5mdla2Jcy
TO5eUoKgHCeEAAqCLxBAggw7D9vizejL3tiTNvSvJwRz5+c3DYYSRxMvVdVbyuFTc1WO+Fmj3rh/
z66EchzcJ06dWemhNNAshirMx2vSQkMa4h6yX6voAoi31iy4e5/Kz30hZ8C28dyYjFHZYDUwPtey
65WUqjN8Qk2ldwJKNyKpP4aRW2Xx8tBzkLmHtcHa8lLhpAC+96i/w8it8enOvgubaEIsIo7kfu3a
n9RGvUQVBgKgEHdpPDfCyXqZ4Or/3EhjFvwIo+KvWo/wF8/8jy7d4asBxjc/rninitI+fyCcJ1dL
rKI9FGxp2Fp2xYFTOu4Q5yofpoJd/oQ7DhGCh5+/0HVrlvG0B3KyXpqEbELu8FkXHvNaK9EOgeF1
uiMTqBBlPlzRrpVTsJgjy4fdm3vhjDT+GmAo5nBvI0NaEg9w99Xu52n2L1XoWn8FJpyfD9uBXGXh
00eXBL5I0B2cXomgmKIRguefnHEqYVvW9lgqIiu6Sn8JKgq1qP0NYhnfF+bCnaPxHXk4OovnTRw4
t9l8HS8hQQOckFdQk4ItU9DZnywPJqK1uO3yjpLVvsMBRnT+9+0wLb37HuPFTfz/Y0U6LP43GSPZ
a4UwDr1opR6VN0c8H+D7rwbsd+eJHps8V0Uc9qLWhQmSKyCe0PYc2Mwa3BX+x4Uhz+TxhA4BGA1n
uETKVE7gitcES8hOxM3DYzg/Za2bzGo052Q4B/fciVN3xjFQ4XceG9S5UoNqfoAOcOZGyD4PJJ45
PgFa6he2cGjNgmOk1aW9a0C+0omia7u41u+g/NVwwDWSuuuVfrWcjDyL25SYpg3vXYtc9ohGsMDY
2dFbT5FU5ncd9EKgidYn0k43rvGvPNbzaDALQ9Duo84xTYpTo+WgZVZYWllKfLYjhiewjYclqaPT
hYWjBESbmDJKpFb/8kosJShtx0YvfHphuIo6f0pJAHryRogMdd8RfJUAqwmREuB2UCkrbXpOTfTt
LIg/49ZiKvPRZg/JfqYlsggIXmGcRdfR4G0TwhNzvujhANvGPhtlHA0dK+kBHfBopNdCwHKseAON
I+UJpAJuaH8rpkTsKyC2gzIICBB+zTQB+BddnRwauKXNWLbY3CACPz7Tvpujc+MgEs3E7+9r2rHp
Q2hjuq6Zopyrhnso7lSvIi5R2SOqFTwpsfVarINq9DwnBgbB49MGaECld3UEB62NGKaF1UwMLE8Z
uMAhjyUDElWBgC+FL9xk87Xl/NtBBCJG5BlgQLQDWlQm3MEvvZ0K29crbiqVF++N9TjGbNnR9vgZ
oLzgM8BainuDbDPFN7ju16ejFO4xh44guvn5bJnPMiSJsSLD2wdWnG+Pg+8yOLi+SCxDiqLzSJMW
0tQ5XKP6+fqGivWjedT76EzjM+VLmubU8ixPTaNGUujdTS5qAVxVSqAyHm3+6Y6aFeA5GK+Rf+BO
EOVVCMbgiaKs69atFLhM63iAtij+Jezo5qU6NHBPF8abuI6bEKdpw7+9bVj/OssYAQW0LXpaKHj6
HB4QWG5IuU9aQdJFbCQn3SZuDjyNNtnBrFKD+0xVyel84dmB0mOC5TS0jz7zrp570jzU1p3crLjq
STEV3v4sTg5Ks3h6XIORkFkKvZzpZx0Pi1e7GspU38bWSAUAmIRToqV41Pr1UhU64ABbWJV4b/U0
R3ottidqygkO7EENypWdZm1sy0GDFc1c6CtNOMnZvPfkRdsNHC3r/e2PavHs/bY/zKiPlzoNIAWe
U2EQ/fyAgAOfoHwbAh/L1Y7kqJEuCIizCXLvjCcA9x0pvqd1khJuSqJMNuOmNw5msLOavu2zrr71
U6Koi6PVsJa4gUh54YQvemz/QxYVW4hZkXArlmz5TE9VKNOS0AdJNSt28FpnhX5F2zQAoq/Bswx6
U/CR/cpnz+OhXJUAn7f85nNxlKeHA2c6YKHEJD80mtoNO2zriDf1tqqasFDTZzQHrUxy0INopqmQ
/Ll7M9c//wYa1iNe6+EOBLAJwSTS9CJ4KJbAHQDl6HZPGm/jUeeYEcdrh8aSojGujJb+66ri+dI+
5LU++bexd4AhUCP54Ruz9EjMnXlHWgqCJZMxNmNcjUuIX4PE6vMIN3dLPCuUqH0NIfulf8Tg50hS
XD1gaALOaDZJIA97b91igJxtWCVsXa6rzv0BexpUwhM8QwnX4NuRw1UwwKT5cV5pIEHGMlR2iWcS
kn/yNsz7KOqexgYIdZ6qwlCpsaPo75zR+dmn6/tbJmTbVgszW7zbCDcwwBQrp77Hw4+MF1iUCyB9
/Ei9sBgF6khSt+PhErSnsu91cJQ1zftB7v2HnDBVUnuKjHlZCW0QGCVHH7b04Vbz7dh/x+n5G4/4
BM5W2QAx1kLz6DBB2iV9ob/LN+9Qj+DinQjyjeyhTLZ683OY48NifSpWmJN/w2lPK9mO0fFZCzhy
VCqE8n0PdQSMZTc2Kq4g8NW+i1wevKBD7hkzpODpzp44Dm0y2H8QV+aJ2+LioOS8Zx3mahNnW05w
hNUiT+SrpSHkyAd4mTDdhiSdt5uNXYqtBD6n6cTJiAGk+58XBw+QYLK+tJWfwyDt35O9Im5T0lZw
mQ2hj0B8i2E9bH3oeU4ggOwRr9lJejbfOostiY8TM7TRGqYNkZIziiqSWOa2xlxoZJ5T6y7ZDhwP
WHy8wAa5WuscV97TFVDTDplM7sDE2yVsFNO1HVs9rrS+Otr6ETQxjwVLk8sSCZAEaua+22WKsWIF
+/uZF7IFAej6j4p5IkfqsXCBrzzur7ar+0U0mkH7I9hJhes40UYNcqtyWceHgpJIGjRsGWNF+171
4v5ugFbMZH7a2ooJjm2xN16mFxUAxwdMVlBS5aXSuI+slh346eMsXxDZgRvcX9wDD9tRkMsqjBtE
QiSaw/4dJ0BhP8Fre+Iu4flRpLmMJot5hi19Eegceq9GqBscVHZa0pFnnIZv1hSKkAIQZokkPRco
DbubfNNJTv/rK9T1pvr+lMdh92h3eFk1SNh31X4JRvf6KkBagEDyFEM0EhCP0p3ePYZILzaQ0kBd
o2ADWhLz/Tq9sNpznEuYZAeiHo2wyASdPfNeMOweFoDqujk4bbMTF7BoJCfj58b4Kp2Z3GbQWm60
WGBC718lxpJS+hleaVwYqE0RXTXjNPiuiF4IwyuursZx0yodsbw0RyOcBhNtGV+lPRl18zAfgBir
jugVgn2hRiQTs/k0AeFw6hEdtuDddByQMdYiwj+QxhmBx/Co0B5Hl/9MPNWjNxBEIYsXvgeTFwpB
qADRr1Gy6O/v4oMivPU/XufK/4AXy6gdFp3uXo/UZusxTRf3B3JLlwtUSExNRY02R6wrFqzWv1kS
r2LvNhxYRJoQEbhXagzWguhW1j6h/+R4mWY8nRwkb3YoFqjf4FTjB68NsEgd+Dnkcfa28542ckKh
8yNe4iuga7eScS6jDaL0KZs43SmT2dl+7sEWC9BDPk25qhuWoOgNe80OZ3CsL94Csjpi9TDBv6Q3
URtQe8yj7TbDqYZTm587TdU9u0ZH71FWnR6tUsxgxY/f2+Lc2zg/PzwSP7D+eMRelFex0rJs2LqH
fHP8qTTEAYX/i49TkP5CR64zSjN16xocHTRWa5a6yKn+Kfd0beqMKRBhMAB/+TeQPscoG3AxcG71
bCcWDFPGB5Zh/6cyPXrtKZner17y1M7jQ21MbH5g8Xzhz7DTYV71lVRLhCn2fOKI0Wm8jgc5zbMV
lq+MA/oj1WflFYShthvL3gxS8XrDjV08wr7EofIfw4JccjHkQHnRfPOyCd/cacsFjEZfJQ0yIolq
hHNRnZka/pYk2Uuf18vyEOyIUh8kwFPsLucWzy8XzhlFgMjY9m9xemtBfW6U9O9qblkKgWT8f1Pm
Gf9Wxevpdk4lihxupmWP+RuYI3+hcl3KfVgKsztqsQMASTP4yHl1d4gS8Uq7S62AgeyCuoIzYWyf
JODwbG2RkRhFvBxVMsvk2v/uynolvhQe1xMB3SkT1iALdKoL2zkxjbxZti7shQWHO2PUxFhDopKN
jIsYFnAV+7qbBAJ/FZ1nXrbUM9ohM7OB9+GDfUWK4t5gwq9iorzzPP2GaqzpLinVoLV4L2uXISKQ
7T6yVudL8qtLVjlIvCpN0GFlOo898aJHLY/CLlItZD9AvBjwBB+q3kfgVDW2q9M02P+ql7nUsD7L
Ccm07EITWl7y3pt07onkfpJbF1Gvf7qQDmqA6gfoRINCjcciTKby4WrE1ixbYTblhG7qI6vLWrBq
Y/vgN+lZf82vDOC/3etOn3+J3OHPIG9wyaBy5oDiYEyShXl/mjL5gbGWzrde6Tb85lSsVpIx4KLv
Ob8JddaY2bi/mB8KuuP0fqNcxkBXifA70dXmQoEwvrUSeQO15K/GfrVb2Or9WXoiLJj0FVFGuz15
To0ep5CCYRep6EHmh0FM59NJc3lpqNbvnZguG6T5vFFfVYAfKwP/gH57jCH6Hb8cnTW8Z0r7fh8j
1IO+CVypkxM7SU/jHGv+peiT0Y3eOlw26Xzc1CQdQAs94e+IBHqqazQnkn2+C6FB94g02jtlrzTK
gnLwwBJ1DuIv9TBumyIv2hr7TgtfwmiYTmHOQKmtqreUGCwZNIgBNHMqsolmzkc7hmTajxB9T5pw
xRzuTg0/Md1+7pNHTh0sSF1HjjPI79TvdROhjsAoUazKjRgx6pQdRg2sWq8273vo4Kou61ODpQ3/
z6gGINCW9jbj+KqawYbbyMfpD1dFR9ZPoWcC1lngJzWHAwmlW570jdiheYPIHhB+sEj+SL5jcRkF
azSty9tVe9Xy9k6Xe6xEn7UrfOIrlEa/AukaYhCLrF88g9KAL4uDN4VuhvBEqVpq53Iec3r3IrLo
AZq+vmIbBIgV4TyCWjFqYushmP77+HmRACYcKJL7Rzf9pIAWIO9UzNa0iMf/F7y2cb1kRMx9kJWI
HCiSTR7gLQzAg1IVsqqOdhVS3imhjf78nkTAKS4t/7BGSCrLCP8WalaW+e7+BioE/19XOSnkshKr
o2+ek7+QgwKW3uWmUX9+7v+pEAGorVpNaVYXXduw3fERHUMDfWtgyOWQSTToBDi9aAccEuVz3QeE
spG+4Db+hKjPEX8vK85yEG/uCco5sn4d3sLgNzEhIT5xciXMe2yiGj0gmP5t69dsKFqYMhrRjLl9
NjOIXFGoYppkNtmZHBMtkBTr8jIzqhI//EMBPbvO0SyJWmVZZvX9op8684qr+XE38alR5IXM9dET
zDmVNeyOWev5S+0tENwnsLtOENZqv7nvWyh1b3G6M38GBk2vW3QTziyzUOaFsnsUy0f7vMgtazrU
MTqD5Ps2p7ySMUsmZwgoKaaPGO6WmJrZ/w3p+LGIMHC+RwCSvRATNyS4Uj4BtkrEiCe6pGxvE0aD
kair2/CGH0uajM02J9Ntu5GDsIcOGf9U3EwOXewQ14NXl73DjfzvuA1zUF0QBrndUDedRflhGEFk
DHMTB4LXKplGIHcO1UcsPH096uXabigorqjnOycmIjp10E20Sw+7cHD0thGVxKVOrsuvdDn5A8jC
TN8k1o4bnCOecvlNJevtUafG0m4z/BSb+bSnmadYHbpfCZXNZqrIKoX7voI+WL/EmMFQ7m4E19xT
ESs+SfXdt4qw3P/DtUH/XIzuqoH/q2Pu77auZN4XDwcD9T2v88MrbnFICA+zo4ikeOPaWWZHQHeU
SgL8CwfdlCw4Vp1MHc8DyOmJDacpOThxNKuP+/YCQmTj032eTPBo/bv7msqkt6Py2MuuMMNrP8MS
gSGwVg0WhUqIrWwS/wa8BeH10hL2f43vGcV4WRBL/6VnwJVGVeTPzbdQmuGgf2t1B9K3RiIfCD5a
wHjm86VUr1h610KmdjxR87211y5sWj8NBQzH1UVYFGP6YJUuV2cfWYsT+pgtbQ5gduq88PB3JVuN
y4ED1t3vcLzXpDUDaQ4W4tcE25Mt7sjxvtgQnC4tQjn/SXOlIXiNGbQjd0Sy1prExFwZLemjzWNT
4R9cwEnmUvUjWRevR5ROzJMw0Zl7xAELA9Z7U1G/+XuRggnh5/qc9SZZ1OG5axEEIot58btB2jnE
iyjGD1YwZ9Dfw5dJjUTR5wsehZ9yTUQ+jfR4nlMPaHjwJKq8OupyhUpGhrljwypXIRR7VN+04HPi
PXtMLv0LskAExJoCSgjtZR+zlJpSw2kty5sqrnANJU0cmZWK/ATAI7bM+6Zu17OF1kgTiq+lh1Xp
fmrxuTyfy0dXpO829xPYLN7eLsLJxWXc4TiP24k/3hyN1MzxLMxmu15v58q/UOpa3uhQSdcszxx9
+67nse3an0MoaJK4k8SAZcmHERT0EVmVhaTdLjVs/SdHfhX+fEfBk4AlZkJ2i0JZ/UmuEx7/uhZ/
Hvdqo4a2XUxuTPky33toec0Om9anHMkByQyFwAXOM4sE1FAq8+BWcJNPmtU2hH+YCfNaOxrhfXNJ
gizcOXye+EiZLxXHspVlf9ueiZcZxjA+ob7VBAvP0iAsqxY+1bJFZv4HeEzsWLp4br7nY8uXoboo
bYilZCo3sjgpxscRQQzRqRscVynks1oApxYHcUgrRyaYAP9iaIz/uA848YKdOYi+oQVwxLr/oMWL
/au52C6inApg/8qR5djqNGmL7nlBToWZp+8Vz0U8QcnBrpzFyaDcDHdQoG4HUWgXe4w1ODFH5Po/
ymFX3sUWdGi6AbMFyXSLty/6uhGimnalUyv8K7s6n/uuqZlQdjpXSHaGDxP0oBg2A80cDDEvaMMM
Tk5fQynvYVVeMOY+pid/Qs+Q9acB2uXrd62z234bfXoyV2FeKi9JGRCfpd15f6+gXjp86myxuic2
o09nzx57YO5Pm3mEdbiUbc/u+Iceb2Yd0D3NE1VplgbIgUG2HwhK8mwz33aazFGJHbna0anfJDtD
VUDIWZHe3/jeucn5URnxRLGMG0YLu9Akp0bV6MjQKYF2OeGZGiJT/jH8kSSLMKG1ZlkxcyHtpu1c
KnuDFvvsbRFR8L4/cqc7+Y/Ghlica7XqsodNaS1nWFY96pqIAxXZkRQ0EySk4pWWBrCT/iRzEOBb
2DhMbGATDWsnfW9BTI9H79kF+CPXcJJqFPFTzZKp+HWPt2lB+zcUCV5Zl5MmOKd7Ss+uEKMtg+Sj
+Q/OoChq0Qksx0rJBOxBgpNxWDZG6H9Y09b76WckjNPHNWHHsa9esrgriG6KOwAgnxl7Md6nO76q
NM/xITAv0BBWSU3ZxpVHjlci+PBp9hXEEL8SpTItw4isnKXPBJkHDepj2TvUeBhwz2CXYnfp9df6
cuYdlgLhEjHGT7CJ6jQSzGV+AhhzX7P7C4Av1Is3Aq4qW1u031ep+wb6tkiSXMd8mMMWiI31Yf4a
isl1ZQ0IBK28j/hHV0SGPeyUyl/DSKSHTekFq+/z2wsuEK+7fhF3AEStaCEWqCxfVf11KR0eq+V3
m0tHH2Yi4/whTt9kEwdnuPlayu1ZdQxGtdBta3a/tReSpcrpfSyLSpvYtzznbStEbSlIn6UJSmfD
igaSos3nvno1J1dbGciPCbcL0TjEhBnEJhEOeR7fdodgex/ZukUzDG+DQPeU0UGhcQuQFIApd1+0
V5/GNYdCy8CgQx2qw/nxMK/UYG/8kIhO5dzx+1SuGHHNegnAnaf+7rKWmiCmw4qWz+/1Dd+rxDam
v1fcc4svCVPf6zSYQ4MYuIGzH4EY118SGk8gpC1aYvtR+MUWd5fYbmTSbt9fcX9J6f7UmajrSdKV
OjhovUxjtJT12njtGQWRtjZHcH0VXvuZdb4o7zUudW/Vtl0EeVDu+SjzTnyA0Ha3Oi3b1oOak5SQ
Hc0WG6yw1Rv6D5/VFSR9Pn0yjrH+Y7XX1qnrYKdwdha7ILH9QPRhECEQWd4isOYE6zHb947Tanwv
ErbBfM1L0ELMUORto+D1FzwTvMaslWZ7p5eb5ft3XyzsdT3KB11XudcBp5qKgoD9RGdyC+NpKtSI
1LdS+GTUkVeNoWniVx+TotQTfQjwjXrESCK0bKccXDu2V89fVVTJ2eXGB1v7D8N1fkuPMV0lG4Nn
OxcjdHVxO7Xuu/gIIzFASaM4DBG3D6wJI5+YEtwMfzvpn101OejtXkG6DVtSlYIY2Q9qiy6bBpxR
siO5wjM1kgO4Yd0FJrjzQze3c7aphNcp20SdB8QxWUo1QvPqAjHrkqaz7llj0y4CVjg6sL2ZDv5V
AOzA07mTItSn18QbKvIrzUO2ApVav7+KWEQXepm8ojKoCUY68wG/Ito2YCByKVpLmAkwtYKecZwg
S7z4fmmXN74pRnDmjtNRDiGFaYopXf10BdW+8hauNQTcdDDpwShlkWy7J01bS0TTd+No2xmU8lwc
SsbtL6rrVAQN5gi/7KK+B7S18B9OAZbplwG9j71DVbBrXlmokkFU7N3cB2XDRyGTV6DXQ55A0yaR
0cvVcwLXtU5jHC08jg8oBjOsVtHvoTEzAnRSOLPPGyVMYiDsdO9TJDprGhzRNnlC9wmmeq5X32OA
AgWg7mywgUmDeE0w5qwgyj8n7sW+H5ok0C0kVqBfAI5+cGtoDMFzfMsfr/a1oLLpZokLJK0acgU5
aj1v5V7/BsJbFIqY65GPGb3Rbn+WyH1KgA/MV3c1GhlBwej8VZO2LoLRX4hoOhyJWvWzaS1NguOR
IvTQ6uCzQYY0zrqL2LJnYPgaIvg1a2z396MJNXLX5F6XJbIzzCgm/oS/nPOsCGDhPf/Mbb02CWQ2
/G5dkjPMjZfEImUr8DsGOvbe8VC2UcOyb9ndTnCHFGRtmQf5B5xLCTkmjbvDV2pP4mf9DytKgr9r
w8qmpRP5sx5yKbOQVCbAiFQGKMsUnQeaqiM6HiOkbrt/1V96PSN+b3QFdlw8OcJuL5ztpHqeWIn2
tSz4z0Lk05FsPZJZYEtz4lmQrvoV1ipXwpsvzoMzUQ9dM0gpdAIOcYQkBVrstThJ1J4LtFM6A9sO
pQdelbeWoCFOms8szA0Fl1IJPoJO/6UiGB3TQ5lggRCcwqB4YFdiIBQNYZ3uYZDLT/XTWjW5/gvK
niH1bT5NJCeFX4W8q1vXeBuqoFdTLCVtUaDkrabIVimZLYcRtNQXuSQAJuKqHInO4XFeV5weY8FK
pamTwaFiFSY7AIsySoHwnCgwXYJQN3j8mlE7SsRCKr7n1DpI/X4B9El0MPfisEHw6VRJsGlS/2xB
lRiiXU/fzIzGSrvhTV2qtvKqMtQlo8tNC2UlXA93YU25JEdAaCSd4EgOZS+JsF8AYKZI/g99v3jM
6eM7xk8TFEynWqL8sKTB4vX3k8dIpf3m3aaHO0EiSFe417W//OBM9gjrkFtkHVtLoWcsCooeHXxT
mxLJOFsVUIn0/kteotX7KnGg1dysc3rWowpKYr67cXK1y5pq+x5wD2i5L7nJ2jzLPoOPGYBj312x
vT7iGloKET6iZbrJ2il0x0SbwWkea9ims15Vx1bu9irFgEncX9jOk7aiP7gPvSbVMO+6xJ9tj66o
An0/XjY/9NkuvbG8AsIHFgk+7J7Zdgg5NvbemBvwm+C3eM0wNi2jeMf2aGiWH1wUuHou9phbAkbO
SOULdzlN3cadtPNWJFOF+CyK32mYax61l5lLgVq51HYOo46cDtaeIFtueQ+DPRfgDsH/xdQd8xid
Yo3Pf/Au18Cms/OmWINLYZxUjnDOvwIOuDsBpYfu+vgs3GRzLaa+iT7NXq+e+U3wjyDCNodAPBk7
b5rwOB/+ihAff5ze6Hjyw2qi2FZwXwgxW9buv7ImbnuaFLDMt/xFLX6y0IeXenA4BrRC4z6B/G/p
K1jRka4rQyHMZDZAN/87QGZgLL3VcOFR0bbly7TOwQxz5dn0PzJ9ijxuKq6o/NTj+01Vi2WLqOv8
4we6cuDC7EzSY7WjrJfrVobFqClJw0Qln6KVrIKOZtBtuajMJhHrGSb5pRAstNXFIuW6Im0dWJWG
m8jsE0QALNXA3ZUtzj1kxcxEoqfU6qZJa6iHpigBcFVFquObkeA1kLC9J9mxpExVKNVNQhyoUVXr
bIz6gjwyiHsezVvER8Fui5tjCD+Dhle/ECCQwB/T9cmP0UtwcZUGPsbUYRIwe512eIYgBKSajgIi
KCu6Aeh73v0fW893JtukGG/BEQ6+w/MTJfDUiWiKUyacJmsEOyjTaJmo9Lerm7Fdj3gEBBvTxo7J
org2T600RI98lXpyn6x026zbJD2kP9lmQfaOGSYNtfd4JhF/9es0Xvr8MueRs9D/pkobvYxIAXes
v0Mby857hNzpXzgRYW5DqmYIFMCL60bkBlQEEhzLeBL1ll9ikW0uENqzbZHnYTbKp3pBN37lUcPF
GXlgKpN5wYPLfSywYNsmkUEoS2d+Bx7ZS1tf8Qo/Ia3FM9mzG8MNWfA4s35EXd7XK2Yyue9mAt56
WQ4n6DF9OItbTzErF2sY93MVVJytkAlBRa1Nhgouapd2+46rm/0cCUp8mXxuubx+S1AHuWO/vz/a
XQggtrIXwl/tdFmlxT6GvhN+bEMTZl165YkgvbpqE+TFt27Y7WH9xqQYh+c9l8l+n2/27/ckX4TW
aUamqqQts/623vfB3FkBhKAoRHa/hpxouFOTwQGuvdq9vwAycVz1E83aeUrKhSmivIalldCkru0x
KUJRMuPOGbSYnIxKk9ha7UcrWO4GCUjScE6Uv6BnjZ6xzr2i7VlIaGbWAH+iotsUL6IxOyY6ZhaR
q12xpJIbuuCC2UPH10YBsJhpo4UCA/vklzKYzdXYsSRUscAxuR7AlImljsTLVDdm4rT7b+6gfkL+
CWAUtoROhz65S9V7k6UoD7P51lq0F3iKMbvpfFJ0E9zyecc9R+avsXl9DYecWsHmwYGv63m0ORZG
sCfujjbF0+AwWeBNPbGx2c8cwT29J6Gpnh1/tawRvrzk8ZekxksSg6nowZaOgTU83qp0D5+xWgC7
toHgZDt0cqBqqoBRIYJgyO2t/6ZnpACGBKiVMm3fuXWZKdU85+OeKt33wj24ghPpwDAsp3PQpBKm
549ErGxMxYNEpB5Jo/vv33TFs3nzEa2M2ib6LspGbAqpVfvEwfujsH0UT9s18GZ/40AVy4L+ZXui
c2wnoZeGgPfJnXy188C/v1eHFEp8noTQbeLx7WVgwGeyYFeO9VloKldzgM8i4bAl1Jw02+IIU/uE
4ulYqsTKvqVQ4AjB0iVwRKncIj1igvv0Vxo+w6WVoyMmNgzVM7Gp0Wpzv5smxsHxH0pUUtb6axkJ
lcu4DeTE4tnPqIp/jyanJ2ho0tzqfGRGez3ilkzni3qSC0w+Vu2WuDIR/XMWDRZj9Ml3KbC61Wby
tsG+QLNp9noqNlbuwJarEJV80NPDzOt7SanGDnEyPg8QPXj+h6zvCOETLX5A8h/Z7csZXVpo1Zxg
HKz5UbWmSQqh/oDpsy9VkMGngE2+bNPI7XJ7sFTD4QRcoHkRC3nDLcKzb+/a47Ii9rNXWcKvXaed
v5VlfvxAcwSILXX06qhDG5aZbMXL0/PkIrg8TibJLlIgaZ/RpCd4lSA+3M8HYYT5NuKqSpbcM3v7
R5NDdzosoi9R6CrgsRvtPhNvOxxlIwKPy6GaVWu1PKoDF1sgTAG9b2+U0Ui5C/QaQ2th5uRwcEow
6XC0ZHpGaw6opYPB7EU7DN0CijXshnXUt8Jt128hJH5O7POpwlDah2KPgnDakIMS/LZvfEX3T5tK
uMYxfe/l/A7aP1H+OO+azTYiHpkKSnx7XdRqH3sBpQp3ShGW83UmYL55Z2XsMLOWeKJ1NdGNXL39
TgW+GNFTefxvpyjYK5vThln0jNHWdq85h5nayyTQnrD45Oer9Jzy3i6t/j5Pv9r1v84qQe7faH6Q
qSCBt02EAb6mPQe35cMkB0vS4iu9vJFZMNz1d1JVI9mtC8yinMF6yq8RIqOyC12tlLvREed14kNh
KuvSM3pyrVflVoRdJx/QNZMhvyMb0pSGtO4XkV4pL2tlQlK8v1MdE3jjt5LNGCZc8kI0gnXdNLl9
W4dn3vzOxCDYEgsrRUr6w82K9YluEIxidSmV0/eOK9T671pX8yaxvc6EMSkeiAccEVaMel6pVef5
TYxoapnooqiXVoDquS9V24eKoEiJiUsTXKHmcWc73h+pdIDZKP0FvVCK38ROGpXmXtxPVAy+djGr
qLLtVQW0BKws+RdLY0D5DvgH15AN+Jcwr+VkBr7A71Q4a4YT+3wMvgthYbDacEQkuzp6mV6qGKN+
BuNmIjEgry1AXj7sQO3hp8mj2PES99a6AU3oZPx69sykA4qsUbqdKdwp2i+IuQWkzU4y3rCtFhCg
/gL3dWa49DWQEcY3+9IM4VKyNz76qloA2aBe0l+8z0i5qhUwXFSapSUJO3zqou++R2mxGv8EiPia
evtH6dBc9/jNJHr7+FCcT2de1pYIP2tkDqoO9vNT1ZPwDEPWBaJAJa3feOjyt9zp6faL+Jr35LbU
NqF72Gq724DggWsgialgsTj/pcNoHTs74Eou03GPCi6XSP/Dd9AuOfqbHGKQAhHMNRpt5RM3thYc
i0pMZ1bFHmg4uMQKpdUIOBNGfYF7SYtN+xDOxil8TK8NQwUcT/y2Z8V4xxaRJaUGJnAyt+q3Q0j+
2gJLGHZG6DkRGv6sA4f2gZs8naGNA8ujwiuAfA8UGPBLCveFz1tQwTSKrZo1WfjUYqIpwKLwdxaE
14c76qhb2DJwma5ma+zo8PJel28ln97GHKc6ZJbiC4UFvkE9h3d6XuBs4KUI0eo5tLY1ksJEudCq
WoMJoJWSv9LMlCxqzUM3vAQocnvZMNBaUjE+8GmHwSypadMKI6jXeSfDmmoK2NcLg8Ro1hiGcQZL
wZfqGvHZRN6mWmramRtL+8Afe0iD+6iTFAax+83quojF/ruXFTwXkbfs+uFdOBh5ia/bMLvAGDcn
zD+PUC67eTagU0m2nXOWN1odbFg+2Mc9MTfrh5vwqh7ZjHRsvkddEjj55MFW++veK5HAWpoMFddV
W+o7VfaIbp9W4mOFFr/QfatMn9TI3ECd3N0Hqo5GA+P4ubLyOKXAymDPgVsW0C95beCSdfYpuDuV
hq+RUkImxy5Eo8QHN1wKCNkCMLROd5syV7IRLtpj2kns97UqrWddWn2xr5FR4kY1pPLpXmc0vXQA
NPK03T98xSqTm9k0LHzkOlEmIBg9fIditL2MDxjVei8Gr4HLsW3MwjdZs4rfneX3iUyrL/kNiPxW
li1HdvZB0ELbHevJyAE6uIIo0fFzUPqcP+VneJHEucd98cZW1cTThJ2P7aC3LKX66tYYhh48TY1F
nIlQr3tjyKui5LAWpET//hAAjfCtg78uVSqvCdo5oFDIUiudnpTzWr82Ne7mVslSKv92iOcyUTeo
ujWAcyGjDBVold2m2+FpTPqqehttcbExq/RrV0X2cgktdwQa50uDe3UbRHyKXLDK6HA+rei2x1ll
ZsU929JyuyRXzm2vOWOp7Wtg1z6xuqlzsPgfq4AsIINsLCEhR0hW1sTMsi7iFRiF61ZYFkUKWViO
GOTKfZvvRyhcyXoDzGA9wUxWkG0XHS1VIGpKprhZtZdBNmRwYgfrDsJGL0B0A0aMNsiiFntkdhrC
Fb5vHQR1kUGTkUXDPljAWkv20sSDQCeRTaeNznoe4INSfyLQTeWXhkb85zuT9uKCFj3E6UXauXO2
E6pxphoPV8Lb/pDw7FcmfspZOw7z08NMf9i/BnGD785AfIZKtz3qEvYSZHgjLt3fH12O4LlXEoMc
PtS+Q+yvFjX6nJW/MLkREYvZXyT6vQacMB3OVwnIOVuLWjheW96+m72Du9DXGtGS9fU2/qt6yGaW
WBtNMwAl58/n84oXIS2dLOZaugXos+fz/QjafTfsU1SAAV1rL0YHcUFpMJCIRgwMtYx5E2JU5JHb
aMl21UB5qjCfH9cUG1KE3/SMO7bVUQ/7Fzrq2fi0DiJBjuFFL6QM8ZnAba3073jn8HvSGZ7ZLtgh
af11PLkTA4rWig7H5AkX2Ar2GL4Tuy5V8jATbVgLYvCxmRtSxu/ykpsIucy/A4KodlPdXtZYSCj3
J4ONyzEUP9C5sgp00ZY3GsIQP93zOti6UIs01v69oJHeeC6/hADJWZl9XsVuoPQPSzzM22iZAwG5
31NBb3H79aGVGdjQW2c+8tEYl0Isexe3q5HtgtRli1Xo1wFHA7NeCEGJ0nY8rfZcyNHw9lQbqf27
fiA0ys6XSNXsCpVZI6KjdpAVMXu9MUYPmECfZuZj/YxiU8L2dwrw6aNPkpelAcIC7fvnIVQNZ1q6
mvFUZ+LRpQ5XFKyo0PUqPP1DfE6ZgdWgW5BLTh4YeExJjCj7LEkwuDk+aWK/2g5fbZDGPU1WR8cJ
xJIk+XQ1oktu7xyqwegoYc+M147uqgsC36GH/C3HuALK6FQckP4+v4lEeNn8vUuwWLDlSCd0Cq6p
ZLpc9TOOeKL4NAg8Vp8YAf+XF8ubkxgDz0RksmzWD/BqJZg+GireKcz8zfEdnunD2okKMkFj8DiU
wJpqf99hqphQrCdAqL9xCCbnGbO6kQxHnV62RHq5VnVpWRsdcJ+YuEaysuKe3sPUQbJnMge7Yv8m
w338JCnY0qPlQMyz+f5Kz6kRAj8mLoMvSRSg1X598NOUI1PqBrBH+SY/A69/3JcaOUOxRe9qhrt/
5uVHzsGfzezdRWaPCJtUrE4eky2o/3Tafe+Avoc87+yFaBOrx5Z5KiGxMe453xFtNpM2XsiHqoCa
1tDAzG66y16GbPvM8Tj02JeoHkYOOKLCSBlAgCA/uDs0wpX6DFtlFgNeo1snnqmzkvUU0pqLNnWn
/8TysZNaNohozS4WkxeRxii5K3bVb/HlEBuXliad7B5OUh7rKc3Sewf9E7guBlvatJT9NRlgvEt/
+uva7VhTHANhsOrGiJA6HX4Lbwb2LN/ArmHAS3l6qymfMtB5eJj+6mp8CqOggfCc01IciK4PYVwE
/cywvPKJ28u//ZMy8ju3iK7YlPEPyH3gP557QQacl4OwVmnSEVN5LTBo3KEysnpizJvqUoJAdXFW
oO7PDSqmARJw6Z4yBeNw6pOpi9Intkwd7K+aB3HBr5CbIf9FnUSZgiw2iz7zP5Yv56wL7qyZ1grI
ltQIYYyTLBy83wR5y0hKzPiQUA4myE0TvBUr/zRp3KEOYZEPv0TuqzVWdtJAmnnoriF60x5gc+Gw
FMHL/4o/rSFBhTmKhUFfm0YZtdRaJULp7mwB64A3HBJcD2Hoa8V6Y6vW4j+gAv/19YX7LHDuPZWb
DKfga6ZYlV31iqesvsW8OcYTXmhwYTJH34NJaoIPAtAojSyxLO/VwIdhAspax4yM7EPtWwSfJngW
pvZRlMOpEz8yXSNdY2XBmDJjP69WRj7ADgO5ZsWHltGd/oP0NL96o2KIP/MIDKGSuD8GENdL65Cm
VTIU/OPc8o403R6cC3a8ZiK5mYW3zSMjv7qi/VCfKqABGJz27TjVZSm1owScK+QnGReaekapW+Pe
dMLV/AznLzK8+k3GH+HfVUApK/6OyuQuqeojyO6/yzSZidXYvynsKLriLdnpEE8Qz0XjxzYYrK94
yPvWxOKp6wjOQ/KtfLRvimZVG9uh5j6NkHktus3UA2CzYJf3XKj6OBxJyfc9R52dKM0a8jwSk4qU
vsqXdRApqOihXYi0OjqGJ0Wn8qGpcvrq5jXDxMzgEpzMarBvFt7jRsX60Izxpr9qFML1gjMXtR4F
XO2wfzjWUzBS88cYEP+oZ2xuQZpx3kbSKzEcPBmty7HWZKDvJbUyUg9IClshIhyu0pM68UXD7Fn7
3cB/rOcn7sPJb4O8qyFNHnk4i4VXBmCgx7kO9dKKjj4asQKjcvU7dPo2t2RJFTnrqDHxo/hqifjm
Au3p7N+2jW0FBnYyx1rmYjYS8igqUz2GYluGOpF4KRQLrj3HIKAd64qCTbORk3L0I4lJeml1ZkzU
GAf45oTj7pmcKhd13YyOptLHVlnXuX7O/EkrYpJHATF7bXKYIZvrpia8yJATr8HNNqo/SpmftEz0
S9+Aq5VOb8mcFRv3A3DMcfTWC//lRKpxJ8ekYGmBPcZfoYrpDOk63iYGtXA9AVL+YExKtkFWK3w9
6Fo7fUPUimKzPpBbZp/926rzt8ruEhnxmrngrieHGdzF2kJyqKXzliRn+l0WliZAUJdbBAxKBQJP
KwSKwhvUyNblM1upSIaJ7F0WcdovdPPDO7UbRZBi1gDq8gtQnvByrirlzBZSgIlEtIWUGDQn0r8A
tZMDl+KMbg6OGND/vn01ECV6HpbJDMSO/gwtnFIFITMxahovAnb7/xOn4+GXK90j21v44D+mzptc
t41Ox0yF0BiheaSyLuqnUGdU6nGMaAAzXDVq0RAsDBrwYbVJDkK3/TFni5INrutgCxa/tdjcJ8go
NT17JDnyHMLl2UFp9DtFxV5A0oUpvh/Bb5wMoqWbJGSyW2kcbCphy/YOpz5j/tOnbSEAzMJLh1QV
KPARDe6AsGbrbEKJwJPL7Ek67rD1xxkLEAbVQa30o0yM3ZPEeNo37zSCQUMuaH/rGYlwKihS+s0I
uBbQb7Z82tRlQb5Dc8p3LYi+tsUqsqsZ0GUmZt1qqrSM9Ev3BqqKyqJo7w/4i7VbPC/7t8P56q2p
+SLpjGtQ/DGUjaeWPj8hXoN9w5e/FSH6DOx8N8FCZGatS8fbsJAi3PVlT1bsxK6Cgp7dGylC3Nl4
4VsIUYBVrExAaDBOwdNFBFlK4Ea7/5k5o/yy6/6PyAZ0ge7FXq2ST9yPX1LPrim85/bh/rvTwRlt
tk9XMbOQQBfxKQYSVzuQiDvAjW8bYmzr8OcS9JDqQ6pQOiYR2u9r0RSRFueZQZCmQf9Ov0d0Zy5O
fTQcWuH75BuYwj4bKv6BATxdFMroZGs8QQ/p04qUu3YZgdXb/Soe9xqqn41szTvqjoxQZAACSSnP
2O8k3XJ2lQ3tsVUvFaghzL3zTOJ+xxdCq564mVLE0Kz3jQ/WbPCZOif+NXlTCy2Yp7oYVJQykIfU
nDde1EhvxTa7cN7O5GBj6pL5oHkONI00fCPAsRpCPsaS+thIdqHmUnJdC9reIzgviMCI670t//A2
7oseWBtQoRKbVUQ5Ds8xBuvSytD9OF/5nIygSaDFfl6stidn+ifButdB1NdPVWonuE/DKqrc5N/z
QOjF41AZE9oT8+2PNMe5JtyvvRgKXOjFd11QgEqM6wtB+I7MrneifR4KHKlfp1be+C9Sq9JvANhn
dxUrJl93xJfxNNewuwlltft+vjGm7q3P395h7fd5fHLQyNReoyvRLQO1h3CkjDi5oCIN0xuiImCX
3aYHBQhfOXJYBcfJhKsNyvH/97m7bay9O4rB1cqq1UD5cLvisxQwvg2emTORcFHu0X6j8O/DIRUj
i1LnTTFiqrZaR1KJYOAJo0B9w4TY6vs1fMS0ZelHt/KphAb8stySydiFJRErqi8KGvSLPjuv0Zpl
UJoCOEELMAW0zJxXwKU5eEKXd1wVQ8rqYcGTFKrlvCuy1mMnNXX/d7RpWiNRpJOmWf56DzR6RXmI
vN9yIQ+0ZULnSeaeh2RV/+CJKjpgvJCPRnrtYyDllETSmGQLlZDKivQsk/wm1ytzDSwWCQaWNQO3
e5BQzvAqe6Q7zTZY8c9EpDm2UT78TPjB6vKyAK9BjMh0DY0balr3u+IS3PbgWncc2abvktU60rbd
56Nu32eOSw2k7zcafYDy2D3w65Lm7ZLz9WuQ2VNI5HPp/ajejMA2dz6DVTVqOYyWV49FWQtSDMNw
sckvl4N9hGEATgnpfDiWI9ClB983sfi+ngJNezq4PPGM53XFhOU/HW6OcCslwM5ja4bKQ4VwKvBI
9mI6mnT3dITBmWxHHD4H73X0+pOY4LOzg6JrmefMti6hrndT3EzBR4mkaq58yxYRkvqmn1uJMPJZ
HfSayvkXYOE8H2ULxG73RwFvPqCfT+aUgG9MmEeVMqwT7B8J0ai3YX6qN+Pa1qN/IQnH4Gbp7XFR
ZUNHyTPsgu/Adgb9nX0rNwWDGsTL/UfndEDurRYwr2GIxIYKbbunoVbLv5a9k0j6kcY+cg4HLcQr
9fQHU6rhdQuGSkOTWNMcIbCSLRmmh0DFGUko9pRpWmvKQ11vrgJ0Itvp8UNOzKjx8aDUZAkPaEF+
t+v+uQPnNVzM2CjO/6LTjxX27kfkQKW8zwJsoSfdeHas9+X0e1wLXSjGyGlFrPc61BqnywvgQc6q
dkf7aJ2/bRDKN5zwKy0GIMpWl/lm8MDw7LaEJ8uSCdXmNUcyKv+aCZkux+kPqxZ0iDhv1pmiBgiM
YYRgr/4ufTD31yKEEUIG5GQxpl7nj0/7y6q+8GHyywkpGOeQWShEa+EOWyytdj7D1Mpd4LnSSSyI
7F78DgMn6+2BN5mv8VtF39tsCHEfXMxONEk6PS9zdhj/YP2penqRYeo8KCiapf0CDo92HNhVy4nW
C7MWUAvtIR6fEWCMYeRsdCfdVrTuX5S5JKvTf3c/71bC1e+pctfKSrCK2rrsw0z4/kD2Oa1wJ8eO
4XaTIZtDgBs/rkfjHSyJUayzPCIZXvfrhRY0Ps6ZStmpNhgoingH/lmkHC+JbjYvYhP+SwdiWFui
aTPnXHNe6LUwLIWgcntRbWzC701WlZtIvi/6l4mRuKWUjiuDN1O05Hp0wdNyC393+TxGGJRNEluS
16c24Gx8xYWz08swabqIeEGeAa6ZkBkIIYbsqv3Bfy/sRCUjeglt9yakoT/GJSSd3vsfm+aCOD5v
hFeBLe83nkp5IEY2XmqP1r7TKRp+DhDJxMy0CphM/jpzGEsOG1npdmUGsfDdLX7tbA7kgrpjwXtE
5IeC+4mmrFfohVd6DY+wzoZPtc9TJrmS2e3ENUDrYGobyuvCMirKZMoIxs5JvzRJXytQ1znUTgGm
CCK7oaxvFrjt8uF1rmzD70TnKymhOYPPKZX43gRD7Oy7YKZiNzI+Vn/1IUF65WfQ0O5eyn8vFNTc
Yx9MBIppLYG3BkpnSjSeCLZc0fMnmxf3RzgL34iKquPYmkNW+jGkNWEMEXq+PDWO97HHGbMfn/gB
A+2YoMnhVN5IBmX8uHjjerJ7tkye8EKGE7TE+/oJJi1RPI3a78VE+aQ84Qp8vYoX4sAsP3wrYizq
3xTgag+EDztk4sD5lhgAswolTmYUnqqvfpw5PabspNXIxhgKUHFr/KCs0U+CKiZ914ZLvNq/1cMO
V0T+jGwoTvwJKbttICX0Fwk4afQbiS87VakDMojl9g5rQcYEa6W8fDxayJS8/X1DBCOoKY1ibZ6a
A0EJPIcjthyQHLBmkuf2pChx2tzbI7mpeFDX92j6e5ZI6osHLj5hdmuMb69daSHDZC+SPUd1kP5w
AiKtVhFNmx4B8vEzCwn/fR8wlseQb9ASFuXdlxSQp0o72tI29EESzDMRLBG2aT+2Bn83lMF9yUjE
LBzVie3xTGSemOGn2WqdOmb/lR6SRfQDPVPnGBVH2+vTx4ATB9aaEFBb2XXoYn7S8mB2ZdmhGpOe
dfi9CLe1iH1uYAvQjq8rx1jvYau27P454rOP3pbW4kYaXfd398GXkyBPsHw2tvT4bpbTXR8ij4Tx
K00Dagghbrh3Bj8xXsLejT/CLyvoO1EDMSl+K8qP2DRcnyjbQX65+4HDb8grEt2apwPptTpIqWk9
X56mLA4p/gqw15WfxVuNCR1RdLXYPafWDk6k/1bdyWS0/kins1JKr7VyQtl6Fns/n3jyJHCQLUZZ
ttuXJU2PvoN+tR2TninIUq12jzPk6+iejMmSJv2UTMheCjxvxNXjQiumKVbtsbHZKx5a0Gx7yKsO
1PbQJBuGPLwCYbaoK1BFsUm8jXQuZCuNQRi12fBJW5EEjgjbO2DoqFlrQYceEQ9Qtmo3rN43TJEo
Ez8ZA7ubHJjiM0TZYgreKNorV0Avo/V2/I8aZO4Zb0gWHoVK8Hwd9tUyrmqgrUUG0VLHaBbFLOhP
axQMZ37QdZTn5NmfDkOkkBLJfWg5UxylFDVq28nWh47DmPQpz1eB4BGF2oJt2vWAwo+JGuGOW1KI
QbeM5hI8m48E8CCogWxOYBOe8G8gNdHPdRZhtcqClfCkkVkVAKS3zm8lWDTdpUALpwe+8ZZgxgHJ
aTC8Zv0XZomgr5nly3X5XrsMorNU/MSqIYB9JQ0D/auXUPhIjEEOWhFGoPAFSGyJJkuicD5cWjuB
3iOsChbXvTLMCdE/PAGmYi3QJSiQ1RJch+3cQrTArsWaBgvAxWqENsP8lpTfUbPNAfY+j/kH0J/V
jF/CVDKWEvJf+JKF49glEbpwz+wa+K/dm6HUrCdtVDyt1lCsDuMfw05LlfWDJSTUhmdsmfhmItTy
U/rBBaQ3ny2Ftsz9iW7sCjlBsJlbKuVdRAoP2+AGr2JvTTuw1R9JcYoSLl6Fbx7l+X9HiBtTXigi
ojRmkfkCk/7XNC4MmX71C/wJbnrlVFhQLSbLyRKZrACLifFqUo8ddoT2R54UJCfCYVBlvVVNgVeV
bJrv+MPLf8MbfSFFbsj2vAijzfG2/Ix+rIqeqnEB9th9z2t4yBP/KpRNXRFZvxiZdodXQOPPKg4C
AzYV/KIi3IdLTJYRe8u2lGTVIgGdDMCep0/kd7DlMRgihIAK17pSxgygvsBP6TeMrrf5Ko+r8oak
IHq3hlRpihevl1qwqKa87jkoBJKvr9y7OiGA3IInKbNXpgWvjjFiNKgTaK2cpwm0KY7ta7laYohR
0A2EOR0xf6irSSRLE231OkKbJrPqGt/oRtYiqW+0W8iOu9xurEbadpHs+qFVPohB6NKWqcJ8k4cB
qFPveGq5MbWOAydRTJWZesKtAKTfhQvNIGlXy2DhytpMQtZnnpLf2Xzx8eYnY009GniYrYxkz0kb
vLwZoe3a/3Nnvqe00VxTa1dKAmgTCTDAu2wVgFSxCMqDEyQgwjxUFRj+ax8JqvE+2mQDnAGsgVn1
zKdwnn0ijZIgDjPHF5K2UW58QT5TvCAfJxfftbb5eTpXhSToRtM6n6bY34tAllsldumXBdQKytfZ
QrXvWqbSfhMK43YR225mrLA8yZl9moeHrMBrJbwlbdooZ0XJV7lnxaNwJZMGdNg4qCIKjIHG5d4f
CInFTk59csBYLBMdLD8HyK8meqiDbOUP0qSnVfTKBLZyUG9Lwh5UsF1le16Uxcas74EUTRG/meBN
xlnuCdDsTrtrwnCoVR6QEqyQP5GvFe10oxktWwOR07N3WyzW4FAZq12iouJ3ldx3Xs/3m+NQJ+Rh
S8DoOln6IBnpBSaPCoQ0w+WzcS2fMZjQFpNKwCyf41E7qf/5jlpivYi41r8kwdq+qSGGxTgfkOa1
H7LthF0727Gs7hGibF25aGMaeuHQmJjlhTMo9A9BS4HZnpcHUeySGPY6IZQSLjY1LRdcem/CoFoI
9I2blOHhlmVMQS4c5o8d+fdUUYM2qbttQI0610q31n1C99TCF7GatcQsIBAGiXMt9cRDqN1HhZwl
5G+er+Dx5dSF6NVFr90hcN5aKftISFGrPZQLjmkXFCY3kvkcoq3VI4q4NolckmVIjA8buAVYGxDp
72mBXpTKLaJDF4jNDEaaBRq3gq0McDLqf+m9TAsxGRdvW4H05Y/ERQshlQc7XARZIhKMbisZiXtt
EkZ0g1A31NzD2yJG2Fj5PVWZJqdsWlAR6fJKDUkUuhhZo3LFCLG5YVfkJIQ3B0L2sRLwbx9OBr8n
hJrl+XZpCN1jGYIV8+5skeqUAdWpKAr2ge1SPaJeAMOOYpBKVIWZgYCNsqmwmFlpoVUbObPy8O6Q
xR5FaaDRJU92w2kIsoYTyzW65VW9WpTbaIzkLR0I4D9Qc4CCGv3pp95F8APqNvRrkwQfl51tK0/a
4YSWz6DJHX2E20dfs1nXJ/Ish2OLGiy/Z90chBKZcyI22+l5/tdjeD7n0aAd+cY4J33zHDwVCaU7
divJx6CRwlJUPWYc4RpyQ+MB9EuCoimUtF0qG4bz7zcW7pk93EHAKlcaTS9FoMr0jsC9S1ooZGL9
i5RqxcaLgFkH2m17yMba+b3TCjrAHavdj87a+K4uFLp/PEUeBnlR7BgubJGBHO5HVa1gdPwlaHBX
I8c0iKjRuIKJRc8wCj13gGfk0/C7KX6SNdQHH7uSXwDy9Ilqj3KjxxR7QlSBnxqUy92ONkGPzj6p
g9SpJ2fk9Ovk0tW58g9r81ZdEZKW2PAjgULTt6pmeyx+W+FNHopNjTJHRKnh84BK/mVEDr2gNDeV
5zQHkFnosyyI+si0XZmjzu/5jLEIQwMUAwUUYbfwVCw7dfmj/o23bP+SGKUtjLkHleZt5VIYimsS
8GSyXXsgX+CQkIio4VVno5m+z7BwZ+XzNFmaHXDVnIJcAPpsmjYdi6EQIBdpnoj7aNr/wgkDvQUt
Z3XqvCkD9S+oOTmmUXlp7VKKGXqHlQKrPv717M7e6hiYhTAaveux4pP9Lhbog62+lgMKEq2lwzqb
NIQIGF3pUEGXsDsfESnK8XCg7NzVQnth+iGwvIW3Zw1qed+HJAVgfKzYVsEhPQkkSB4mwT8Rk3fa
eVxLjy9nYqij2vyI7MAPyMR2uS7bNDw8AKq7I5JA0wND25a7NMBsPtfawEblTZzwAqFsRmNx0IYp
xgfdkML9fI8QbuAq4k0xsZQQiO9oug3lC+GX+9uAw2gxjhArju5KrQy6N9S3/aO2g4rH0Wlfc9Ar
t/GyoyQkVcSRlQZNhTKXlJHyjBFyaJ6nWjUyvVawCiIGOCkWPrzxlkU6Y1aOqg+7UPzK5APzSl7F
hZpmgJbJM7R+LOAcKY5LvXnSxjD6jAfF/ouPMWY3LUztbr31vHda7qYQ9iVtB/VdgFfFX0FmacwW
XKzWMSD5MQpvUlcy2KrQmQIv278idKBKOXhvFjgoPmPHAn4dmSjmHG3xerFXlDoKK6zoZfH76e9/
miTALuqiDU/eEliwIf3n90R3ZW7OsOdCSopxneox/E6WMo+BUIBijBQ7p1pGdvxmI6DItAw+8ng9
Lq18x586zo3OEbxHwCVV2rPWXtp6DdDLWTTnSg3Rp3zVTphM2urkeSbDAJxmxOAvuqrE6dPkFZSI
CuR5HLNpn2HHykjS4NredDK3RlUGS8oJmC0Suz986sfGhwwDbsvBEaK+94SpYW/HEU3Nw+uIphDR
Aw+lh3cZ9FjmKN9nk3WAAduQWNS2jhzXaYuDksoMLFnORUv4nAwSCtQkYDakrK6fzsqxLdXbxu+Z
IcrB8lJWOFUTbG476iNHsxJlVI3hj2/6G2+2dt2NF3V/c/lwvh8vYX4gVP2UCUrX7J960SktDf/x
UuipDc3LvoNgfzBK3w1K81OiJz3s88shYi5EbG6ZNsau9SrGZG6LyZYzp/vXrXGA3NQA0mUKRquj
6GVST78jCXdAUcj+LWq2yqSDLYCW5AeNCA7UnuWPXJ+UVuQh760r2+6u6RbR3c5EvxmNqVWGPgbZ
ZFaYmxhhzYmrau4hfRnrzwjxBd3K+EgIC/PZTm6kmmcBm2XCbUdJWkFFvo9b4Wep7u0Mksk3ueze
RGC15m/0k8foBC6QdKKEf60HYmeEbBVuV7M3on2LjwdGg+YApOvVcLSiMNA2Fbfw1XfYpctfwOhD
4ieQ0z18fiVZxpG4Ge0HVCTLTgsNasgNHWJkU2u8paaf/ZSTzvEjVZoAlrIyn7UuUQ9iPuYtvvfM
Y352qtUNXhDY+SK1HRsp6E+R1lknpZNdFEg/NN40DF5GRm1T7/sGj+yiCTR25LPmkHwpWK5bbn+7
5FeEcA/70vgV8Z4QqweyWbPQ78qbcxy/HUhtQ2an2oXIc/AMQLqk/64WbhnZbZP3ekUVMHaImip6
4XjdsgVy6/Wvz0lhZMAQPAsE5Y0939Eh2CamGDgizjexV9Mmegb6MniHPw9ZCGWdtrnmV8W3z5om
u8vGAhAQeusUfvUVmbeNb86Z+oYjnbsIkfkawY3NvmRVpxZG5RkTt69eUo2yO5EO7a5JhNeN+QZ8
6KMMa2WOU4s37p6or8yGRR/5rQXoLwR5DBtXOU5fdH3FdpBZ3fQkMd/ei82hYua71K4cSP7XM8O/
WrnznunNNvmm3vTE7l3OJFCEh/o8Z9wpF6KulGEPZPCCpHgUL/rpIp4dikLG5ELKn/z4bWdEO3TX
LRIZzDG8k6uCd+RMP7btJmrmKHOxnxQC74w2YsUEeJQXL0Y6vxoZBr41Hngjyr3E1uDRrDEpQ1t1
IQMXywDxlw3vLDRqG9+BZXUmHjA090mYaZ5eGtoEtwQfezKeG+3tVv23NQVUn8cXZMb9cVjSRnjC
CtPkfgpSnJuAnmPMUPUGHilbkQEXn/c62iFpV+vCJb3TJVbBHyy2euCTfJRmaS7hCOEYFEagat3T
j/9hJOewEakIGdV0tuU2ZMSMohTb5CbYAUMD4WmNFoZgPdPLfgdNe/3nEfyd2Nk43TFMZJ0foXO6
M7MLmeIOcafVlhk+0Tg4YrSWMSp12w8x3pk6S8rsREHi9tei/0mUVHIC+lyV7G1I5eNla0PndgxE
oFnVzo8pUEk7JocIdyIRDbqwNXkzBUhdSQT4hQDmquVLbX/SoiotuVySwYEwNmmSZZzARhjqzP1J
q2eSYyzgW0Z4dfA3O8T1n3F0zlcGuaVoWt64yrhkmEcAcjUWUfMCdSUvKCBEVaSv1OYjUEOpcQ4t
66+8nkjamZh2O+7nmZqsRK4UHQEItGr+/2Y8Ikwt/chMtLIewtW1KGTe0T8VH65paxWYGoPeXRuY
y/cMcN46SJF7Upg2ia+RCxuSPQc9DuOuT19in0PiyCXzowqE+rKP3J7N2Iu52dSw8UFMNbPfKsxq
DiPI+JN5RRdGw8/pUAaRecK3KrEoRcPEQe/ryx5m7y0gn6O/xkM/Jjr4+KhwQPY0UcUiJ8m6/cPY
17tX4eiZjE1k/tKMcRhuQqH8Sa/tulwb1hRDEK9nWREAJ7pINDh3MLdmzn2NP9wMuJPRpOb4pArE
7nAC9OcrMQ9HwMoXdCBfc8jAbXiTk1KA8uTq5DDIw4xu3y0MqKyfCRGk1DLczFqIoF8ZNRdOgPCG
hXQJqYxnXPKCODCKmX9h1z2oDbpaZMLTuzt9BLMidKnXyPOIOhm5WZiuwIbMIvdASBzvPJNb6wxq
GuuDR99KcSpwehzeVX550fH3eL1or1/1iry5dtv1pW1z89XiC+56j3r8Pl0lGXB5wdLIX78ukcRH
yJTLPttpm9wEZyN8obKOgGLyFCCrxSFlJSWNAxyLrbwx3jK9gwlNJZ7dDWcjHA0JPW2sJS/gwljg
hpILiI2LyEXJ6Qqz5twFQH7oFAQlH4CAjWeMm+lJGFwFQdY4Ms3vKI1zwUXqKl2ogFXeS+iAlUXW
YtmAS0gesl8RsZr0RFk6zy0YQLqTwRaelp6SWejTdP0hYYGqGGxO4arCXikB+4jZslUb/6Vx8Cie
qDZBAhN65T2Xb/WMNPcm/ShA+zWTCuqniQc2gwfz5s70bAx2pKVZc1rEAnKZjXSjt4KSxPtpL/kd
SmCVfB9DAXqQt1esmoU/xYCEb4QHnNa+aptd2+8qSFocQMe1QHv+FpDmC4VIeMXx/vMmCsENnBp5
QFapvnnwFMmiYASSvk8jiMut55vugSMGNTZBkXd3l2YPAKnTVvWK+Cn7s21cHFzfmkw9F+4uVo1F
sUB7U+8xH4pqmW3fGheALzojehIJC9MOjzT9HFsInCKEfAiQ9EavWXITtpIuTQyx/zaK63wGCj0w
ZxnF1Yxuj38+LH/DonSHZVCtxemGZ8AN7b1vDkPJf0He4zep8e7sMN71PP4IcSSKa3u1pZc70t6x
gRf1YMZqaPIJZ1t//c1bEX1g+nZMv6jdXrUa8ZUXYdr3aWePehJDX5FDw3O0ZThPLqlbFKdKC6I5
T6vu+8IM9gNmBWY42jG3lrXwUWf9BizhGcGI5XAmxvYbuJBX0EyNbw9w6lssR5ZlLLb7r131NMHv
VRy8XSNIm3yGDwrw+VQn/VXjJ55MrRe3nl3p0b2cE5FzCYhmHfz+cKCndI85oeRhYbhj7+Ez0cCw
xvB8sCDSu6HqRJMxp62kvVpDsBsyRGSF9ACwvIOdUzWRX1lpzcCPrg65P8ziITOjaJY6a+ZrSp5b
OC9Ldca/xCA3sNzuSlUPFmuKEyRCH54bG1UWpBxy12ljIu5syjMMbgVBtDQDOgFOfifmT0zpMaSt
fzFEkVTpYVjP3YZ/l9Sx7ZknBvX92GzqdtkB+m1P1NwJFolkGuuKSThbAg+q8lC+DC0PEIOKYmx0
mOZY9HjpeP7Tjq/Q3U3wLdnWLC2BZaiBvRdScdnRQ24uzqoNsSKGT6Dm2IBtVTwRwaiJBu3E3DKt
153JYpHYpBX6zEkKNAeuFjTcJt9qKWTKbWvJHYwILfZjkTBgvTDHBmB6B9NtVKG5ZXv5QtI5P14w
PWE3B7Q3WJwobg0ubl8vzHnPkdtL0e6E1Y0XKIyEaXZtwEUnDOqm1BggcUP22EH4Bw29WMxOqdSx
OuZZ/C54dDlgwXZ87BoNmKVawlagL0VAOWxn0xvgqY9NaUY62wBriZ+wry2IWQnf/bURpxQFSTWo
YfM1uuJ8apjSuxRx5xp85Ty4WHBjIIIEqHpeM5O/ChYwnC4L47dLqCOZZqLfmRGuAQld+rR2F939
rKrmuV/YYp+zZArecLp7xN9+mK3RO1SYwhH0G//lTip6DjuWGBSSz3gjPzEmXxmb+/tBOu1VrPCc
flKSCJNAaQ650jJR/YAj0qL5IeSY0LvEkmAWtSlO6Ffu8wyZbRuE0e5SvMENybe8baXBbHe16yqt
lJmISuUh/pVkD5VwG4rTAuPW18gqh9+6lPKNoZEFas/CXnyyXLQVBef3W9Vqli+6YJFuPYHasRVa
Vz0ykfYmNIRpSg4YYpoNJTUhc1xwml6DSRCJU/mXEyCcg4mJO/Uall6aLd8tZuL8uL6Xvr6CLKUV
O8dt2B+JuVrCxAgJE7K5PTCP18GG8SJziXIbS0aAgk49rRtTNTXnjPCIlR9jyuLVT+z5swDnyq3M
x2EFfi43OjIXQei80dX4pn4AsPm62YF+uWeYvNhoZwGxAXHMT+zSGulBlUXKFsMoQHtQZjNAu9vC
XgVtpiwMOVNbN89wCUi7pzuM/EoPHLluqqDs1GiMe98KPeSNJkQasqoZnKgwlZ6dNHZ26obDrcN2
8zuHQikwMbM/BFGmmo9bFlS7w1do6ylqEsI8mhp17IvIxjtILKdHZvg4kHDrxp03owvAHiEebu0p
5cyRwpRVIwgYwZaF1S03vnhbXnwpkPPec46RuJo9/w8uRk92yCeahbsrL2O1dW7+E4yge7SRJ/of
e/iYZ9m5Hiz6zhWeyUP0r0MTzkFFXMl8OVxTK/FKLZ5U4JkG4XH6I+sSu7Gpmp4hSPGATrbHPvK/
Xh94i5sy4mkSWIaR/fHzlC6sdDeJpIyQH/bbPICTL44I/cwaiM9wq9OjNTyhng+tc0ij77CTgVuS
m6sF0Qfvwt2irgP/d9t67qUaIOyAbb8rlXOb4Zc1+7cqhI+WaRrTAwcwQ+OxQhdYgkXeu0xjWNQX
vH1sjfBrdxnMBacQSfP0vvWXzErfx91DDr/iCuBiHbXhmT48fVEzkZ9cZdHktLDdZTT5AOfT4Aus
uUwGUBw5OiEUASyM8n56beleQUuLssOnhBv7+ToeBqLALKX3jq7DjePcuWu1LtEqZatSzQCvM/gA
4PstuoZByJrKOjc2lzPlmh1AC/BIdBhol0e8KF03bmYlIbMBTC4QMaYtsitmbRxAb6RRjSkkqEMU
vRe7oCDiAto5xnlfRm5869N1j193L9SKQ1cQWLea16vR1hYRPcXIXx8y1uwHgDGS14h7TLznnHyv
DcokexnFNke/wV1O7l9XP/c0R742hTzIF6cIFut1BJzeiosRM8A1p7gOUhV1ssTTSuXBGMyDtKD0
te4eeJemnjdi+BTzOCOEUMdwXlMQ6+3fg0vcvntKZhA5YfTggMg01H3jgqKfYtutwgum7aJiA4tv
4albTPvA2Z4J3tPzd/MSlCZEEGT+vieOF30TRaXRdsTyA6Dyf7TV1sq4s9ixMHxCsOLBbI+ECus8
md5crxEKtg3TuWCoQMpwpxP5VcdMUBU2AF4fuqFljyviTUvK2ZxsKUw6lp1nmfTTvPfA0c8lKAeA
FYQq/nCV5VgSijwaLv4Hbh+qLl2Bq6+DdJqaYpA55cnvM89Bh2eK+bh/yuYa3R47ZAXhbJHTm0Ph
5tV7T+h+zQEaO6gXxiwV1zEtis5Qg2NNYyLkiObYtoGCw/Owx83jgZwN8tV+l72wjMgUsfaRrIuG
wdfnoY0pP145ZjAmHaiHuBMgNNKr3W1tWv9IJNuA2Lt9qH8XA/GBU6s985V26qXVfOhiU7ivuANj
X4Gj7hLNC3KE8YZ8rWIrZPUvRgVSmUYKo249kCMidpyEHa5kDKH3MwXQEZdqJg6YH3PiZmKuzDHJ
05mY5K/s7lZH/V2b/lPH+yRvgmJpOTRKAiCTTcDdatYujvjqc8wozfzrnSGCesUCzDq1n9+aw8S6
Yd9FFsWVSvSyWQeG7CqwOWHtUSFxQmJGWmwLyysNaB2gUcS+JcQa2cU+hYTQmoMpYmht7xNZv8XU
n7zbb/gXf+q6qe9uQthqvJJehpLDxtb4/FJTIWbS2JnNNBJwqNRvyt4qFJakMwwyb8jNeZ2OZCwL
4RaTj5DedXVDdomI18/7GmqpmMGdIxyI6IC1xtJI2n5m5qWu+nEVfzcA+sNqNQJ2OjcLZnF0EOMR
Kt+yJ+RgnjsikDquS+Wng/zoLwDFksRJPxyDCCRF5r5ALN6K/aDHKQ7+uBgdm8Qk4xsIk6U5xs/A
3gwsOKX9GINhVH8WMbHG7Me9+UYkoibmCCYQhZZwjTo4q+SdIXCxtb0XNJUjgJVVYhbxKoePxquI
JUJ1G50UcDsGkVUfHAc8sRRcPLGgLZpR94PDL/wz6IYJyVKilpW13uOAfbmjGZNNrqv/wg1krJOp
oBV5EdU36fGl5Lhe7FoVCfBFK373SYFaRRTVefnm9KoE2edCWurQc7J15d+0TtbSAdPVZDYYlTsG
Iytl+bi1vPpfxZfx4yrlVSsSCXjWbRRXxANfjbRl+COYRxHuRL9CbJAjACRzQIbvUIpNuz5i6H4G
q0Yo0OLLYgqDLjEXQphCEK0BDzWtO0VSGkb8i/w9MhJDC/myWwn2l5c66vsytHFqrVqIIVFsdNIb
IPsNLydpAJgidbcHy5JqRLj+tzDBGHgRnf5RoIKaJL2div1hXSAEIYUODuSoOTq175l8PwuOn5TK
OD+r8agSbCkv6Hpkqzy7Xae8KerBWtx317ugMiThhXVetvfY+PoPl8sfD4pB8WeGV23r3Lx2nVDh
InjYtdzKe9pXWVjPdK/PBoZ4N3BbGpTdHWu8kYjmVy9D0kSXseEsehZo9hePy/9AhMMY76TCJMsq
kXrN1BNNGPM6tAZd31j/vNhS1cYGik/4l0BNl3mppzAMFJs6LC7tp1D+DlK8Be5eZ3Xh0lljAzAq
y5apzjXOSm3o2aYqakh8dHG7YUZw0kb7yULNcMatwxxtZYfsuWMwy5D5OSuqP8D/EK8xNwMZXvHs
nuJd7UCCGEEUGBoWqFAw0LCreaR8pu1UcUU58ATzBEdeIPFpmSkFls/VcfU05Oz5tT9O32auCrHL
loDYm0gSJCrA4B8LeKwARAm8B3gQWjSXgEbj8fgmHNUu6Cn5FicV4IJsivyEzaGekuYTKPEfZIwf
DKXKGKfY/hOsaSBF+wiZqM49GoDLdI3gAZltCvGVfZM1PPyVvvhdDqra2DIdIxGrA0jkpPOR4oJs
9GqTycGpil+CsIGVqXVssdthfgfRoV0LOk7NuKmxUtsaFShEzmUNYN+tHWX5FIrhNasciH3C92oo
8UftghzraBwqTCl4PkpiuWwNn9klI0lp9ElCkvFskg8meS7R2WY+EvfafB+iZUFadQWSWyGrdR42
how2OjHC71fr2EUu2fS5YdMYqN9FCABLk7tdTiNS/IcYymLGFLJoj8rl52OA8efLTJUGcQJyhVFp
BtSxzQk2XZ/PnqwFatoZjDXuYU+KR261HnZQ1t7BB7kxSg2oJEvm3TgxWzZeGlOsdewQimfjXEzM
DKE8kSXQVZWUEm9CJLQlX8Q9NsfHm5bjT0NoZ+yR67HTXO+OiI+i3c9tIeK0GeTRI8HujXnQNMwQ
r46ny+NqvVO73hZgKwM2tAFtC/gSpSk7fm0hEnKlTDNqTyWajdjcdJoTuV3EHmfyHiKsfltun6FR
lpV167EYCzT/nY/LGSbi3UZ9Jwk1YZWwV2TPI61fi3wDOFzmDKjlO7+9/2Hw7ZCRw//lhV3f6F2M
1aUITGJTJbcMlNKhKSRPI59glqab0TO2jHpsxz9/Vl17oV0WMsVY7tGKnXMM5IkS8SMJEEpQbJM5
YTwbU/ckfl7+yUfOjsJLOaMlGriF4OW+ByMl7fE3LNHWK8XHC9N3AFb8VKgK8zknPB/uRMaPD9RI
JfMp3CCgexamB0rc7DwC+KRj/YF9W0xingTWeeCC8Ug3Pk+AfdaUC+XdC+KzabqUqrNNPj1GdWof
T1eNJPkgKL6PGGpyT69pPKQAGLjVLA4e5rSp5a6G6J+Q24dTsj6Fm4NqnNZDN5qXdg0kY7N4Uhml
cWgBIZ4twp8+E56er8apE5ccQXjXoHu6qIA7qaEI4f4PjTDu+sfkm1hBUDwVtD2ZLEGjhelsVSS0
PUWR3O8QDKYp1diz+fQcjRN+eyE+O/9MOVHLG05mrXVyNlc+FvDod03oBW4hJSOOOZfFCFsyq38j
bKGSKW5MrfSsRmkjP2fIpTiof4ZVuYxcDFrVH8KmunziL0U66uiuNJSPR6AvXWc21cAuIA3dcA08
Sk0X9wiRaomJZJw9PnFKe3ez+9hnGGEsfQMWuGrvueTDDQEcZaupBZr8TIDrEMtgOM0kz/XElD4M
4zZtH004v3VfAOHAzeFy+MzR22UUwDXD9Bxv1whaB0uLkZouJ3fVYCeKDWFO5M8ppHHTxhBJe2hj
HlkCTI8dG07zIMDCXWXMJJcqM14z29wIKh1d6WEKfV+4e97WsH7+HrLpt8jQDFCc6a/0RtqhAJP2
IPg3DemJBJ+ir8wtJYq1xSXrdZ/oJT6s/9flT86QHx8BUxRl10VOEJxbSUCQ7zjBJsKHkV+UDpZF
xwN0yzX2i+LL+q0XIt0/eza8PyNc1xXuNS/OhQbklBX+c0uMcO5KTEMs+1fEbiNNolimCShZrUNs
bluJ1Yarf8u/x2FEg2fXb0AzhG/4jVtTqLpyhL2ASULsylj28ihLDyIS0+ECNG4IwuHj9HOPuJnh
MewQie6DW/5UMx4Ao2QilQGYJaJ/czLcdkpw629o0LKOTOBw7JRFn/l3vKiteuunQGkT33Pi1CaS
0cFDWgV34SXBQJJAvXa/WEoOKzEPnsChKgPRWbz3TGLzuEqwue+WPrfjkFMp8ZLcJmQMmD1mQsLm
KKLKVqcwsMXLZEWVspCbUUgIYhJTqAc9tF8PVPN4Ithg2q+8wV9DJBGvBusPCF4nNjH9UmIVSKL4
AyTVkNe1qXD1Uc8wOoZNPUy6shbHGqV6LuSIou9FACxcupEiSXsApQUsJw97w55An2Pl6Kfu8oS5
M0PGPeXwf4P2EZCik8pmgfSeLXIu8saucYCLCxYKgYmb1JsUONGVA8Q4TnNNHYHRDx1z9x1VcM0L
zK1/TgsOCY8m1pxUq1W4KrRljw2tw2vW05xHoD1VXOxaiL+tMlZCXvA/sVe+gVrLyBbA3OBiJWbd
9w+cUvCcJZYG+5YquFZInh9GrGurFqefgG0NJzB/m3JVmprp0HWS1NrLCp/4tpmYMMFyIWzUcntl
OrguqVuxhnTwJ7jowlsGCzu1lHFqQYyFJhl9/Hdc3kL7Ids3hdhM+K1t2PzXsk/u102UAJZqFbVp
/kzYBnV5BqIyE3ika8XZXpugYe503129pxY82y0adD7jv6zwgH2Sivk8hloSFlCr6FqkG+h6r4fY
E89JY90EtXMs5GslWC979TErsAJKAGQNJ1M5X3IrUl6+tAvOZwp5gsnnW9jOg1As6bHuDjzFXM/w
BXs7ouC6sFZ/84V8Db8UsZLVS134WIkuAbRKuW5bgBzEdTgpVIOB5+z1zwf03E3WhZXZQAJ2BiI6
kon79Oqe3yfuCGNaLQc4hFdQgg8NJh/NB0xPghFNogTvGNDVnegwrKV1VDHkE85i/zpsyBiJ/Ddw
iSOvnnu2kCgS9YRdZ3jmgaQZwIswQurQabxOCoYTS1MJgA6a7F+X60TIkFmCvkBIjLsvrsJIPXL6
qjG9tM6sxh6LVCC8/eYfJIQHwYZ/r3yzUE407Ep1kWqVlcRGR1mYFCAhNgbmPpjgabPDfk+aL9GS
3pzwj7rnofHInU5ZSh4O/Wb5qxtcmHG5InAwzi1BMeziJtI9EHi2hdajAOJF4Weh8e16sMGBT21J
my4vQ8lkTw+0igKpGD1x7zsEat00lPPwdRsXFdWcaAJBU41Jsf1YHCIaCJpVnh/hQ240P8ZRFLr7
blGC44/vwlNf+AXk/gjyHLBRaVQoJicQ4stFomvdvjsxKMBSzrQlp4PX1TsucwinSQEopN9jofED
n+p73XpDtk+riP7mQ01UnRkW83V+UaPcfnf3LpqXFTELwqvkaLknrzEIxXflsNmKLOsvarrj4Mw9
7g+ZBs/hBNGY5YHpChJGJ1pJDrfC6efVAni1SC9Jc04R2d5nccwWvbiziByYslOmSjC45bvWUv3W
A3FDViM+B2loNYMUc9LWriXmNqx8UbaZNDiPSUPthQAsHggDghJYO5o/McOtwCuCio7FYyz4LO3L
0r040tIGoqTZBb+OIoej383Ngez8VJsOl4TzKJ+CE3MTC2wmDGykabuqcC38xTnRdaaalI2xx4L6
Kvf6ILNsPdlll6C/QlwiBBVk5OzTkvUSB4+1pIkgbVmF8OMySi52js0upJNzi4K6QIqOas58kp2W
pfa5z2Wicr0kHukO4K1p6harwHv5ozdRuJDarZMqcs+tHEk5hDEWIrzrvAKNMkAa0BHj+SkCNkRw
3SYFV7i+i4U0KKgXSRJHBRaPENLUjJ1Lj+muOBg00PanXcRYL/+IvjcOyXTklfF25CWwHvNvZzjz
5wHGlZpjYUYapkqy37+vCJILyDSzEsL9BL+bwu+2A3lJ4dU6GgXHW/XiKSo/A1aqCPlYKACqRN9o
njEvUcQDvMA/yMssYbNRwhySli02o+BMu7YhEwRulSb13xLxClF6Imc48WpeIEAd/rMRB3bfZlUz
x4EA/4aWKRKBmF2dP6277HfjP/5QjPzQJ3PeuOs+zDE/x6Qp0Eio8YJ8XQxCqo1aoxWKbgTWmcmp
UwK0TPLXt9XcFbAh9WBOLIJW3s6IWceD4+ELBSEmYBBGwnjOSmgt+DAR1Q52QZ2isC6yT+5NYlsj
lCb8Bk1dFVPgXTGN8eUcQwL+qqP6nFO1bW2aGezIaEhlok5jOwuM9clnY2VI/mFRMcaxKLev+OkA
91obhT8DxgRU0m1TuEaoFwocz+hSeNTZQkPP7yB24mASDq/HaH/OzBY+tRxX42+owicwRlTt/dN+
ChhX8ysb2NNcb0dg+oZJGPCvCozLrJVhBP0z42KOyl5kAUq3EEX39sxxJlTWv5jCzNV6KtI4RceT
uyDpq4AC6fVc8buZ5Ggya/YDjDXNCW0GuNgu+O13sg9X6E9ST2aYsnZmql2c9bTM0ZvUeOYHfPk+
eeyF26ZB2ASV+tgpK3jDrzBVdwebog+9L5EkwQplTtpFx+XwmV/idTfUSkPDW8lqKyI32OB8+8bV
hzTfC2W4XamvhRRdMfsWWPQmz5b3kSTkkB0/adHspbdAiS8qd/ng5BnITA+Tfqrdvay92pJkttQs
7QAshlNz355jaCLgAPoP9eNbgHgrgRJBllNZlGihwzmJrAtikBbtoUO5AQeuQJfL7/FHlI/6Wo5U
on8z+KJ+thFd3o573Urh3HKRyBtH33w5boSzGN9Cg0DEfCFU5/OYrlpx+o4pGFUK3TdiNIpL0Gaq
edHf1z5IP6Jnmo1jSzgPUuI/hOC2GSodGo94b0aMrWjgkPJ1Yw8HJI/KbwWtmTerHThskRn/ZFPl
yhcwexqxZ5CkqYm9ju9h7RdiIRuCv2lu8915ca7bfLjYaXpQKGKl4Gdgv9orYGRpqWCIMy+jq1Tj
SfL9z5hQ6JRWQhjn5RLNpb06EABQ3s0KCEN0UjBIKCzc+bgAxz0ixCi445o2tMc4bu/CHFmMhs5g
dsrCGtJGpcQdGqI8YsGYPHS7KGEaqzWvlV4/mjPJubdZc1aRvusGdfG+W4WZy1DZCWIBkv6d77kj
QJ6d68vflGnwrauasp5X4mIOLlDfIJ9HAAdSzft+UlSB8WHe0Km1iB0d4qRJedf/JwYPulwsllgN
WMJ5jVSwMGZKjXaHS8mje5xCdtzLt3AVy753/v7xhsA3ckMRwuIqG6VyHKFnElY0taJ7326lKocS
mX1wI/29240u4aNAK9L/7k04RfqDNiWWycBxkH0Srm0BX89MuSEK1XzzKb6F9ouWs5kd80rNKuMt
xhrfK3+iNVGmRex+2RSAyqyugb1uZqQiAIehk2QcxPqXLxX3VXTLgBIVdhNQKbdk1VeabepDTHEC
oedbN4ZLrHAeG+YDfqO+mmD38uAZk+VAt51grvL/+XsPL+EASKlR8/3CWIdGDI/qH/Az8snMfS2S
iPDYzeufsIK5Gy0cnv2wJje5cd8BMjYZAlQHVl7a+fdRlZZYASC6RF594dJdi8/CnkEapNI1xO+V
p1jv112ivw4RmZxE7KH6Z9UU2GW44y6Y4rR4UkrnX3qOyX7FXK0Oyp4wrODz6rineWU/uuutelPf
SYiKeLmWmqM7jx84qA8Qxd/ngRtg/nXPabfafJVaeMcnJnLeZ38/3vSRusAkFP+8tvvyJxCXpQDZ
xMTQivude7ytNPCAHle6xOVL8iUvu4SxRra8O5ucmFbKKgqaqjLfGOXOJtrQXt1p/FelG0WzuTp7
JTzaJZlVin5iUBJXhLZsgZvaHEN2Gde8T3fiRJlw2rMsUklQGnFBUcdW3+AtL0N0mHXIn3vONPjp
W1DvSAIGwV1a/r/9scDyW2XUF/W4/4fyJ2/3viVHNr90mwnF7UmiDe4Q7Z/rxIKPabj7blTPT9Cn
sqqWfNFuwsuJdRKPYzV9bvyrW/MkIf9YlasSccryGGXdpg2HtrYSupQveA4vy7XnMkF3OhjLhx5+
h2//TFI2uY/76VeTJ5tIlj8Yz2VtGE3LmORISLQ9u2ids0Led+61UXyxMxkcAMoYbZ8nX/MqgIKs
5vrV3ShU98ynvuVWvCEZbh2B7YRM0GFKQE/IOUzsifEuIUF6M98pp/uIpwdb6WlptNkZZa8VHEUo
wkvYjGk9CjdnUxKsUAXq2z+15MhbJe8ySARX2sQzge81U2UhUUNsQE44EK4XJOKn4MEFZGi224CR
Jt9PC0pcuI7JcLRYGIDu8YOyjchuSxUm9R0NJO8yhMQELJAoOTVbRV+nOqk1biDZWzEVWUOu/S0+
guOcWzS+DJEz3n+5Yu9Ji7DIGHC4jMxL2B/697N48Y0DB3X2HPWAcQNX2UBLRfem7ufKWlM3JZO0
5Vw/ycT7ei/QAvtHrsrkQExaHEhS1Ep9Cxu1hMpEHshgg9C/WpggOcsWSb/k5hFem6WSRegbwW26
2v+FSr/65wZUHbas7q5vEVi70l63f/2UF610vsY3WHV8QvFqP8guD4LmMlravLXBAt3OazbclxcT
iVepmk2cvgFyQzRkui2yfoH8pZbUZrEqodIwOkHEqMUedwDtsnTTFjGq0dr0hPr6q7wZXtWdXpEK
dG4nmPJONwL13o58MANJBfaN7Nt0SU+P4P/jV4gwIMjMMpkcuT9OawPktnNbtvS/NAEApYxtmwvf
yV/lEkV3Lh+o73pXRoYcAowINpjmfVo+IVJKXPMPIAxprsVc2uTMpIZB7PhWMlWCooMN9VDeP53B
hMBm1sNXTR5iPAF3cTQCyC1QyNo0L9x1W+ajtxjUMWNaLay+vf4fJqukimfQRWvENGkdDnny1LtR
OE9Lijqo1m74c+7Jsb00Cju0f2GqoZBzBSyQNN1z2iOZTN73kSwlPSqoeTZ3br0uNN3yN7kUTgiK
ZvmV08/Cw789fOPp57bBStTFzjGcd+xZMhmBgPcyBFmCj0swnORdV2vRIQG9pZNpWnYC34v1NzET
OVOlCEVq58kVhlqhJq9QgtrE0g9kz0m/JzaA2N6L1S2nX0JhYnMRvRiDUMyozkib5f32O/VcDjVT
hW4QccCvzz+KXkYoyXBbUK82gtcLCVjHPFAdqeL8aVmm11EKJ5cq3mN9GJwRsggAGMXKs2k09DJw
gbRgz8vXdHF+A/Y2EIEq+P97n/VD2Ao//3GTw+MYW9JV/NPqMcmd6BJHX7LsFH6MZZ55Wt9tpkU5
IfA5i0z8H50tVd77deQLg1kUr6vRQC08Oeuv9zwfh2vuDPPOHpxbuieWoWJ9bOnFIdSIU6kvkqM1
pBKbcjtYyEwxTUpdaUUJkg+hFh5PjZ36kxv9bZrJD67ni2RYHad13T49LIxrQFdndv+/UIqjlG/Q
xqVlsxMIR9sfRupQti/8hDIVtBkpPEzVh/jGYOWwnAd4rZGnlqjxKIs8mz2griLEzm3CHwE4LSow
OOFI3xyLFWZ1BwozRjgjEh9n75ChCbeHKECl4dIqRXecgUa4OTg8cVH3zRw/XlsCj5bTucKIF4KV
nLiuk7GFEqL41nLa3Y6B66KU0mV2OvuN7SJqaJ+Ps9fchQ4mh6EHQZZKJicG3X3GDNRaB9jTvzOG
InNtwdbh+ksM+TFqR/WPKE/9vMMxAq7yvwxjq8ewf2Oi4bwNYghaMtExESZPiKTrqYa4Oo2wMAnQ
MPT720VXU83PFEAHqQFaT7OLT3wSuIVyomXHPWGY/tGY/+KlW/2h2yCqGfElhfJPnqvoRbNa06Rn
u+F2pl64hRsmEvMwWnDQOcbDsX+gu2aF2Ss8tCl785Rb571eFLH1jE1gthSTBzGxFRdBukaUPIN5
6YdwSzRBl/0TxW30xTZsYN44zobE/vOVYcL2GIU8xJdxBTUgDBmqde2+UfG19QzNfGqSpqo80V2q
P5jfpP1T7KWP7yWiaeghJqGF7tHtIX0wVtRX9i5d19TbrTxEMDTqSv3l/XaOw+/P78FuuxVB/YYq
idACXwbX4Wzxevujpwuj3wPYlj70uZD6DkTNO3tvUhoDj9MxckDG02JGMiF54d+B88w7iZXtCiKu
tSn5FsgBHDRTh0UCPuw3pWmO64dsj17E+yos1h4ULPzWN8lF/z67h5xlHFbI2Ez4g3ALuNNqN6ml
FCa8skPvz6R6bM03E7CTs2CThTWDGDxawBUhOCT4qVapSjRQWl9FVyEaO6jsRjleYFNCJtSOnr1i
9ylX7CWvZMISfUSaY07jZlMml0+NhIP3DDwv1I0T5kEPKC/RHyV9zD7Fu4B0GZsTfw8cyY6xH24R
PR2zBUFkDFWv3VeTuNY2CUO/JH0++gwDI5TJSv86Ok1j5xJZciF1NJ4Ff6YRW+lAYlhQtExRQTAX
NP20XMN31FvssBmOANYU8TOjWXIj9hBpLHiGeaJzPzVTl4x/4RjJ7QxCuEIhA92wE/9JCQYcKgFC
WinV2CxMT7y06/JO3uJtyXTpuhP8fU9J8msIXT04bOWMN77FqGtKbJ+7r6YDt1fiPVyGgCUMD1pi
fmlAijJcBVPie4lmb2kvLJVHS3WoPtHkhSJVquWIYYOngyuavFIHFmp0xE0SbvH2Mke+kypj0cWS
bNspdfajpJD4PEFWYNMNJz6qr2u+CZS755xh7Ns4a6CsBGkxkC6/i7oVwy0knWEvV72WUYafG42s
nbJIox/hYqEQGHxGo65HbpDhecMMbfnqgvzCpjmNnC6nfudO4qMESL3+Hk/KMVL44hsdSniuaV8P
CPDurgVdWXq8FVDocgt4rB7vQ05ChV3W0hnjR2WBpyIy79W1YfIc0/B8SOTb7sWhAkPYkhVV1mJd
xxtS4LC7XDlMPqcktElICxaVc1Y2w1T84GfoWkXs06UmkuZG1MMkoyHibsbVbjojUbTB12Q+dmUg
mOmqUUxxbO0gCQRssD2P6k5MuoV09bFQtWIVDR5lY4J+3LDXSv9hEobcrIDHKmJpqEaZSuXGVQEe
j08Oe8qTZDfwbjybUUBdP2FWXSTDh+o9+OmwDaDdgDRqDG4hfRvPxW9CXVN6+Inu4oASAJ+nmzpv
R2tAhgQmnUwAXe8pII41ozKpElEszQdfFc05spyA9Yjn82DIW9sclYTQNmhu3/y5klIJamG1WW8Z
alRxiyYF6YEx78w4Ar5ejFvsWWvAxlz3XlmKxHdWuVjtX3xCaAu5Lz5S4CRoQEQFd74u+pE+07OC
TRGJCQYIycZ8vzuqkYEu+qgd4NR7EZZmS/gYCHjbmkzZukxbftfc5gqehXI8ucYRcY7XzrHcoyhA
N/RYLNwB04/SpSnOPYy/cmi5Uw8QdN76RXLl+YLNgWD/Jqywg9tmnkxt0/4uoYWPS1diZsIgzlie
t4sCO68LaTLKB2Rn4lRrg8o/xSEg9f2vuijjYXTbQtn6K3xOcbouMIoa/d2BA5M+lsBDS1fqAEBY
Mq4Y12iSc6MOV2r/9Utqspto25y14FSEO/GjtL5xwOr50xYIoMi65hpweoCqs7lk/3d4Exki5dvk
zgROP1eSjF8V0i4DbHq2dhhFk5zugj959JLH2WiZJC7Cn8xT2AUvDa1PB+E+Nar2yZFUd61/HnGX
tfamZ1lCbA4fGcVN2ytsEg/mun5uu0Ub849D9ztWLsmnjoccnSViVXwJldFT49Vo98QhvaDILSZG
D2nkemxaD6RIv9wT1umLxh3Kxqu3bEzkMp7GplpjGtA5ygkrhKjQIoA5fDdcN1T+ffrTbJGrJc+0
lxuGPk3zWx/B7+7z/EMsXT5UsETs7TMhnZSFr1ZspXGH1edncvLRA75NEmVjmOxr0MVBWVbEHWHB
rHJ9qxKkmm9dbEfpeclnegkcr2p8akyqfZJMAV8e0b/nl5p0viZ29GHfuRp9Q3FO3hl6UdyzEaOa
NkkT4296Ur3FTMql6IGwe0UR8HdCSUPxNxqPqW9tPALfa1E3UeskAP9CRGJx2Pyd4weumEKHDOgL
F7YHJPAPC75UPR3DGoxfkvQDXW2gt9FxVl7ypEx5RyRg3W1ExWM4fy/d1bKapMPb38fvwsxPWzYA
QZyM1wV08+X4E849pYFYoC6Nruh73wZ6kFbo7KZ0JxqQAMeqMOdheyDgLNqDql/VuMM4fQSN6gyi
ZEe0gY3S8TbVKYO0GY1bGysbjioqmeFaRZ7dqorUBlrpKBKJwZcM69zDTQH1Wc104O4s6LvuoXni
ByERphzZrArzr+ZYMFmw747Qz90UVUmhsFf8oCpMFZMFS19IVG1BVTmgOfRVmxMh7e54tjOmC740
dWq12CpHAooVsbVXKIHaMtKtgTOXzuqOdYzmav1vZhKrlkvcd9BkZU0uVqp6vn0XO3aSaQ6hNIBj
dT/1deIDFM46MTUQEjPbsbtZP3CID/wGQe4Vgz8hzGcGdetZPmesGbxmz5mJPZ87JX78cXwNk+4G
eVFE40+ouCfi0Wyrq5yjEDXJVXV9cUuNBQUXD1JWsShqCPU9GWHBl+Yj/JCEx7Y/WHXS8wz5bo0C
mKb/IvHdwggf8HqKfxxZM7M8SDnzh9RXxqEJh40F4aaXT2G3X+AsQ06PqYgDf1RfUOojXVdQPAhc
RFivYBlYDC2GcSE+Sc2o2TaVX92q9bRqLotleYVi9hJV4HWvETflPfc1ngdV+L2zPPqX/ySuoyEi
2z+I+j10mmoEuLPKqUOEV7b/bNCTwOL19FuMH0gn1+BUaEHQo+b/56nFr59QQC18//S0pyEtXTUd
EW2hJ296PPKVruN9+9IhpGPmpRTK2fjDRyZicHzoiOoRBVi9U8syDcdyPOAG0cr5zihJp7WMdzV7
gADGUnlHj+Dc4yq1lHX428d8WgdUow+IU2WmG2gQGxE6GPd2a3zVlt0naLq4+dy9QFKVV93S+UWj
yn5MQu2L2dkNrj8+V7JJ9HQnotSWpMGjON7IZ6z4OciIAg27Dpal3p2TZ5UPIctv83i1FYjJ/Tjo
Leeu+v4gYuD9jdiYUA0KSZf+Do9xyJo8c4pyvVFq5rydGm3GnvtCRU4hGgdDrGrwA9rqenW/0yzI
/tanTs5ATvQJzfK2LE9owAiYP+tbuam7PpmhcxTomlc8Q40/LOJTxI2h+uDhXPHvT2CPwZa2wWGX
ujV9gmDeeFLyvxoeNmh9LWO/QWtLybZeWWgnSvJxpggDZCutSl1+3qsT739hEn7PDygSlX/4Uz+U
0w8omnpSy/PXc9HLUEFqaH6tMtR5gZpZeZPpTtonSo+QNZeT0+n0g/JSZANUUQb24hpqLJVMtHLV
OFXSPyT92D/aBT15qDV9+FKRzQeIr7WedOxBrFrpWyL61chG+lRfsW8z/xo5vfParxIdAHsAIZA+
sX8TijjZ50SrejefIdqlMufNO/EAlBRuuXrXjg4GtTf3K9E9gATZxTfIsHCnV85qgktFdMo84cAG
MFmsWYT4Ad6rNU/d9MzPGliamTUxCZAtYUUKvT6LFv9H/DYmAYTzOMgH+GmNzdCXJ8IOfmb9UuM1
x60yptJserHE9lDfuXhs34J5EbTI9DJdLQiSUy2+66sklrDrYfEM8fGK37ETZcAxMTeTXUrPr71s
dEc1uR4HHhfB7qCJ2pHV7Zw/Pybs8ZPKIVBwEjffYqh1MPlbxq8IXes99WFqgJqcbPLBwnf6RJYs
EygSbDDnYf/lPmsp5DhdHtv+xFAbtbkG5loQwaWGPRvFDEnTKH8rpKVaPrJIveLKMlUpz5bO0X9C
qAf4CPa9vlY/HUjNiGwGHSWU0qQ9EnLuZ47UbviQTIZXTHPcVbxOMBwzIa/5B334q3oCRrvS47NJ
eeb8YUAhhE5aHqjm0ryLG6zLkz4BKPcFZNoYzF7sw5dnIWH2ocwpZtLNIkrVCJ+RKPQYfqTtdd66
8mgs1SknQW/LydIkmoxDGwfQ5KYPZzCQ9HG4TYVxNOHCHay6FCCRf1I79gRDueYEicTZ6Veb9fa1
UyS0NCKp+X+HUaPKqivBdIRJRfMcBxa9+vC/NxfokcQ+tOARn2P0T92oZYsBINLdGeZSJLjqdN06
ZdJ6ydLNQskp4Dz+ldB1v1we7M8ya6ND9XxbH6cZVZxNXmHb/2o7cVDjBrP5/gpjQf30jJ1EsBeG
yi6SOjmMczQT9YQCs78eqHRt95ZTciL1qhYNf6pJ65RULYvSEoBdDcmBsz1IPkcr8dus8Il+MnTH
zzfjpXsbr1cZ2nKKnTcbfEMfZEHsemLzLnSp1Q6O5mADXUawijLpE9cvYXOLNHX+C5xjkav9Ln3K
JxZQyla4pxXMldsFSCjNFdR6L0XLsjLg047rGQ29Tx9BIOgjgyJAKKmoeQLI+c27p3D6vHE7VbFC
KpyD3dIWONxR7TY1RDByWb8WsgBLam1v/6OBKnJ7VN+7fIm4+L7HjhjTxwDTK2awqXxVPm19lLEY
nAEzGEcM6QNj7LIF1HwZhbwwjmmeQ5ALif8JKfdVN9ajeEqu+p3M1ZSQEnpBh7/daTk0M8FoMg2i
AnOZQLFrIa6m8p2zJ1/Nxi2aob6gjTEy7nfnfKnllj2oYSh0Rn1lQgcoJW0f+SjY5Ao1kweE8CA7
AdfvMYBlcybIAJz1azYqncxKxUSZbqZSMGUStUIoWEvfnRspcD/e12gWzZ14JYpXsvztvf6y2mJm
toKrMGuMz3Wmh2pN8esNfSsed5oTYrt6MIfUnRxqAO4iPDi5/53OphpvCSm0Hb1ZKcNNY0wionAL
OGr2BrpfiNlhiAHrjhfRESMwkT+sqjDhiDM1JFnH9vmtaqmVdWkLncLiIDmlRrxxLVaHZvAprjRf
1r1Rjo3Z+H9tIMDAyqTEhNODLPmMDfgrF8E1K09z4Eo4k+wEq1IRaUnoFtgoc+QeBh8+qv4dWRml
tRSPMwfQ5A0iy1EiHHmEBNE79llpS0dgwUmyVny1QxChED/P50lG9cW4nfhRJY0gVKgi43qmsfIa
giZbJKoEyI6bxtHUB3IB0kp8rLgcaVyoP/zLSH67fDqO3lpHkT037tZi/cQcjNdEhQwJQTy1+JkT
rpZtzZ2F7G3MD+Z5EpbtWarX3WOAddn64hQLGjjCtMBoy9p/7OfQ9tjK6CgCSW95NZFighDJOMXj
XRSP+HAcLyr/Pgv6jSu1j5PzQvao9aWyWSOF6uyiKKhcV3hjBxxgCPfYb/n8FM9oHa8BltZC9rsV
E7yME5p4DDdLtOoYS5Z0hZDheOPg+znLsRon+pzaX1Pn+hN96lpB/Jhg8hqksX//NSk0RNcnqn9O
QcuAxMC4M6xUrzCjkZYDdFeaRwIKuEgTy+dACgdiKFzr1/5y9AvfDV6PVkHI9ylZJwZnHn3UnPBG
SvSdd9aakEjFrD0+9QFr7KzjulncKefYsioMe0R67v9ZC8QInbpoQQuGlLRX7z7QfWLIT3F3gLLi
98xyn/EfR450M4yKoLjOyUg/2jLPO7ZGF08KV8Ak4SxjEmn9AyoUWujO3nyETlajNTI8i1EQR1fW
bntXz4PTds57Dx98e5TL1KjEGGAh61hZ+41Kdyfdx6QIEFWKM8UiqoYG75LG97YRl/xgoFtwuam0
VafDrI+Ngvtl0627JJNXjy3ldzVOXBIigxB82qd35OL7UiOCnsFEaxOuPHuCE6AzAiHSp+bEcO2y
8lcTaR+L5FSaD3zb/XnwubMsphjKbRJYMs7+LpRM7xfyex8CIEGboxSWBMWaxbMbpo6jqgU7fA1Y
6/s6Xd7ro5MEVsMSxc5AC5sj/LQVjed+ZOnnLzV6AzW/iO3W+Id/hVxUD+PikApEwVQFM1Bv4tH5
cROCoAbx66rRjvXRVEc+N7nBJGcUuGMIXKLT5UUyfEqhvpeS1O8y0CpMG6FOGeH7wDRblNK7loz4
Uz2GJJlpQ6maU8TUmmcRHUgZlGNtZxTOY7vlHKKorkXzUxcJyd3Jral44Uu3pfZqunO834dS5w1j
CJ1TJIzY5YGHsQXT61BrFrl6Eej528WzJhuWFEIFp9VKDuUP+2NOTSXbVtNzh9WUVKBAyq7NQEHo
g7M0R/3Wgset09kpCx+ZshM31S2Y0ZPksLc0yPw5u+7K2Lotb4DKH/QSK75uNjxRnYal0nICmNBQ
WIUazsrhPnTm1EM16NAdcFpSzHCVFuOH6ak6prAJm7Wd2vS6Vo6i8MEVwiano1QKQa0/EpfFLWnS
XamMI/RxrDiF3AXeEH8/QdoQh3H/FFuLmF/LKtyp3olaQ0zCAwMd3qZIkI/mDt7xngsIIOUHnwGz
AgTIVftjHFnkDfUyb689AtTrrTdTLqDbWK+IVBHyK32+3FAnNnDQxuxFJyTngEbvhyP4bHu8V5q/
pLyAfNvb2NHPN+vMsTkEnCLJ86rxL9c52j+mPG91feixJnA3Q5oiaX1pknN902TKOnn0uRdewhlk
MkmBDd42Y7JpdS0LcuH1Kr6GWNdRREJs0CIn+0i2Ldq1Tu46M4URMoqsaT55EMKAsZibsYN5Ohhn
kXFdg6/p4s1SBVynfjCY+RIZ/vmvcrs/nm2Ru7vH/k/GeFkCscGinZI96SqgZy0Yyt50Z3bsTv9S
K45mYgZopMGRb+4eAlCEW+bAJktIL+gIRRP+MpCAluot7KEvW3ojF52FinGgyhsNUfMCBx3lGWE1
nRa/aiUW6Ee1zlQ4K6TXfVtlSrZ6Vp1gtEQ/KnDYIrphqNp3yslYY8Lg/7U+Z9OvCrOdrsjnes1l
PUqvjyREULocOXMFKk7pAwKgcq8ehb+pu3bzmB+EdjpkPkI5gM/T8joz6e2AHeHSRC21WU+Qarix
KEAH8zj2St6N+kpm7dMvSm+Q/J62rxM+vCGvDoS50j141XnzcA/npF1/vqBjU90ZL4WHeQs+TOhm
gjDtN97Ub+BxPMfQv+oLXrPbhZpE2TOXHd1LiF5xE4ztL2UXI3Pgpjj2ZVgBvxkiOL4lmhrdL3An
II8q9J5JwtBDyD83JRpE1K/fJsvGapUbLnMM8eH712nDqoGsim7OuSYhy9A1j9c+Eyw3Tu5OGuKj
KF9L7Jk189nOz9bjuaAwEPp5ZJxBMRdfBw9ySXEdW9hemNNWy1Hls0N71D9+yhYwBy5oamUI0Ass
CIl2zJdC3D8mDFJO+FIZrJz7GLb0l/FqFOJWkVDfWmBZPWqsXnwiHPOWbkBnQv5+QbWI6jXoWBzx
ST4IWGBg3JVnUFudCt/PJ3UErFiQg86flfrd7eo4SJOqTOPij+nXycGjnF3Hm1XaMlW2+X+mSrpX
QwQF3k+Wzzp0722MS/dERHaqrlNnWj4q+RD86iSqL8ZX9sLN6TQAWgcKFLi3jsJSOlHmoUpFKp0S
KPoS06uzBGCcBMhQiCiVMxx3wph88on2Pin8vPDD/ApShZ7L6sXlXmLuqnicuVLpFyPKiItVWa0l
TnfPvKIzIp+xHup34qJPXGG4DJD/Q4sw/v+BEYaZhVOf6sbPwJMo0LBbxLboew/aMoB+S0psIPPz
GidRKRtLWKJxul7uGxOynA/YzUXJYRB/wkcNmhsIakzMIdcrmf6KJDDLzHEQDIfLKVBjvkkJX/Fs
ACgl6T7HyyqoBFc3XTn427LeLvYLe9Zad2mM9I2u4sqVaqba1/PEnXT05v4bKzWTx7AalQaV8urv
elLeeLFFOac2zon/XtVz1jzbjzG3YGThmYDwizl58wOcrULdthjOvMAooQVYsoa07k55/IPaY4Hd
J+JMg2Pz+nuqpmeg+PBJBuM+0Vt7KGP8f8mwCDr9EodqQ0J0qnzlFbLdx4qYoWd++Olvj2U0MsLh
PdNCfwRLCwMpqTIusknVG6TvUCQ6D/ekIQec9YetmFw2bq4F9agB26OOBU8AOlJSzO2fkr6zlcpH
i6kyvoBWV8dZf0+F5EAn2WhFOuHCHzDQWMmFb2XqrQODYc8xFfQp95zaJHYuYeSf1l3dMTq2psxi
Sbzl49NvFPk444hJcqgeMvUwd5VENo/SeiAj35rcZG7uhxyZmslVzEwubF7CYS0OsD6OcEzPlA91
cf+UGQXDlX6I/1f5a++SR3wFkj5HGTDjgUBBBiA0jiUESwniOaqqbQytOQ0QmORgu66mFffBTnZT
0wB6pwo22WZ1zygb415uX8XW4P1PEwO8v8AiiVoqATvNnlKCmRp52fUApzKQ1V/ouesJUn2KCaVc
3casv+fdy0V39H2fE/pD+bgczICE5md8JlZ5Rz1XT3j8tCdGgwieZa7BS2G1s43XGyGh742R0VhN
z+G8sue9amyqR1x53rA9fY70ZOcKpMJvspsn23bSlaAMB/3oLHL8Wps1Sc+fI3MlQ0oRrgrocU2c
gQIhOch1xo8zFLyotj57yqWPLqskaq/HGfmHwBagjzekfpYfUrTCe2w9rRHkkwEe3dOsB46CutQA
dPVLCLrEyHbpbaVrATU6CE64WcNIChICK9Yr44IPJBaYes9urJ4+XMl+AKPAQjhj3dOGt+RX2KnC
DkqzFn4DotVQccStzfSJetkkfbLEhaHuV4xgiwilG9GhXs/c9sTGZ1tx5uNcxYdmb1IFq2Q6Keke
Dd9kau560BkxDu5auDKhsToMeYqUg8zWl1n6qp+eP3i5aFtIrkBH1Oe5JUvG0LGR32cXbWcbgT+L
VHFKM1Ct72n+BTVwcuxBV5NUuNOr0cytcxjLebmTG5iWnHcjUjDfuHypI9HgzDOWkSczy/8n6jqZ
KHxH5PEYpvXqIiOriJL23T9O7odHieuz8YvmAti0Ux3wp10cpBDiz8u78q1UWuXuYjpESVzgBdXl
zLB/n6K1W9w3sLObvhXCHTz2FPsKhzXk8aZr1/dN7ycmois0VVysU9qoo+NYWFddMrqSDqyqt6Bj
xZquyA2Qf+PF6q4rG9klwOuGd4kuHN1MUJmApqLfLpVVY6NOnZbaWkJxuUWLMBgTE91jQQ/XjOWd
2UIrzl4CxdQyLxCWOl6O6Oj2CpdoAhr1KdJSV+mDqrpOpifZu3rJM87eZJJO6Nv1fS7RlnxGLngS
kttL+pjMLUz+C4bfd9703J80Th1wG1LfCYdgP/LwOb20qxCHGIymzL3vOb9oNdRYv65KQpIGiPRZ
Plt3tRiJdCZ5GlVfXtB24k69JBTx0GoewfTjMITm1sTKnVSlgu96Cn0QxgbGWlRxLMtSZ7myc3tC
+jWManlJeWqnJrmxAEOLXkMmYxS11pqCGxmfLgwIu7XwQjARl0ncPcv3KEIYMXte7OhopukV3kC1
ZOii6OIWNGDxX9d0UQfFcZAo6xGU/7GVkC0pwmmzHbcD3jTBe4BKM1Rz4jdpkpbRAQJSUFHKooGL
Akj0VAIkizuwLPrCFFxikK/bUFBX0gHr6P/DJjiPz+YN2CUvgeQh9iadyHYM1LA6cCc/nFWb7UDu
9fwIc/aPYiT8ZudsbRbAeiFpQSxg4PBy53NkG171kA8cnu2NAwyIZfHnWUBht3XPoI4ELwh+cEyj
RcdWZrF5Qntnm6L7mOXVMhEfyIdpB84CrexZDCEXZgTqKgmoaONTRyHvMApt+W+9rnVe8brYpj1F
rNw2GqqIvfSlnSNEYt6jWRI/zdYMyifgNOz/8jviRS99nc/zNdReuhuHlcup53wSoZHjOWY5lsIn
fMk0vSPRR11k6cP3+3Z+XfQxRGucSgM5DijZOevAom1HtxZ62b69DiC52xICe+DfoNc/DiFH7kq8
SncE5yK0J5Jn8wyZsd6LxZiNL7rSFeft1k3Xpp3m/7BpcghBTnXMTR9bjW8DTUvxYU32wTDmjyeS
HOrwA0tfemK+wkGneENiEu0lCyi2TWyIztQZsDbK+OIkHGflsrBOel02GIuvoH5iGQp+YsMuwm7S
kcVLtQQN4OoRaPnlFfTU8vSPlq2YOhuvMoPhj+7YFwXDejxfF7dBsXPrHKYzH9gMVzEZFpCUw1mG
GG89VBYdff9jcGoLmE1Wbu/EjaXuDMd7h7xvI7ynjEPotsJNXC0rvX2vbTym65Q+pc99UNHsCWxz
Oxm8nyIacCFBoFfxSIJ+6+Dwwu8LtuZyCyASSRLri3z2P1jlyIQMglQVSdZ9x5Y+SWVDInky3qbc
7yh3lCDhT4c5bgJHr7D4HBh6HiYSu/83iaL1N29xg4LmWCnJk2Red0yvh82aQ+junO5zr/gK8IKF
XpAJh1HsW1f2FmDMjRcHQHoQ5+iHJZgMRNxMhpYWOlUZ50BUTTSkoaWuZLD6wdMNTTm0nZSx6Um4
yb4pskL3pFP3t17kEZZbZ/oV8OxMoQKl1SOQGg8MitghRyJdlzxT9mLG7GgCNWJPqyB3sOz+Gfmq
ZAWzbdTEh59G5SOPJ1mpe1GfC4XmUe2OJIxHMuku71pi+mguf3E37W1EAd15BLAivdSD6g2irGA/
DVyPurvNi2k5BkPW0XtysxGtnsp4QTYeP5wcGNl6ImZbzRjDdG+xzN1u3YDjYfgBZUxYqK9+6+nD
3y80Tcl+twL4Vu2iZpUA8o+hUgZ98L4PwZumIMY15yuIwwznyGGbyBrFULf6h9FZduv0XZnsOEXq
c8f351z0tvEn7Z5N4EXb69yyO0fI3S5kObbrWrBcxEYR2itDaeEj/P3OT/kN9HjbM+I6F+szdSWn
XVpn5aBESUibL/8XLKjRrUSR8SfAnQF+smqBZzm3dUmrQtmkbKAWG8ESVZud9PbdztpQLWerW3ca
1Qv9CSpw7nN6mXja1bb++cLGxF9CoQHeiy7k3TlnVhCgyNNdGVIkUNNblP0W/Y8S2EjjdqMFHfKk
25Cern++gChIcbcYc+Kbmmj6ggwiyRli6B3zsenbRpva1U8SwpqcynJjoaNjsuokZOQj/o52u8WT
/srMWEz80h/z0PaVGOotTGwxNmT8J4OM2BeuXcDbasGnwOMOIwMZMzz1+eCCgfKnAhhIk+eCzHQa
xrvubcoD/AVsF5dNdDOW8W9rGkl1P/g+s+JwEoezQDDZUai9pPMN+SyvTt9pHEBJTzt0G1CC602t
xUVVlGrBwr0vra9hdvt+Ci83aMFOwaM+qaBw0UdM1doCCOkBVFHGZm241CwE1uu9E9zZl6nfJv4K
ASWLbgA5nv0/e+9KtbHwCXMWx9OzzlBOy8IJ2F0vy+BNwa98k1htTQgMw/bfYR17l9mXRj+RSsK8
08WUXJpw970B4zpf9AN4BspuAOpTdh0IHBYldSaQ3pnmha0gqOnSVKVRtEXmw7kWV2zmYqeFhQHX
jCdPg/T/l9zfrCqWefTS71DBxWrZUftigRjJZ+ZwEsUKTM+sejMgJ7PBbGMUd3KtMb8m9EoDO2g2
w+72+CYZesa1onpGfrY766LPIiArGJ/rZ+FTQyVM5dDzXStkCpQDuMxV5IbvyJv0abnl4TEftA4Y
M0PoRLbi5GFdSmGtK3zaSNl5Sy7imhP896OPIxNjRKkZlX2pndBF4WDmSPqf+6IwHbJwXxAcCAhL
02cFvP0jfQtFTYcM4cQSGx6aZJA8CnNELyAQ9W1qasz0CFnNpWaiZ73cFyF20QlUB14+8Prpae3s
vlGdo71KhrjcUspL2/WP5HF4ijtGrcdHiUC4vaFh+a4qpcsqNPlYFU5mVthDydGDZkBzpIzMFRLn
0EfGqSFQpoMkTDHM2+78QJkLEqce/mf840sc7NwXNuCHjgrewGPmJcGQw3YRu0+5E/lrsVakcfC+
D+53tzyU3rhCmSGav3KsXrhUMQyp6odQsqS5zH9uP+bBd3Urf1mHitxW9hKwlyK5nx45mJbwTb0G
jaUOoaCzzMhknvEtIj6ju2N13/47Eo7OcJv15DxPEJM1Kv5f1q99q2rzkEcQc28xbQL5h0hT7f2x
tSRv4DniQOmWWynhU03KUPwIkcGbYbXtd5w0u9jVC2fx3hR103QWFS0pFsMaWnwY5R16ItHGRbht
E5nU5wmToBHzCfyfIik6DTxNcB3ipAi9rO3CsZlPI65C/qfkm722V/W3oaVQ6tB9QYOdWRm1h9fG
bfx15tXaBaYKcDam+raeJzKQajArQipQdLOCsrocgmi/oGDmXL9UGOsGCiO70tSIz0Epki7Y4pB4
f/+au6jLbzc/vwEcHAzIMMFukOynD8Za1cdrvqKRD+LAEZ7iT85h3d5nrcusj9dDr5+/SCTwOQlG
80kexafqVNO8jNwnaoWDSDXdI6FLl/Y9YR5/2b0kJ+Lf8wRs+zS035IrRU2mX6V/OKeQ8JXPl1V6
aoKw9EmZeju7bXykI/jNJwYS6YaYwvJpQLalms8rIKmXPiNmAGJ5qk9rhN4L1XNeoojm9DhcEofR
a3fxh+DI5JLwHJA0541rL0jQ593nQJ4Z4rXdXXzvtUs30bZwYstx0i9SKgMD+BDEc8k3yO52bi4V
i64WW7pb2lmzcZGqStVB+wcgbO2doEORJ9oAt3897Ewyrwj4si8jyoNC9ZOTNvhXCI6ssujXWY7q
UFJC469yTC4ANeiFjkmz78JBrM1J5+IGMuclt++DY8/Rlc5098c/vcSbbOuT7WG0H2PBhjQTZVr2
iSgGXBv/PH/mlVJRot3XXvpMhdXArXR+LAw1BUJe5Im0McjpW+sGyIHLdWXKpEznz5pR+Gti3bBj
8wTStcUld8RU8WYXBkBRbqaus0Jeu9LLQyIiZ6n4DOYuBdHE/kBf+Awrkk8UQgeUd7HHPbEwobYW
9jIexOphrlbcilYprlul97ie2Zh5sW7hkVOq1wIyHJoHgtGYaeM8Z/0c083wEM0hIb+/6RERmIui
jX3WoyZWArSIMFVTuZ7GQwWSlJ6ZVWsbUblDZasjdng9FLEavJStRYN13qmBF/5yEkkADdCS4SWA
JXMGRbFuR8JatQVheJjPnjr4xLDE8F7JwATP1eSZePXbQ+au3zA3bjUpvJFWDpJqdN7IJ4exkD22
7D27tfFo4weuRPWgwxHhEqYVXdNxXN+Ap9PXx1G7Bc5urHozXZdBOJdP7LAIClqA/IMzkQzp14Wg
QqoHW+XygIi+yJWDysj979PNg3JZDi+vrhs8D/nIFQTsQ5bZmkd4C80+T2sQ80+PmlEfJpgHdbUP
roQwTOeTkKm0+s5x3yeBMF+9ViMJNUh24vOLUAdiBOQMIWcZFo7ENnBxk7f7qeZmJLhTPpeQP72D
xxn9yB6J5PX2l7tAlCratRsFDnAx3CUcBqNHxal+pzjw/DQXaT1sKrfTiCCkovuZxrdNgiI9dcQq
S6JOYi7ac3kEFpMsxZmzUpenV9k1D2wR52wsAKICZA0VhRWRoqA+at0QEof0yNL3kwrFQSdVtNBU
sBJAjsTXQrRmeu62dYUHIpJtl01JZI/IJOZQ82b8xOMlKcSQSQ4vFipieqCBXp1GKbJ3IJQj5uvm
eISO7Or5OLY3M6kcXn7LP60xkLkjXP5KaMYJux+cjD0Gqwagyyg7xtEe8cNgi68x5UWWECZZ49si
tK3Ly+lbA/8wE+zNU3DcaH5vCgw3o+g3IuYViChkhTMBRFXA/GdxdLCvgeqho8LCxjkxWoZYuVov
MXF/Z5qXHVE1pX6g68e09D3ec/vJ1o0PpimEuRWvbnz9kdfWcX8BE9K+7Q//3aY2/CxG53hoOVL8
7qHW+EvVpASffctdqpy0PDmTvb+8qvdexV6MHFIHTmY+kksuehq0KrM8OZCDMvCb5r5ZGq+VWaex
WMNgzUeLhub+I5qCILUCspBTF9x2dgpT4bNVibltMPBPzWf7khaoqw0BGsXZBUybuw0Z5vK5cw93
2tZlu3b6UOhqraXgaxLLkcIIcBiQF8NAKWO8QTyqWlJ3xaJi4+s46CkWPtKd2q6NB4M3gMZ8nHRE
SKRLs2u7BD6KujKDmhvMHBwhNMui7CQ3+f/EfbMrai3ZdGCLBP63R3Ymr+eHG4trrbIv7L/Ra5P4
mOUx8azZXUFZmaLz9UUWn3ABooIo5Yz3de6gvl53/5GBSfxaj12CHIgyeUKuJsPnkCWag0tsp57D
JZ0bSNbuuSUVKI5WvKI16u8J+h7WBcGe/Pq94F9Tmpr78kCpEVejWp+lodbmdiLJH8YR+5IIO5qD
TLaQdt1h2ObWGCjizwCtbaaQN4BIJB0LpZjxV2ofBKyQqkV6XgZqKL7PRPJzmmZtomptC+Pi8Y/t
3KfAm24OuhCHOMoMNtRP91YsdYRq57mmKN+bpBX9VmvnarO1Qh6EyCieWGNbfyhLwp8rdHZE1ocO
8JBsLSmnLEf5QLdaiMM3sRr5/G40F+WIVdxR/0dU/t+J9IwynL3P2NsD7cIevtL7OTgFA8BomeS1
MfRXMgsIsxBtR7kdbFU8o48t4n8+MWM4GnOnovJ6kbdnlfQu6FlnvMS1dn2+859bdG5V/GV19LcL
JLFa+gHg7Fia04K6TaNiVC7dSMZie4ay8EZLVdNAAGgo92p9n4+wG3MfKr2Sky7J0nBB3Ga+x2lf
M8HwyTvgs5rDSVKda6ZqJ3oD+NDu+IhXmpy1HZF4jIa7t5x4V/vq8LV0tpEaZBsQKaMlTSHmYXD2
vlQnM73I/wy9Klq2yeZDu0XLgYHXlSQo4yf7UbgP2SQaj8X91bgPGWl+nhLvB7myYUBE97U827o2
bpi31L6gFXdr1xgMTqPAYRST2JdgxXM6Bem4yCavqeuEZ4fG2/iL/hmqetcxIKCjpGa9cwQ/E413
hs3hwqBAX1DQstS+rmZn5JEBqKZFCWwWkqGjnXK0TAGHY4iRFT36WdA7mQ0ZtLKb3HFVj3qXB+Jh
o8Vv3Y1lITEyujbh94iioCj23mfUmc+g+GmfUJc+Ltf6V4ZxEo9qPZTpWKgpequZSzND2TNcIFWt
LjHu1hH4EXqzk91R2mJtw5ivcp/w/Fk1envl26M4f6pLcCu7mXhen1HurgqEx0gUJYCmBNN8bsoQ
tjgJGJdo2cDEHL1OTAzUOWVSuWhk3NWGX110UkYj2sTlKMIRd5SSxHDy0Qn2GehGrBsndg8aRtQM
AaD7+srmeMtDGiRH0RHgEjoYge4vuIvZMIPKH30ymP7yzfuuClgKy0FIrWq05rS7xvyUj8bF8w4/
BRP0pNVOBAWTjZfJw9lDW2l444gtUfrhfweOPqbjEJyjzKysMrrfUX16KlCQH3yofcZYnzb6Mf+P
FZuyoS+tKGCStXFMvHAoPXCbZUZpvM5wmS6Uo8HnAmwF47u7l2h3mo33x1EpVjdndm62jXdvP6Fd
GlZFxNbIDAjVAch1CbyHW5a/StcjsdXGFGxTqPpxeLMFf+/BlfXD96E6JTMILq4l1YGLnw7GFTJL
VnAdJRd9SPs3gEL/tpS8SljO+doaf5OHeX7pyUSxNqt62WVIMCAgmCG/oXkSP5WfhgRuKU2RoAkq
9N1ken0rvuF2jUVdLs9OnOC0AQC3iNu2GPTC7XnC8MG66+nDuD5BcZNECa9NHJIR9NkBmbgXdjoa
wAIU9OI9M+YDl7onDXL8vPi37j6sh7aYKL+FcpdLRjA9818BpbD/y+mIuPA+JQEaTbEjKcW32k8B
DrTjzSEk7kzPy6lVb2UGxl2zcusUsHb76sLFLG/hSEX3MFmI92Rz3RgbtSGWQYsoWEssNVOfCML8
EM6AJkn9yrXqNoqL9t6Dxgk6GLTMSJ5fY4D6ouPlQLGLQg58Y++RVOFzXCMVcusUlyn/fUoxOhCq
0pwbrAQ3n06m/9QKho0AovP6+jFKFC5TtioBX2IkKdv/gIK9bDV4fSpGMmIPjNukGqsYCambuznH
YKNg6WHjrW7BWXtt5b45sXKlCa+7wRyGNEy/kQlWrI3Q0oW60cOA8Dv/uJWB9tG3nDRCObkdqdjo
91MetPXLoq4TQleKniTbvvjpPwxEIZUitTGTTovoFpMFFuMAnupa7lhapIdNEko3cThTNy/gvbst
SMZstZVC0a22QSoNavh6ukqVNwrMJD1tDvn2xeo/GU+tmVYBeZVgR5snLUAfkA4M28ZgH8jYgmbi
uk4Br1tLLJOP27ld5a11VVSQysUKe4+luz2EziwWlrjZIRnk2BUCfrT1qW9UBINmoEt5ErplNynX
ySQJy1iDvW1lKa5Q/qlF0RHLdLy5BrIMuVISTP78CDhNMIDhZnpjxBCdy1hDhgKhPIuS4xVjB3eK
hPLizCdx7rjnoT43lxdaumKD861uTJznoUJuUnJSSy0FCDG/lcUkGZPsFbpKgwWsT5hIQ11Sw5YU
PqPRFhojy18hfffUmhqArKO5/3er2tQ/qSKK1z3B+oOJCVUWETrPOIhS442Yq23f1CmQqdb9QrA/
+vKSvpmwsJicT1Sp5bdeluk0m1bZ8uJYgRltzL3kfuk0yaPMNfItbvziiK3AVrfFT7ofzYHyYhXI
XZaXi5yZHa/yVnvtYkITjKi0eghBcT/xtBJS66H1tu4R2Cn1xWyiRuk3cbnTIJVat3Q63vxDaUmX
FDva9zw6TVa7JDOPwLrELJTNW/jtYdBf3NgqPmby6c+r/m6Y0NlHTb924x9XrGjNrbMlL+c9ym5S
ZNLsm7GnBqQRgFLSZSkOjT3Xsa0jaRsccMw442A27HngioAgTrkKHAF8upgnPjwRmADviY3vx+oA
95xYWV0tj0AXbGRqMu/jmSE792oT2hBwxIm+7yihPFUWocz7rnXBmyVhW0Stmb0kVFgu0IeRL92s
zAtG0V8Ey1HqJrhNamscsKtivkdJ1XnNHuSrSobbixR5x7W/lr+y6SQK/+jI0li+yn6HedsclbLd
hGmp6oL3cVMvMVVbdtvSPZ11BE9wI+vNAGeMLlCT67+4D+4bi/mPvuNGcG55b2ZO7s5MA/L4lppP
36Aw+tlu9ghaDs57uYKpTsznoq4aUi0nAMacT3fIsIa/3hUCLIFcpWRSOAj4LQnQKQ9Om9Mz1ODx
7ap7kn7iD1RvzvmBAKEG8vg6ifKTEJvuSm3FwUNfMeT77QW49bdAi/Wa6vRqv8KIhvTVcUdF01jm
fu2lO+pxkVj9nG1AznDDyo2USla3iY++mHVEo0rfc8RQEuYeGg49PmlfAEF14ayf5w+G14k0ITry
QLWQA0p6zLfNfWffofbgepAr4h9jj8G7/sQqZlyTbhw9o5WBgQVNQA/0qb2U8nBrdgy9MxbkE2yR
G6KDsDGTBQXRvNQy+HLwduUeR/gmnIG4oe3DwbrB+IvyBLsdJTVWcU4e/lAj5NLqqt7iOGeDJiPM
UPh1jvCDGDEZ91FjO7E0e6Xfp2tREm/6v7TFyXXdtMcOCdxZ05Jd+TJLk/sXPZ+4C5MyKypRRARC
EpKD6gFUI9saR7wtsbzG/3FtGTjiZFiQXrOTMjqIhUbnM/Razzhx8KtB880QG/eKHSQTnBwVSY0/
SdMG5zCL7kYDUmTJ+QTQwPhpeQmBzHvxDRNZxWVDjnO5AqbIEpZWA6tWfdpxNKWx/OaZ1KB17dcC
e64rqQyffB3GyJhpsvqJD9f/CMSghNk3mHQ6zd8ji7lpBUUm8lpUzZbiI7mTExnf2WvE3ur0TSAJ
TiU0OhUU3HVVLlpiCRtbS78l+AMwDigyCxdWRlhCv8xn2G/UP/FKJYfw3CasNYhjSjAWUcdzGJoj
+ZpQIBR5cHacc/nFql2knJfFmAylMQ8N/1RgJL1VUVUkHN3wnthp3J6pVXNzBn7+HcJmZIS3EgKH
DOVpmUgohUDzH37Tgz2cYL0MW0l2oO7q5g7kvxOsp/wGtzBzOkyLg4a+5LW3NuEJ8rQfn/Q7FJCh
d71nU+LWX0cnFQobFZjmaxcOOVWG6SuujFamIpj1aQsjI5KZTJY32d4vr/CtrhiWs9qQrOebAbmu
rp5+poiGhBx6ZSRWVVJzJYf+z29AChbZZ2yoVxLDMSr5sBvKSkDtDLHWf4mlvfNDZrlaaopIB4of
Iet54JZwe6AG832JZxhoWoB+cBSoYV8K4seJ7DuN2xw90LCFOrayQxWZ3n4t/xELhwv86PUwZFGJ
4m3hGgJs71JWiHho13YHdMe/EHid2mslhBbT4jeQw/tFSU6sbTUxEjopJs5Wd/nNuRBdb432gAZG
7SWySNIgvRGX+SJh7SCHZcpM4l5qGuVt2nwTdVpoCBCSVfK3EczjGgEsIJbgGAI9J91pg3vz9ByG
W+pT8cD/miIdSJG9ZVhXrKpguP8aHkSZukxYe9XOfpkHmorYNjkUt55uGMAta47iBNk4RLS03jx0
XIpnOz/ZnXk/5+vFj1VKcih0NsJCOT0qy6z8GVOPNVSuVK5kFp1fJf301TkbNOy5QgUYF5Ond2iK
rRF3HptGCKiwYbZvnpCp0TzVgzRtX5MwJgCz1YGB/6FoiRIkQSSzdw5w0LcwgdeAQ+LQrmii8qJM
COEfcTjKZ49PuS+TyOrJyO2cqHjYax66nhqZTP51QIhlgRvE+ggWNH9CkO4KhqaictXuRfVVwlIF
wHV9NmGx4mk6Io6mpmDjX0BFgDx2UAIsJoWRtBAzZg4HKD8OqFN17K1bzznLjKfwS7O/KcnsOocr
w2sZsMCBh2GuDOeUyBDqsF9HaK96o3XXHcZUH5DCz92Z4R+YvhByz1G6uucabXji4V+NcLVbkNUf
oO6XJP+gbsxADmum7CNzeUiKwFKVzp/L1x3SaiOFwrhH6SvbCaXqtZRqar2yvAI3vg3zxhr/BV03
Gvu1vqUXlma7u3otCKN3LYkUk5m7goSTn/3ad9qnlHh2cHkaqgsbsuAdYuMncC6jgQ52GmwPH7kp
7qCnkAth9xp56f2CLc8ubOC1WZFasEK/DruZ1ZImQTzjtslPAPSKvcnQPEREVi+cQem6A3u0RYWj
KZRKlxKONZtlZrnvBPoTn3Ebifi8uHzV8gmU9dPvJdApANBvxL1fsmvtyr8nqeWXMovxS5bfl8as
DH/W1gZZzICAodB+UBWMo2F4up6fhcDTaSSDCRJQX31mw9w0O88PcPjlvB1aCQQndL66rgOsbrZT
5TaUi5U/vBTNlRqKuvVOqGGWUvk1hj5oGItbipo1tYKC0zdtdqFyWOVbxJQgIsXNwR6/9KxbY7uT
NMZhGExrVxKrvHA+If+L0bwVe18qlLcXHgKmDnrz2X1Ze/ieZU/hSfna1Hhnn6OkXCCYHORgcH84
y6aFpkdHJ/UeCSQ/3gy7+MSEzDFWGasT8CSmeRakX/gaGKWVHB4wjeI/1UMDRO+AyFMQt8gL9BuN
jDsRSZUXyh76B5YZLDB629tq8Ye2cmOoKb9rhpj06uwbQ+cV5EdpQD0E4FqooXb4BDETD03phX9D
pKWI9IrthPyEDIRJpWtLjY8xxFZQxIkB7BpWcGrWomT7G6t8BPm/t+24XatClU+eaN3rvlK73D14
zOm03oHNfLBQWJDKjjx9zDEpLrBHzp5Y+DY8wrG0TUDAYvhEYcGxaiuNWktRY1UStnFYFUZUCxRj
IecUD+jzuo9bMm2JuPji1NqxG/f2jvPeuFj5tEksUSP4WP7r0hJGz3kpAky7SYPwpo652+cH2HlO
mA0iPGYhZE2+wN6LSEi4kTHoEfrE9lbSvrKKOAE9L/KZyg3dQPwbPOZ+5c7qGZhTEJhACATOW1C4
mqCagxAGFL5LT7kTciNNv3ONOsHaBwFvHKB0B7MbIYpD0CygUaD9xDFADHx+HFzxdxJbwtSWZ6Nr
zOVGWrMWScyc+ZE5BswsPDB1xrP9+FAOTnliwJmVdmYrUHUdMudBYae2MlVGqf+WG2ixo2Jy1YSu
pVuFeZBDeqWL1rXVmz2QXusRdm0dEWen1Llox5qxtABKZGoplMYexLeajyHhZVOVofIktkZ2OPIH
wyBcCDLXy0Ys437jABXuoQgg/4HlYi8IXfuICXzKuu9euQ3S+FDbsSzHw0Uen9WFEOgmI5Qy11wS
aRu2VEZ2Ma/ixY6Onh7DLIf03FvW3S86ZlJUHvgmIf9CJhVbRxfDQ3kEfxKh14jb5bbRvI37wEqO
QdGtDwIvaEkDYgACojTigNlFwnFUVbnMMQs2r9sQ/OHT8m95a/j2fGNrPzTiQX+9Y8fSp3J928gH
sQEBndP2y1CLlYNNYG1dA4yNZKID5K2FcjXWLGPqVNEryRs/XzjddFZXXPh98L3ITh9prNewtA7T
xMPpMW1V9TQGjo4T5imZeeEX/C52civ4rJIpT3R0yxAlB0J1QpIyim6066/tiPBGyQLkTcBPWI1k
BA7XJbLlPQhfTjabzUFijjYFNsJ9kmCc+5Y3E0Jgayf7J5B1DZBF5ngBYWXzjm+uZ5PgLn3PO76J
S0J2Y+uLAhWNQZeknzPCkAiInbVTQ61enibhxQTArlakUenEgwKicdnZ467hgCP3qpUYC51ZBy2Q
dLY6XfNq1yUIhzWhEtgDWVwnc4j8bo5WhtKed/3velee9cUAjHsgbdeHCfZnmIrViW1D1394nqpb
gDDexTB3p1Q5l/Ucqurfru/NNFWBrJwfhsnkiUuJ9WcA6ZhmuH2Cf1hLJqRhC2t9MPZ8JD92lcrL
wAQdIptGT83R9OODammWXw4JD0VoN6FWUXeAgY+a1xMGdntHomK4bz+QZBdrNr6CHDFZnsYzH8fu
Ldn7wASFPtxcMkPCa38izSbuStW7FSoJ5c1LD20GkOiSGnHL6JCLK+1rxTvdTDzbjzQaVIcdcwyD
lApjcUoEzLazAAXqEGezaxyqobaviSFMT8sjfpzj4QnXtgtFVyH76D5bs1ERhD+oLCJ2PyhhPmif
I8o8hSxOcdkIjvA5W43evPVRQ8M1yEDjldypXCwX5br1Dr8jZkanNMlXrYQF7lbWw8gUM9bdpu+i
+o5YwiLKb98kB7rplNFpQpTHIStNJ0YB4FQ5LYLlGlppJ/tT9YZbX6FkcRfmmhuMpT7ReN3kdZIq
iXav5Fspb2UO//uP7iYAARjSm3t2t15k1WpH1SaHL+RyP5TAmrgZhjxyvoFQLxnRbNCF6gSh150H
WYbYKCJ0D8efVrLepZfwvQsJM10HPo5qgKEw5J6BboPnboZhOvAejOpBNFyNgdKCYPHXPQECoBKy
zqoAavs9DwnPtt85v7QaXBiteCfMb0XXBuITm5ThjC1y7mAl65iCZsDRePm/B7U8fMFiXirtXpVk
Gzr2URuerJwmmkDCRCs/uYheRRAhJZEhiM7HbohhEEV2t+YZl2vyzmq8KamQ9A4sQ45OlxmyUILS
3ajisVbpav3pokw41iCAYEoPxNeRrIoODPiAuViaBmpB8O0N7R1PZ+49ShicJyp4LiuEQ50om9Di
HFlNcSOBsfp1cM1mUSSaxx3EJ2Q1yXnp2PLCNvoZXhrGRtjdexAEVtAeTz0z8GAamRQDdjI29zmC
dSfpxP1H0jq3BI8yqOe6jr/EMqmQ8pK4rqgzPi9pd+EHPMYdm80TeojiIH9ShVBeQz4/xWu8fkqY
0PF0TDDR4CQ/xJ9S4joZ7rdoThvehgvjKyS0MPnS7UHmwW0b+HP/JnvF74KBc0pYazRPhOlC1X54
9L7TevertG/l/b5hFTtbc27RCJS/EKx2quZ/yhEAbqwSSTw9tsAChj9Hkre6QiAE07cDv4DpI3t+
fnFOa+8aFfvJIdW+HhhyQSwpGvC5bVBtk07ScgeZLEDdEV2ZupRkBHZzs1thxaL1nBvebB8Mr2qY
Cqscu1G0p/u49JYHmjyx+Zox0u5qtzWUllLUdvw0TijtqWCl9brbM61qKTqSBLpMskyx9A6PXvM3
xeN3+Cr1ayP4N1DjP0zyk2Db66tTVZdL61KuVnjNZXst8Z0EDJpiYKpZO2ofSJz24ciw/gV+uhJF
ngGxQ6jh5g1IluhulEX9ipET+yZ9XUFFRvbwuZ1gRSUwXGhTuGsw4d9jIaTjuiyGy+BiiES2+4SU
lp2QlTFGQIS/BkQWHr/MyT5RbZqET2voYARKuHuKvfyqUFXIWqxEHuwXRAUxUBxzdpPFrCYGk8Dq
mjQ/YBZ3NL7YQb7MiDtICGrNmD03d3eNxqmoePpZGeXpMQoq2TZrqcaSKOvpEtceAhyP3tyqGUi/
l1kCZKN5ac2zgzLddHX1xQuto7RBYKFiFZh1HLtrou8Tf/Zv9DTQPXjGkOBWkdaG830n/oLGs8nL
zojq7fIXm2Ce18AX2TepAj9pVmTqa7Bx9+mIR5jW5UWgpPC5+13Wlu1J7xrFsCWlNSePKfQBsCpv
inleaWE9jiejR2b4v6l52q3960d/bTLejYLNx8lyfSWkl8z69C8FPFdSxnE3b5GH+pG473lpPEGT
gDjGPl9VwYYkxa1QcNRuKK5knCQoSNZmnw3WcAx4AeQeRK2YElOvfWqWoSzxt11I7ZN8KrPlr/yn
ITihYzr8416Uzd2kP0DUKIkQa8eqLYJLW4XNBKK7SSE1/1Ko36dDKDcOPBPjRo2l0VzzpvnNhVr0
YoHLRwHBTwqY5xYrt5RHiHVJXHa5GZYLZTSB6QGlx0y6i7edPaB4dH/B25f1DLxr2vSCFcR9NADD
qhoRqkgzNBMusxHRrrVTsF6Giexkd0sOmL8LbbBP4rxPpmIlunTcyUtFQ+YXJChtTI9191Glwpsu
mbcc1JK7iv7rU8h/6iWn9DAkuCpEMv01fyei2tinOvynkM4hOOiY7QTNygFvK+M86LX9Yta3cAUk
95MC95OafmKPbGBm/wDKkeW3rDmaHiAnpzomLDS+zrojdwnThlndLhSXpZJG+BwDrYF+HdoVrQ5G
uW2nEhpS7s6jpnVDAirk1NrNZLKEhrqN3t3hlnrScegMqpFwKIhq44ov8cXB8gTgof8E6MilT0Jp
lvbkWy+8ttsBR4JUkoYRlN8aO3v0uN7NZXhvYgtX7MycCDkLaque9CtFBHKTa/5RyQdRQVQ9Yehh
qjIDm/JN5R6qE8Jusrhx2zIfUeiXuT2EdzTGhoplg2PDOkn79fT5SVB9lKxKf/B4Oa9fAlp9/fzl
zptEvVdRUYP0a4JxDhgzbKbMvKaKDq5xvJGwPclX1fz2DTtlg8LraQDlENxqcUK+FBMagg4NPkTQ
KaZlCOONvznKOlmpFLfFV8kdgFrvrhhEARzh3ZCMNcUbEZhesH3rFr3GLiHGAnd2TKDlEdKkHYdz
LoEK5s0StAyjkxz+ObeK+z4cEsblca4UKbFysA/X/jEI+wBUKM7CN3gfTgDhsiD4fxBt3L1t9whP
h/3/Raaj7oJSBng2l3dDVejw9ghi0ZijC37Tv/2Yt2aXs+JhY3qjcA+yKgEUCIwF5FmjXfelo9Ap
TGIvk8WBDNeKyLJ2ACw8jlyrG26zLJc8hf5oxsvUPuGMhxVnGKsHpy8jM3h8OUBhNpiSLJBRUqCB
Vf7rSsHfJRSZ7RL5zyQzPikhma85AO+x9Qw1oDDTX3MgaxuhOgnbLOUZD2z1m4W00M82r/k9UFMN
CXGKX+xYAZtrJWmCUtnZR8y2anMJi9Nk56aXtWNsmkcxJgRxnpQwamJ0XFaAt0kk3yldqs+2bhqM
P4V9n1FdAuFJFpvnkl3PnKJlWPhI5flbQ0Ra/vIFDHs2IZox4vLPA4xyZuQwD/nuYroRxu1n+6/J
tWJIVQP1UvhobRz0uCOwsf7fDQcdt2fzTfcYJHMSqiGbzgfqB3dQl2kdlC687GsFGeV7zkPTkDe0
/QJEfW3QNAXBgkaJEptsMXslAPD1KbCsjPB4DAGK5q04KlIaW7SXuX5UfUqs0qoTBIfNhj8CSWTt
MAYJQ577+NC4KY1/DiBL/QiqD9v7BvVs7p0TYfX2k6zRftGZlMgLQXb/CL3sTTvbtKf6i+frRrZ5
rtZL4Q+44ziQD0WPCrpZ9tcvmtWpeUJOPo+VlR6gML9Kc5WZIKUnse3gWcnxwhVAmHH201X92/Hq
QmKNsAMHcw7Q/0w6jBNvqxhz5HE4UZkyIbMJnvJljDrG+ZS65++Av1zUWTjg/vmwRFCG+8GnR7F5
je1+7laWCUIGSn+UP9flXLiI5TksXrBZbRxB5U4zWRsvkN/gUrm0eKQ8IqwEhKEZbda49hnnPe9r
SodNV/bU7WYRzxw+WvK72K577Ook6PZGppY3EBbd0D/BOkilYv6E1uslDn7qzkQg+KhdTLQX71wH
PQlLhQChoMgk8EPEXo8v/fcIqfKgRixCSFTKbqNyBTqvH8E3CjILKmgoOU8Vj0N84ciuciC4ghOJ
hqWGnh3Wh1Ph5Z1/0D3EbpLIiDSHE1sjsycOgrrWwGwwOQ7SFuo0bVuYCcYyZJ7kaXQfAQjAFPl9
h4hstHC+WwJn4We3hHeE7HjLaNYyOdk8iMgIsk6D79QR9WdI76gOvs/Cv7fnDlzT43IPKFoXREgm
4eQk0/vCLitmKdWZoaPuWQoJIeBvGQhpZTvwkornrP56LD23pD5LT/6npKkX2v2tlDHpL5aRo+zv
N4fAane7G/B3DSXC+Ow9c9STT94+mSBHCgCErCX16GOqsdPyFMhh9xV1/IvHJeEYmH/ZxqihQLNI
1vZq7JGeDt9kWxPOSj3OA57MjRUohg3ca4tjqaQ3/c6HRHzKIEfs+Nt0Qv8MpnAIV7JjpK9lfiPb
tF+UASG7fI6YzofRBDUI0ab0t0ti3LS96x058tYqYMsP1dLRWEMCLLhBIRrUBuSkCIS6KqGLzX4m
K4Aic9b5osNNp0J/T3F58nITijPM6fyVQ+sm81V7zLv49Q1zdVBThAJajB7+Xmx7YINj7y9er/ZI
xieWGXv7nmhG+S93ij3BH6DZO3L2e/JM+5dp9YvnrqdEX1F/TLIMFcHhr0ObhSm3EWcyKJK+UAAD
//VwRt7JfeV1mwsLIqEwXnOU+/5sbF8S/6aTu7+/Ql0YjsraA3akcR3h1EhOS9zxQDagJ4oHbrsV
g58AAok3u2J8TT9UiF6fniWXuaVL1n1z/2Gpi//hozApx4WgrG21If56p32HkRnR2xy9G6pOIcdb
bL9akuDtrQXTCtn+fS0WRlTEtTH/hLVTGe0lqa4pV9e5XjdCkzw1UcrFkOehBlwIbn7Jwd1cF+Sq
Hs9pQSJCpMwQuTM5rrr4KbYUVOgqAtd9IvvOKZBu2pz9Xl7/WfeZoDCrd/Jr3LQvFh6CGGDcvrh4
EEJ7MYfH0qzOWXi9O5A1U1qzJywl7CmeLsh54kNfy5HS6ddZY5F3TtsSltl0wy5ui5eGKmvFUlCX
sIlRy9gQvWT304J+20t6wa7OzV7TrV0UB5V7T7Eijj1gEsIA0VhkEqhQzE3O3HcdZLYtQC7Ppc7j
pRI8MgHOL9ky50CZ9J25wMRGutMUg/N0uYQ1g6VUjc81QBXD8qBcOQIf7tK46/cNakjKWc25dcoP
FpM0kHSoNqNU6HG1tsRWy2mdHwovcXJdFhT77U+fycNhnW80mtf0XyFyUY+LlD9IV+xZuRCg2kyt
kPIaYPQoxolZuizeLP1UoDzH+F3rpVpwbk1m7nB/n/L0dTC3UM4YWj0Guj2CRdEP4nAhMkgr2DuI
RoWjAIFycWvUePCdnB67FP7xufBy9bnyBPos6QDcuU/2tpaLSwugUGhqgjQIgY5ZDRRJoMvfKqum
uUWSNRffQzyWhzwtIKG6xxoJLr1hOQbVjM/zrZydGShcWA7ihvVzKeKsGdLTOXm7xE99Gi7ug3Va
A9Kx6sQrSI8rb2QkG2XUCu6LOjvUEIQY3vSmXLz22NEYQEbWjK7LREnVOLwSXgXR4HD0q6q9YlkW
vugr+Fr4pPh+NmmV8eGeHFs+/H7RnlatEw8dpF1VnRS8rL6+EQpeHjyyGVGZPtsaWPuV7JobtABt
KeOUiYSPw/q79gojOthxCgnB9sXZ1G6Z4bH9oOBZOHnx16eyRnREDagFUJ2oHFD68vbckY3WvZm2
jPDLP3wTRzZoKK+YbgSPvI2KsK9E5dUFb6XnCLPueLpofVEGKjBAcWz6uO8I5H2wGEr1rtvDd/ka
Y9tlVgnH12REsgy+X4/yicrA8igda1quKTPSxLCa/7uluALF64n1BBdXc8maOdTpoRCpv65DmBcB
lOgy7rU9DYIE5rd10Zr1Am7CY8lHUcnLJjtU4S4fu7l3BskZYAw6wsnvrpBpLcffv7Q44R9NiylU
mScfHFFDRgNsTWUOD7TCrfZOWmLi1eSB8WygFT9DuWZGQ2aSVJgHtgQh4b05RWVYiK48JV3Ue+VF
wAF6Ax3z/+s1m+rs5bPIG3DqyvEiv1BuzHYxixNnyToo5sQw0I+l1AmvuRUwlHhwomqVumwm+saS
c3npBfnTV/KJUiUmEy/xQ95wCfJd8/DdMtE/euQ9meDNwnIazIBp2/ksLS1AaLTKEh1q2URN2dwf
I3cMzLLPuKZJ39eg/SMoHMrWZ9PhaBFBVhkf1XAwGqRu/FPMFixOVjkYeBlzEcPp4FbTd4M4edAE
3M4JnM/Wj0sqWypwPGpQX6bPYBo+WO8GG7NmeS1+Hd1RWELNYIrNqbajw0fJGOzjUFXCINEzNCTp
W6HszWyGDdXcxGumQoswzS7doDZc5maaIfv9lxZAdwrPav1cKFys69s1RE/pgNinEfDEC5PNUw6i
z++5gaYrQnrxt6qKBiKPtuakXcko6oE19NVN9vjBZcZDddK2tDhn0z7xMRILnVhMEESeGlLvcYxy
jFWzGKR5O7lUceuMri0V4N/8X/u9oyc6aEPROlgo7MqYBUShKbrdIHYYYXuGYI7mHrrf7n4JgFEe
l8Y6DZn4A6phScBHIFVMND94Jq60qsyUIJQy9Ezva3pnUO4M0LMxIvrDPCAejRTY6ooTDWksg1C8
Ph4sTqn/5dlt5WoViTSPrppcyMU3/fKuXoH3Dt3RjlILHEv0pIQarQcPgPCanBS/x76HfcFs1gaM
G5dFP5qif67F7ayfIZjTwbMK/vCGz1Zc3qfZ4A2RC+yWTq9GPw8zvGlRkc/dyd6Hk8yCajMdP1TG
VW+9TMRhdxcnqRLYOHExx/PzLJNgqtx5VH2llf2dNY2hjZL9ly1vLbRrK/dMAY51xYhM4g1opxoy
iyj22TcQioETgA5Qd+HL6Zopplt4mjDs6pCDvFQhNDI9UkR4dmTjp2bCTXkIBsQONZRsPR7O6XuA
JNCWJMsLPmSjjAtHH6nYDDYZDUQ0GyBWUvfqQp90j4RGmt06IX6YoopzA0eOdEJfbNM4WnppxvZM
FuUJr6eshbFSNqTR+dXaubOKJ8RktU1BbQkDlHm8nEdh66MTwNgTzVNyFdehoau6KEk3ZwSrapdg
Lv2/JP0qUS5a5QIETg/lWpKodLPa4DB/PjBMoZUmCnzIaojKhnojzpGSA6AdvDUOO+G6MxS42Gtt
4J0QGSwwx8b6ZsjyXpTH661xIGwSMWygjJ47itB70WA3LUKE/232AA1jImLcVZgCjzHtyXv1M9Oa
bKUiXWxPLTDIuKsCcR5C56JNDXcGS6S41wWGGTPEgMfi1DoBAvh/R1qEVyoyAFg5Ic2zACKEy6V8
u3tv0fSjeIl4TBW8cWrCVFfFVrq7U9rrpWgnLenbx4FFYbFDRGTPmqEek4BHaK2Gvv0Cu8fBrh+o
Plst0c4zViL5s6ZJ0QFvidglNeEfkOC0i99ogQ5rOvjTx50DeKdGw/L75iyPJ9s4xnXrtH9j7Wzc
PYv+jwS/jLfeqS3VudsIAWvXbEVr0/ogn6/0jYtRkqDxs6mUjQfjxt0UsZkwWv/mCJ4XnO2S1Qrp
KAwp2sdROcA4Vs5gJip8QcYcDcMBmWGnFYuY8XZUmq80e6PZtKO2tzL0B4I5tN96O9COWZ6yJ3DO
XtgU2pB8V4Jjak1CtMycUHP7mL3ayPNiflqCb748ws/nDPUSd8Wdn3kwZMvQujTQQSYRl1RGQy4v
/GEdl2aNJiirgJm4knlioLt4WIxfNHZubSUGBSrMleJfvST3Dl8vT3rGQMVDlSq4BF8smI+x5VPX
T4UnbA6LS5nBdaixE3nKDLabIVDz0DyFmkAuq6D5fav3ilfdb+Mf2bcWvZFNDmnc2dn0Loa7Es3G
NX6HxeS9fIAkKvg7ruU2QQNJ/YkdmJJPSU1O09Cf7Y/aKdAJgksCQkr/JzP7tWhUtQT1bbMMCSE4
3jsnMmWGni0Zqi7+PghEm/PGYrGa/7u0Nl93BK9ty/uwOWAVVpSxWvuwUvs6VIMI6fu8VwanBE5S
LQ9BQosQVgtBoPB8LwFnc0vkQ4al2SSTkDN5AUmxMaWLh0rj/Xi1vx2pyENlNqAqlRGL+bQjQxIA
FPzcdLUD+oV8jiSpPcp4WnUsVwx1SFZDPL5z9FTEu6WdGp4E1g0Zd+JVvmhF5XTkKGJ8s3R6opje
Ef3PDohVgdTjNHmTqdgLQsMGQSPpQzPAROHwZR1MDFGQ5oKyb9QBvwISngaT2Pt83iXtUZCXUIGC
YVm4I9rY4ZtvtRn9Ma6ATMwwVH5Pscend9GvSAVR8rQ3+slYHZApoHO2VYxfUgO8OCfGLeygZ2Pm
A4TiV1DyT3pHigVggjANt5RMMuJaC8V7r22VUgPFl4lA2Rm2Ac4XgOjcM45OnB3YQXZXKowyTTZH
ZV+dghOcy4+lmmcsHZVQHeaiI3KZWmExuAWUaeFJUfK/beJim4M5W0CeKF9bTEG7nMNq4jxkCO44
hx3S9zheYIUPU7O7FE3ryzgzWhjjwRdo99/XvrZZb+ElR2ibqn8NYAmp7ooDI0r4AGhx2zLFScPb
oEUDN5ABsFbDsqfREIc6kYFyypfmXJN8s3oHl8roBq/c+KSc0iFtfUc9jyq4XbHJoaW/7oTyHPTl
GcHiim0Ftru/pnY99IEoadq13dEJobngZ2oZm96PKBhOhFAUBXPdNTY103db0D33beMGKIN+oD05
qeFjQ7vCdZMfpe0MZuG+Qilc9IM1ctMzOES58WFNUxWdHcZJxAZP3QZAaaUWZdGbe2fQf4CzzJug
2BAWfNhirX4reJ3eWv80LMr7y2CRfCQCLpD3sHbH3zOQBeZ8jAGw3FV6xOexeQM5tBcQFYA28lr5
8NPT149C9d9VIQfGbWjnAG7aVJry7zgPXH1xFzhuJNSU1dqk1nPZtSdVtEd6/+U7ssn2IwPhNigp
vxUY/80mIXtsgQgHWBmd3CRQDBUBGI4JliWbufWYlK8aLgnUqyPQevyNJGlExjFVbgCveX1qX1qv
vlSfNZoUP+urhDWX/Khs4OfJjU/aOaaRVzakB66Y0lnYbObEUye4FsdMGpgToNjokd3WrtuL3rnW
P7KoWV+LXcuRVBJQuR88cKNnEbjzwB20XevmHgtUPrYRi/VIRb/8Sb6GRC9H70+7sHDZ3q9G6/4U
2y5IqEDyW9tNjJCllNks/WnXnc978JPSxUi0zl8WzYuA3bSNE7fcacOa/B2zBxVSKJzE7ip05xiO
O93lyAOzpofUik5meUoNjxm6lr6DnwoR2swSEJUOg6QPA2LSSSLwC9TCIqXgLRP0xeCs3MvEpD5o
Zxpe487EM+DBqfuPJJvHhsyWrWh7wDqhqsVuvUIT1dUfsw8QboACjrQASclZZ3+5AvOzCALhyWbM
NjdIEXHFrZbNjogRHL4IKw88AYBrFGVifxsEddLrKP+zQF0s8aiL0YUrJu7tOCcWzLQDlpvNbCtB
PbqLN4raEq9MWGFQvyu7WFQs+uK7T/jMEo/BeWKjQrU0XVK55cWSsV/Djz6XO8RL7IOOxuZd1Y8M
fBq4j/tpojBPxp2Vh9lD/fpDjjtW9jeShCzubWVSeWgjcTyDQ43bpx9Bh+eNz5XuIIHb/Ju/IFB3
EXDzYJ4WEd9ZJF2xKMBoAb8Fi0VWo/FWWnWwljTauirBhERHKHVlUDisCCjYR1rkZj09A0+BlvOJ
2cpN0Iaj/tpbnUlu2QH7PzsjTfUbb2dYQIP30g6ZIm1zVKhjQJJk/dXIAZYMeRpQGxxqcuyQX4V0
MNfhYFlZetgNZXfPAxdJ88U8sz8iuQHKRFu9yCnHtnMS53LEW+ZGYuzQ9rLGJyDYpFvuN79twESt
IkTr3CFahAKT0KKAwsNsFwG7qh0W77UhvMXe1VOm69AvLBU75X/0N75ZVO3bPFoQFMJh56GDkVHG
azIKGPtcWrt+q/52h1LU0YuTb3Im08adOIcMJfDz1kuOhg1sEgiMW4MwmH7yuD/RIfsLd99AedL2
ly6RIxym7bm7a0sDULj7bxqTOyFcX6eem10VhCU3iN7uXl30WZt6cYMxZ5KacTAs+WVDrIePF105
3QZmJ5++JwbO0IXfiT8vPXn6aNbn+fzvtwakOUqPNsCu2j14805JOEk21h2NlMKh70U1ENV54g1N
UXRCvPciF1QgvMlTiolcVlcfSmi67C6SBarXjXcboiXbLIemZD5V69Hfa+Lc2fEG0O7Hvx7prmzp
I4b24Yz3tJq12ymkEbfGEOJcEJBi+Zsvw8yCYfXzSQ9hSU8qxY7L/QqIfoUFRVgk+tBfX1qZcTBt
ZJIrf47C5+0zTgJbh8WJkSOBLFt7ckUhthVzJxrgrYqaEh83cjTQTRN18GsLUMBm2V9KSL+UyEVE
chGkilszbAgqvYf6aiEsAU/cTQFsLVSly8IR7Z2H6S2RnD9WUkIjeWmSwjaNRgttS9qnAcqVyh41
E6mdY+ur9H/PGVu3krjjMmtHwnyYij1l0A1zMdj21EgwF1E+bWSBgJal5eGCRl9N9uEuKEDXxfo/
S8vDMHk1xic9Of2zB0XQyBUtKkIOj04OLvNUoXUIHk9YSiYZFtzh+mnoKrOPzQUBkRgYLpXLVxhk
VqFXPvC8PL3e4LDhgtYgwHBu97WSiHYT8Md/behQ7K3DiRg94wcfTXbNL7gAkUPCEZ0x3bpk6DVW
6DrvQxiQkNIJK9htos9qphobTnGUV3Z49uqtRkQ0VP5EFcwp4htbv8ZsL3Y6xhKcBc0JGI5vvy+k
Rz+jBjjKFB/AcVmE8Yso7vbY7bNz33igtSJK1blpZzG+T6kCrI5/R8S35snVSf+T5edBVUEWwOiy
Q+wDDHv7xzCSIxK/KSvq+3bY8AORw8zd8ZidKAsC1h9hOHONpLvRaFM2BKXzhUANljcvnE64RmWF
NHA234Ff120v827KUSQDyzBjn0LUXMOr/LcBnmi/o9Gh8yPzHkpdCrOexYT9dLE+boY/D5OWVvoY
D8HSmMoxalL4q6+uC9o+sNQ7Z+bi3P5feFChy0WiLILUY2Iei/gdZ6W8ujODRGTznorLsJ/oJjM2
rDIca85UmsO+hriBTcBxgRm/H5MJ/IoPQf7Jhc1RbJTNk2DEo74azkA8+YAgxqsWp5DtV/xR6cT3
g6PbjBndAHcLRSpqEZ+FPENmCyboQswl8+CxFpq6INfAUEKNzRPFcIZQNxlDfI2RuhCA4V/brAq3
+1XMi3janNxwlS6/rFL2yVaC/ih9XU82hgtnwviym6p58bLJToR8TLfwn3Jn38JAyxG6sWa771Af
XqggLhjZHqwvgQUq+cKgwF9yXc9keg77H5w/hPPPvoWiPr7auGKd/1desyYFE1uVvCSjVciG9tLu
kjJjnRaJ0wW3nx4nGKCLS2tWKAIF2RHKsquy/6det4FkK0IddDpDJZbdkaxgm941hBlf5b3bp/0l
D3RejEdrpoCK9fiRLolIMQSeG6tvMnBKcBsfhGe3MSM/wnfV/C1SwQ3aXhZ09MczDb+L7eNtNBiO
p0xjU0M7ViNcJZULUYsC/cD5bkU/YTDFkDmpVWoUf7ZkRiqCzF/+9iE/DJ8BAjfudVxNEJs7gEPt
RR8V03bxnzqhhK3Bw9ezGj3xraauhTQPeDz0pd5j5h1DhO08mK+oa88EcQylLmNaDLOElm7EJGx7
C7y1as13PoRUTrxegw4deY/gXi55ZtsHXNB8oicJ8mD9A0FtuacG4MAWo+hnHiejWmVnoeNdaT/b
8D4ONZLwqaM26PZPyl36fu29R2+k7gnYm/04sfUtTMZg78qGDZfkut3+96sJwhfmQ4usq7hdjY+R
RQSkn1pIxTqJXSa/T5TI9nkGudbtbm9qZi487lxYOx4NyaYwO1F1ey+plvgRYj5iS+7RxTVyDR6g
K2fNMymoVoJzHwBFeaerErIzrjJEHceZZO0scQhIXmahr/1ld/xUZI9D//oAxwE3H/oo0HhRRyLZ
Cr/e/xjaHU8CMnKQBGTDQnmeC6LBD+UDnrBBbqCtLYsFsy1qgPCnnfAdCFJ1dWEowkvOu6N0sJVO
Utcnr84RjU4iLyJJayoxbFbWFevsvYP1r5S61vKo2mZzT151O6X+/9K+lDYpEJwhNlWTz0zdetvI
AcXkqMzu2iy1xrWGS9pw3x1G9YDVu3yhHSRb6bh5MGbirHLUxBnZq233Cr93z8jJBqD3gLGuL7h3
mULHq3sMZHkdThZkM7hZEOlVUoYwghwkikuuOCxPvHI/4Dj46M/H3rPC+RpZ77HHjSDIiICnkCL4
YQtuB255/906gDPfhKkfVJSUnV5eCLl5RvIY3qsw+Cc+XcPRxXIGbnXP11o0KLwd5NbElUGN3czq
OUR8AbE7kxiuYA9loBvMdqCjgUqmQfCxfcdSzOQXj53AV924isXBQdW5oEcCXI/eIXiOf5uYamtJ
uS5mTFyvZGYC6WjVWUP19cqUwfp8picyjzGOvv3hDjT6oV0dXstgHMeBB5lYoNrj/GyDaROAB04t
0XUyZyF0rjjydrocpVejyjxOYDA8xwBn4hTCTAJhQyV0KljOslN+TMIRLMRCJITeOYMI/RqNjMYH
w82y6U5t2nprwLrW0UnDErpt7VGyWTHIKtNVgnzNr6ZkCXjsd+h8qw0FGjMAiPZ1pDwu74bHaL/m
7rPmQe1xlwWU2Hm7G6u7G0VEyHwhdcud8Uyv5fBq017HzGxCU3dShcxtbO/52jGNsaQxnl38wi4t
2xXU1m9K4+8Uz5I/3xDq6ULezRo2STavZE7THrS3t4n/dfWSvALcSQO6JVdHn5mTWXThecjsDTBo
zh3bx7tV1E6CGLqR4kM1xFXsJ2k9OSV9/zRG54F+TU69OA9r+rbAmXa1Wz9uaKgzcFJbMS+OmIJs
WAqcSqSQFTUmEXG4cjSrIYFMKcRAf1f2qb+T19DDNexYCb3vrO61H0FnaI4LIolESgKk69J/dHbC
y8wDWW+qJ7SdqhSj93hZ2NZX2tmYCk2DCrBmvqgmVqw8q6ktqKxefJnMq6nRXRPI0CqpRuNNfRxl
O4+iLWy8SpQFfAYeXVvEF3ao0djmK0UF/0kc+8KQrY4rxjA7GQkIogN8vATCdmeBjBVjM8y3IqP4
f/GjV/yKQ923ku35A6GvHo7ZXaYtC+bJJAGdBQ/1jLeKfS1OuiIC2rCIHc2dBCys43nrX+xddbN9
26/2te7Haw3cL8KVovQu8iTXlMMPBVWRGn5x8LgEDLK/cLwqXFBF5kNpz3hVEjQYaEoTMKDBz03h
G27z8rjbFFTxm4MRPdhutS2g9j2oVEb+xHEe8d+YWYxcS43/VRG/YxhXxeCnyetX+ij2uX+dc8HY
H4GtRWgtSfFP6H6ZrnMirKsJ0r4kqJnUaX3zTBVKt2u2ALQZFwd2MA7soMNG9RLlz4qnbpuVen5X
NySFtkMPMmxkMtsb9gVHkhAj+ywcagwBUO5xZiZQVqryx7yh+qFXgCGKW6wukNHUqGn9bVLesrlJ
OfYfLl9nLVjAm9TX8IKx8K9bTMeDn2M43QYc0aAOCgzkIIPMb5s4ipxs9mg140GrJaxH+sRK5zjO
Ok4vo3oWZzDHhmhp/ItbZfWWDDji/XC+LKVPHoI14ncanjS6q0WW33XHiYex5H3cqpYDyF2/nr+I
jja5DSICnNd2nHIH5uCh7j6WYp3xQ+pHEejGO79oL3zXekm7O+QMngsgiEWwO+uhz3LyMjDPJRBh
b1aR9vUmn1r0+y3Za/pm5cpCnmnP5dlQBfmIScy//0WuYvLepEyzaXCaKAWUmEKFKuO79WC4bSvm
MLtfyjtOltZHq6cd5aP5i61F9Uj7x6LUZOQ/ZVjJQj/w0h0Xc0nmXf2KFpnu/zK3s7tVmWGiqiv8
vq1IAzUxw70hNMAV0kCPaBF/iLZlFXohKbXcAZrKkkypAtIJOmCu7yUSqzrAG353eqanaBPTIKom
usu5G2vtqunoHUloxo8TeKCM/yxyx2zkx4RuBZpENKUis2d/1ObccOGERvu5DegiABk0XdQZw/G/
Uh8OsRYpNTOrGcW/Cbt1lDWvPq/TL7YT82WFh8nq+Itfi+qxMzUhS6Jze/Aa5DU947HDA+0KQwRI
NE8mbudRfkUICIYjiGdxsI62goG4Plu/3bnEZfV/mIw4MeIwKu80vpm+gCwMJfPWc88hdlqQ3vyD
6OVbh0HUyGVYuCpeygw7tzrq73mmtiHD85ZRaLLPGBt3yi6VFWpFpm4jgaJetVXHmOkB6K0IPGb0
NuOV7UWIpDzTQAXKc620M6qQ+FgLU2ak91LyIvVOAoOreFymxwxR8O1UTrkvHSTOJhXeVneOkiJ+
AjB/Pekn7xwYJJ/akFkueoi/o2/8GgSTewJpYy9GynjRMyK9307dC3CONvsx2fTipdMSzs4Kq0gb
8PCS7eIlfuudFDmP8j7Ah4YG8MEbscb3BcUrjal0GEpdSm7JU2YfaD6pxpwjJ/Ir3fZgl4LDQfb2
REGy0KAt37xngP6T/wZhOModSR+58qCTjenuCrfxwtx4HzrxMhwdXDlB8tswxtGiNjWevSE0t/lV
IDdy4ikmD1x/YaUtxxKYjWYtfK3it/a8p/QFXWSlgFNCFcHEGJ/vXZUrGBOxzi9Gom21/ZczENc+
hOpMdr54DP/ROZa9i3pNosJHilvMI0XBMmUpO3wIzGQT0tiEJWHV0Yrc+RpH+iYZrrmVlDSYeLhg
wQvIfnBWWhvZeXmUVbHQ7HfFZNc9u1vCL7aUCq70NkcwGpkOgMfRnXfQFLIKCYiZ/ld66peVS7+3
yJtTCwvZ5iqf0JQUR4tkrK/JiADLX8DZou49wTyGKayYVKPrM1/Dd9ZsXh0SGCNGNpsyLi/k6FI2
GTh+QwWT9+hnQjCKi3Fx6bDC0UUweTbvvofEdCdDcGVkMXX1nTXGw8qwMBDb82meOudYkRuJg9Hc
+xJA62af01nEt5vwApIDXU0aj1r02TKOpTHGofK3jAn8RHj734P9E/3nZtEihKo/6uqWXL0hM4zJ
lld4VesH5MSLJy5UVfyqdhYFPjzMOCSHA7LQXoo9zH2BF1KqFIWGtH6DNPKEWWe8/Dc7dAGnaHh7
9kxQYuAMucLkc4lggojxWk3tw4ciFWYSE4nDEhrqCrmdP9H166zs7eTBUh1eXZnVU7Gfp8SBNoJ/
28nAKMHvsqIQd/rFuE8iVmtz+eoXsycnrUJSARCnLpdCqtcpyhzUHJGuXcQNzbc47+SOdltrWNBQ
8UrbwUPY+mhvQvgiP1VkUZP9Bnvg/EVieJCru/huttzFhG7hom+WfkhlkfbCGZYSVTLaUOOF5ubv
w5ZVJ5dRanTf6cN77Utw77BP1/faQFyIFwk7lzghcKbpxKmh3HHG8fV4aLf+79utbEa/bN9HB4S1
caqcRPLhHIziS0RrfQOp19rZaxUbSg6+u+JMMZI2VY6F5mF7QFzMyO5EC5jW0yxKeAu0ZQDJhdJB
07ZWhfVNPX8iUJRqxq667nNBTBs/7r0H8vgEUc/Jj2+FVFawcWqRlwQS0mqEZfI3K9dcGSmjsebL
fezmI6P21BjXih/FKkFH8Zmil003vZuKXB8qDl1XmVYFvN5Wxmqd6jCRCtc8rzdz7U/vwsfH5Xk5
K4YiCVvNzoGfFXSkyDAgeM9JYhIwMiAzyiI9IRwr7GHVEEMmNNHQkfj21w9WZz6WSzQ7hFD3RWZF
1DpRZjgP1VykXtxBfNXDA1fMIflMwo+CzOV5y0vD6f5IksTgjPyEzkTcJBXkwix/xEGg8fPZJCm0
9Q07FNRZAHBPC9MdVVPPnSSnSGFjy4HKQr88nnX2yNaBp2xmMY7zRa+TrEG3/TaN8IK4m1GLhgdo
puvQBfZ7iCbhDJ80HRNeXuHRAjGYesb+AKZV8nZtJ3+dlW6/Z+09gWuQ39SU32onV3Y1KDk+QjAq
/5By5WNHVI5nxh7FLLJQm24sQKOOqXix785eNDo375vMDOl0O+QZFl/4bq/hPCG4v5i1pkp+yu6M
NhqzdHY3EFOoJwRlXJo+J27v62UMh3dFEkTlzo59tYVrRCL2+w/oekTi1ucQJKzCxT2qud6pS5Kh
lWmvRUzbRWBVzm2F3yH7f2jBNw4Knr8nm9Z2SW5rwIVnmhg3BnWx5MxA2d85cAMVVC2S1Ns0MNdM
u3vLKI6WDNhqPJMrN/m/1TTEtJoZgukuUSMY1jArmQ+6E8a3yZHo/hfkPTqUeIZ+zL14c69CsY7S
5d4K5LnaIKPoB23SzYdDmcfnGkoKoSRaNN1tiJT+E/QkBb1Oh/nDReheDTsi1ltwBjdmSD4rRd5+
MEHiD9AQlLrCidtoap0xnBr2SsxpYPJu22nOVNWF4UjQI2Kv3ybx9g5kceZ11PQQhwZ7OnZI8UBW
VcEj5cfJFk7t/1Bl8wFoz7J4xb2wMV0OyN1vNixfN0Do65lh9LczuVqK8ekjdOUFPU4I5yACZdwi
NiCJGcreeY6BGzT07gAQXVDzf6MMbhujuRVP8Vq4+DeNTTlTBDtEBVOGB/0lxWM6fbij+h3Z33jx
M1Iy7NqpRkHu7ab+9ZmK5eWxUyD7dte3FKL/PJbpS/vBfGtHkRJwrLghaJOFe36NJ8m8gf+UwLoh
fD5FlPxWRJBNDGSACzpzPGFHQKhzlvRXpZJhiT71a/PsgRFK9wUsj2MsG2B1OKmo2vsKLmBfUzzc
N/A6Y0WwXCEMcdZUXu7O9Bkj/xUyb3wtcvAyDogeOIcbM1IWZJkLYSxvCHmfzP0KHJRlTy8EPxMG
dakvXd71eDldHfHZbzAyPj7CzWAipV/YLOZsKoE9cx7Nbinxj/+nyEc1PCbfjg57lJaSberhwAG8
RUkVBQdpK3UBrQ2EIUJVS7td402BiFpNZLFusmPtzi/BTOG8CWHWD3mDaCW9a2F1mthlwDzpTkBp
TiadDleFlLtNacoN1r2uxGf2F8CBGCJ41OnJvAbYeVYbfr5cANbnmeUcR6plwwvGPhJFSECyc46y
GURVeKctB7qB2k3xInxxvJD4ZXSdrahzWkEAG7dq017vtyjp0Jnr6onux0+kryxANqFbhfXN+d9o
mzuQzej4CyH2Zc5ev8fKf7ivoci42BULvYtDuk8ryIwvo+8QsOTF/037QhJcXe/UfRdVufO00TUl
OyCkpewFqs4THp0JGk/RJ+EZouUhmXMYdwXRlz40YrSrUQ5l3VlwiJGslqwXsRfP2vFcKuaEoVL1
VnR6Cs7ykSmUucLwveD8rhRP00mPLjVuw2Hd+exeT/1prmtnxI/67qKTAWZVlYP979jtWbBopmR6
p/fLJCE2IYeXHlZ3CHoVzfLH5FBaJvbCqTSPgutgTwpdl754bJZijJ3dA8eND47oWS3yBvrzKTi1
zYI1t8AbBlYkAK8wvhHWR+YZ7sbkpMwLd5ZWW2XhYu1mxVw8OJVgXSulBQ+o/22VCl7rNYKXixTh
dv0a/o9gFErYq9oOtIddzPv1mnsT0wrMpJ0gpF/CzO2m/wO2xZbmsJe2btwclvVlYkjiwTgBv9/t
zzNnJlA5L1MHc3i7Y0HHsNaL/zKDb0pjdiGQethRLwNB2eUlv3J5erBcCl9wlCGf/A6skt9gL1mQ
EE7qnCfCtxDJ3mW6mA3GksM7HztX5mjIIsoR7TK1aMuJkJ0uUY15BI7eIDBE1u0v2uu+GP+rr0C/
gxUSxIGERDTjKhFzXwB67wZSkub6O2Rg1v/juw/AHBOmzSBVmn2lW5ZPq+xeTNQQnQDuo4hhx7Zy
oyuyrsvnqdLwp4jpw6vRq2ha+1hT0kvTLIXXg1F/Shx/rnLaGQ2pTgusk1bnrR3OHrp43MC1LkNj
KxrHMem2E+OlQ8a2cR7twGoHDc8B7/xWg8MwTfi5LLiwR9ZTZqj1OsbOCz4qoSb9hPhKUA36a/b3
ceMne4YBouAGR2CpGFGAC/c29COrkLUZZQQA+YWwR6xa6RfZ9ln8njWRab7cQqhBFzCawg0nA5Uu
ZGqgTFGmkaVZzVzX1+LXnE2fQLuvk1wg8wHnRiBfzd6R76glG0ETW9eavPBTlzdJhFlGllawgliW
iCRBfGSG9TFv/IKfZJsNV8iiTG0TCWwtDkg7iBbjwOz5XxMCSPzNDuyMCTsbKpQ0RYlH89mRaTKB
9yq7GELbiuhxjtw0tdHMzh+RG1qB0qDd8+9469PsYLjxn844g3kjXHWKdjvqtz3ySaLV71MGrqK+
PlbWeNJYRKOm6UDEsmwjvAO84ILPW02yxaPIa60q8GlChcEGpq3JtJ+x3f3IKmDqQEqPJeFECRpx
NSsx+qsvdLIwAtZ17iKCHlA8yr8YsC/zPn996xQOUsj4EcpCef1Jp0PqdUJgpKLVBnAGrtPDEK0H
Q0kB76Z8+p/x+cZYqSi48ZkpXKElFaJeNnD1j8bbbWgjuhTBp/QNk4yljLyJjsM/6ApAvbiq2h2U
uqP5cBWrKKqM07UxNDFl8m2ZTLBTOwTg6uT4cJ9n8+EOULRJehCd3Kpra2I4Y+rwmlhLQogsLMUY
V5ci50/f47fOT9/2A+kb+xIDqExA+JC0pe7c+Uy2FiIo07++crxPDM7dLPdcZ+3SyGgiKsKcerQm
UEbtBizLVqeUrp3pubz5udShskVlnAnKO1b/28qS2NCGfFWsVFgv4C/KtG31eQpvUFIbesYrnXSI
zeRrFo0bnswOeP5D8pMnRJynuVFxi8NYnufvgnzKT3qYb5/Wemh6o7LS9imfVbR6Kv+mlQcRqRaa
dnz5jx1kU1WcspzUHZZYiCNZV5uiaxDfS0o2gh1n9YON1a6X8eH9oGPuSsuTSmn3+jViuQ/rSDV1
44o7H7v4OmwJ4pJhHMyL14iGJ2NNPW4pW3Iw5jOGkAUwV+pQu8FUPEd1UNP1BPGajVVD5ryZAFN4
RJwIZFG8HJd2UOePD5r8GGJLy9pNXxxRSFE86jm5bLQ9AowZKUhrJExygLciJecViiSPxMoXfLj/
TKdh+Z7zn6fP6wa79GqOC530f1owEUcDsxWnISQNxewzkd6Y0Xl2ut3nzq76Unz30zSDO84gXzES
l0NMeotv9Ofi7jJJy4FCHYOeRJrm/Pfw6w8QCl8dBKHgh+4v+72lUtbYA+daaHeUxS/W9Z4UHe8B
OhXikAL/0UfWGj6kuCvVXNSVrKUJEKqmHuws+sRDUdWBjkCs9v77Sw4W6nGCz+bK52spYsCGSKJr
PsyK7u/DbcrD1tiF4Nndlbwct19EUXdrqWHlgdNQJ0abNPj3v1KchoDY6ohxupImoFYxQBfgjAN4
s05VYy5DGCaJxQjPiOUwhQkaLaU3kfSrdtI+rQC5HBUUp6VzM8Au8sLorCWaspE8bF7ZSnFAS2QJ
MEfBF/Nx15hUVeWamTLHigPkfxW8QgMUhqsxA1U1doiGA0bPjdfsrnGxfhDN0l21FJWGoKrN0JhQ
UHXcO39z6dQgq98JaNmKObAzw9vB2uzMcQUBjygNaJiMpFoAB2R6u6SRnu95XOfVq8dJQMG/APOZ
CKnyfqBXQ3BZHmGnXq7rtFDROLfgG8o//M/8+Mqtvsh9erdiKwhUU4/hQbER+pO2OF6WFrhVOKop
M1ORr9Gb7ZIh2ewLP0NT+ewksWCFfSnStPR2Pn8ihpHPAxsNjON0zSnvcE/62v+leIMH34BPb0IL
E4vXmke178zr3Jczh224xvf+rt4JtRMiIKzyrHsdvaCngw+6mSwuQzv8RgnpiFa1gd/xErZQDSzg
a+fCdr+/W25x9+xaYkMt4k0kLI+f6mHrqoT7WoHPnongW3EZlZiTo26oJrP+ClQSKAxq5zDAXETk
fTwlj2DwwSuMDtU6TsJ32SS2Iwh/LrUJDPx731dorAmF0Bsw2mCPzWfF93/7xLM6k36BwZrHRVC/
WkhLoctNCq001ZMLPD1o9dDlxffFkfiIEcyBMgQKSQRil0zBEpPFp23ZFx2xAowBEp5zvuWIcxlJ
fNQjcYVfarpdq0XgOsruHH7BzvJQPmL1O668KvMIRUgpYtEMMdm5vN5kW6pWBpYo5pXYWgHGRps5
/10UeQAzs8Si7tGnVjsdkqhXjRgysAe1oOv5/2NmWOLfQzosaY++370gDqwVgzTUUg+rY+BhJSeG
IKf7/C8V3z2VkAj9T+tX7JbQwqoGg33Q+asps1PL3SMblaj0Fb1PNp6Nc9NVSi+q0XlfVIKe5Yf9
coqh3TAy4XLksa7w8vhisD7ahCURwE6ipj7JTioSRHgc4xrY8c8waw8vWvGuHtVs/zjIhVsziGyA
R0tZyURCOhIvRp9MUNLu8/TzD90YPhiQ4rocmvBKcjFDztWz0+5nDzPdNQ5YBUUVkzn1Q6LYuxSL
X8GgBDJWEBIbetUN8Nvq3N4qvv5GlBXw2H1g4aLxZfV+sNkG8ydW5VPV3MteqUSCZ3EWb5R/PfkJ
WR1Wrw3aQb3F3SwGbO4ivfLawvxySx8KOlN0VEG8/K8NNtLeW+SkJQL1sZTfLanETqh5peQ7Ebdg
usWhxYXOjmjalx6i6vcsVgoJi3f0iUXS1VT3V/qhIxB+M0PGxAqJ3siTO3CkmnYyIKBAV7d+ZgO8
6DXgqI2/7wxxBPbpla/XpMufBpgVNTYAKff6ZVOgw5ZWJd7/0cKQpR56sNXJKnPf1Eie7OYgMmXO
VTYZ2PZUuM3MQxsDc8uVcI6z9EtRbaSU0EgXWFJTc7ULXcbo/c15Bc7JBisWK95lEzHIpMQwvFih
sbRwYjBoCUU/eTXli5eiXqgNrB5/vWHZUPurAqmAYZk3VxOAsOdpA6gk52KzZ4sV4m+/lIQ2XRdw
5Dzoq4SWlmgVeRz3urehMekzEK1vEgomo5r48PZ2UD7UU0frg+I8b+mTHvjSXUwOpd7Ytos5hUtg
UpNf3JxuDsZz8gf25aBcxQcV549Ru1UflOTHETDQOnMfs7lunv0ssfSV4TiFPAzEPKwtgkppzmKe
x3d9LlQtTz5uzwPApOBCaFCcQh7mtthwD2kV3lebMCvLwWH6JFVkVJx3QOdsI0eKaJEahJBtVt/o
JmvcC5do2mQ9bXwav60ZKy0j4NrzpnIQz+grzWpysG3V3K+6h/D3gsYtJEZIk+GKmV+6Sgxz+GaQ
WS1HKoRsK/WTorfildXuj7iY1i8DMuDtz0Mt0PnzZf6UC+D4KUXtiWETvvwCW2YxaxvgNYdY1zcY
HfhG2/QQrF+aeYfU/Xk31FA0SDoD9Q2TnB+m/pAHFWEdcP0k4m7ELhnWrnYuYlC2bS1VmrQqeUTt
Ui8kEzNNqdSEHTW+sIexH9UvaSe0VkNcBxldF0x/KHtNv569XADROgTPIDCPxV1DjctTp8crL+MT
QSx6X2CsxJLWBmn6JLuT853lBX27XNALgvN6yfyPvZY+v9HZDOoLycCnCsD4WPckY1iNxab3mn48
BGy75QtCravd7s4Hg7XwPBRJyfDPvU4GU8EsGz9YdMnBv4ycYJKehQPmTPd/TpcWisET2FA8s+vI
xzf7w6AUgis+B7smJPxZyC9XCWyrkt+B2TnnKwK+PPOectma6d76CobUEdldbDffVJWlyqXmqcwF
hAHcfwUp67vAu7gRCr9DLut221kBb1D1yN4UcdWCo+9D39zhAJMQ4hw7wosVhd7vgU82ADHGeCsN
PmsgdXO0lkxFW7kQjWCU4unVYuhNffzU+Opg19vKY/f2cRon2kTL1/ACMlKgqx4YVuq6nnMZPYjh
d4ypJ+HUaCzID41vyE8Ixddl8dpHPbcigOhYo3cdlyLo4HnJzn0N6n2TWdFhF/8dSP1o7cjR3y72
8sjowJ9QAMJBlpGJlKea8TFesWcg0GSruiLvPExbdNA+E2BVnGA3NprDwLaQuQl1Xcbh0uYiyMQM
XTeUqsYqO0ko4RHUnsuCyxlCGyFdUkFB/RfgPKGAYuQjpiKV+/KPQ38o8rV8mG0fPe2vweeVIu7v
91mXCs6qJKSdXheynH1zIhDG64L1IC2bFj0s4HTJvV3RGJrfRL43KXrhzDIpqWfqleHQaK+tmJ43
fTfyVTWCWFactcPHAO2LORRy3NqWWO7GnTaBbr9sTCt9GfsnlH34mNWyKzY6wVav+R7CC2VY6F9H
lSL5srBc+oKwVwF4se2eAf1+9hud9+VV1GqgfZD/EuPq7Ik8UWI7L3hYriHkWhpgW6LyLWH3d11V
sVIQdgKs/mULBCjcZr2HU+9+PtBM0XcnJA2shAxp/App5UV8wmmoDZhdzeMPswmv3gf3UEam790W
S2iIHOHDOurswdssJAsuAuOhNdTsCN3reQ5QL6g7kBDs9WbvQS6j2nN1HHBI0JciLe9etLS/E735
AGsjmkne/z4KF5R75YAyeaLaBA4I6RAZBcRhahag22+foM1YvwQpDvOQ2A1jSbzJwAhV+iKQZeoI
wGztF62jFxWY+1TpLgbf5x3rq9dKT+Av24NfQrX6oE4nAqQVrDLhRb8IzfLhyGVjShHpclb7Vpib
zeADoMLRJNieC43vQc1COKYtIkrOjEUNhFWyduCpDIRXEYKTN54fcaXquDJr/hEwm1SuGZAHfkHK
Eqkabvm3Nde3k3vCcQuFgw9DEFTYYRj3lrTT/ioReUHEMv6OiEEjYrYSgcRfy64mcC+LdphEFhZx
pR2RWnptq9j8QHHB4u6NjgNqMVFzWbN833IL6W71jja+j6Cj6dW/cU4ZzppKTbvkYEGPBlK5uFXc
0c/c4rID+DSA5sOZPP+KPcMjV8NUfDG3uNwSan+6j9IpmL/VRt4uO83IuWY9hKP6o0RSkyE9tLpm
/ZcFx3vTc0kuPVQV21LgEH/k/ZDojgEfk18iH3q98+/Ol1OANLXCW39J1hJHCE7uU//y6VSLm9Xb
dsKfs67l5WCTk3FlVsdwaPHENeeApKTnbOFYDhJqDeUJsa6SpOAIai4swspfjkPYIw98fmtC4vQT
ZLKZ5+3KH9AMRndHwqiyj4xqKm8UHVCFYku4PyojDjJtgn/quvyFD/LcKdybc43Ze2peDXqmRzwn
TPFV7nYudaOp9RkOiv3hEh6KmLc+qcjlFYBPR6gQ8TePCzZDgOA/Im+pQwRajhtqZXp8p/QYLZ8K
mn2/FiJmi5+GeNMtqjJBMHPJS4waL9rNY/prj3HkPDuciyloZ9nhG7BPtKakUrSe6e2Vvil3+sCa
jUs5AVLI2qcOVhIX/qOFq171il5vw8flRezCQye+giaHA2whcZWWCOy1uJQBnAPwAzlA/BsezgVp
Aoyc0Wl9bxVAfPRWuVz0PFbmxPEzSp6j2kNt5i+78Ovlj3AJGPu5ZNW+cPpiFYwZzv570MqHskxb
HwitozrtBqd6KqwSvpvsrQq8erUMkRnFibVGPSvmgWJLla1/RLVfsyaIGSS5aonBAeA7RXC96iwY
1WIC8WkF31h6uOGJKM8n6MVAt1gzh9cD1zRwynycDJNIBhPxH8X4uNFr33Jcule1f8xUtgfdlJHU
3paPl9ohiUWAe60DAca06c1TQPew61TB5MqgT6JxBK8cVaVK8tok19uEQE9XWMoNpcfQtx0E3FCa
fE9g/1cWyMy54SX0jtKMIFPiVG7mkL1klHny3nmr3MOis0ojhtTxfqL328ibIwxCsRo8DNJtqqYQ
pJDA8JZ9hucCmEZQv8/MsrSNOqcOICBqAtwVq9aQ9UwaW4q/JfaX490xdsdn58W5kAXnEaIx6706
ilxaeF0Gyzjize+FhQx2HDgqM6XH7oruRTVUBr5i1XXDuxx60yyGfVM0II1cmdQzr4BafFXN1j4S
GHJrEGZUuU60/GGYm+JnLCwPZkwxsuP8RjTDm35dG/ANP1j2Ij244bgj4twMupjXBzhrjVf3ma0w
90PNqqdR6CGG3tZBqPmQlqzVJRK+aX8XMlTFks+5mD0pygguW2D1rGCofLHC0vISBUeTLPSa2MkQ
TR1Yy7Z5M97hfGEOhk8uIhni8TtAT2YhoYxt3Zp+xjCSjVX7b0vu17bp8Jt1eqvdUaPzXNPYSjt4
dJiuvJTnsKHdvJJkQiscdz98XEUdc45jyOmb4zgQM26W5hSPJeVwLnq9JcMGRC3NUcAo+/DP8vD4
H2IWjb4BxabnFhx2B9cqwUkHdGyoUFHB0pthEmn71WbipEsYgLUu1WKhM8lSaueDtJ2fj/l+uCFX
XSaYe2u/minfU8NgDNbuC8K8BO8/bBCgqvOpBuPlfXyeTJku5iy9KRxvS4cmaigA1N9WeF2PIuL1
2cx6vI4MPOfFx8MxgI/KA+lP4/FBXFnpx8kOAu4WVmEM8CL7kZjW7N+Hnz51WHMr39ZrDJWueQEM
/Bqu3jRZ8ZWlZ0MajwPYpJIlu//GDi1+YynqxCVzEvbgPyhGlSlczqPUq/gPZXe28d5CfY3kg4kL
puWKvQ5LB9z/anGHXTxZUN5GRM9yfuDjz1fx52qrLml/SE8gOygaDlkcT6Pgljks87yKv6zQm8qt
H8YpcqKnI/md7Vud0rLapMTvaIHhoLoKAUEHh6H8DKecDEL8tm3lE3lTUeX36KjKeIZah0ppN9Y0
VZbRsCQ0dm5SbbzLHHWFCjQpCjFszvWpKc6vnpHi5ZtvZclZyZWuEIfn6qRTwYWD6mRUjBUZndft
Qm5PyfAP0P5tn2ho+mVZqCoCGV45nhr2sMhV9PXdR7SQCqdw14eCLLRMIctzjp3fmtzdH+0M7LOB
6CDl2Gvffm3mz2z1Llmgn6yn95JU5IPAlvfGBj1AEFifC/bYT6MacRccnksUKgE0eyi8dyXt+XF1
91goqwtrNMfPEh3j+tNXtu3/36bT9cYPzf3ko95RU1hrJXod+hIOFsDN74W8nBCSv1wPyTuH6p4/
g89NpqugjAfx5tw/FSeT4uyHRYDGUdVqKApzUF8xOMHTZ+Uds9vzYeEhvOysB3P6m6Lx6b5eMSpI
SF+6ne3ro26ifwXDzQNuAgF+QMQ+lN4xZiBAuUU87ESZKCPqIjX2PZirjUZ8ZxWDRBVghS+jgUYz
YO5Cb1FZFCefd4+eUzwTGaBu6n+DyHzodGQo8kVprQuXn8ioAgWV7TcsWJor56kaLyLMqB1S7szt
S411p/rHY487jnVVBlmNpNm3H/5CNuSnx1TDEr1dYNmIdRM00jLPSFbn4CFv1RJQMv+PaB3a+Y6z
zDTjbYKq6wkCtuVBAr3jxnRR5z1Zom2u84C7enHF+9qhxnuwnR+DZtG5Gu73VoojN0rGBQdWRXEB
/Das6AN9Mb+QxE8m7aoR7nWmAz4kluHBxMNyYvbQ/wBW6DMYLkq6JqXevNQX5tMc2+7Vq+9t4Scv
77/sM1hQWqjXF/K0oEYw07Q1IA5AZdajymqsKQ+DobAGLgkwO3MRVtcJPZ9OKZB1UJpxQQ3uEuAR
3RCz87sV2Q5DmmAWnjhUOEbHddKwmKTE+ow/3RnugdHFLVD1rP6sOHB62s8eJHEJj6uITeaVWaRB
cMWMSmt4uonsRaAE0vu5LWXvz7CrvkC2kvWNDv43CDWHOG08ewJ6LIjXy0JS8Jawnwnfgy/McC/B
lXSi7ZeqZ2BRZNY6mbuG58lK9eCGgKAW+4iqwUNcrZH/blEECs8zvSRLHjbKOkVuPSOENCYtnU98
CduMHgxmbHzVjG22JDJVUUZ+Vvq4OcoQ6A6IrJy/i79gVIw0Y+Mq/OpItFZNOJ0hhMBNzU8rMh0l
Z8KY96pyKDoKFJWFKe7Gye66jqefpNHaKJjL9oWwTol/88nY7PGMOTgO/IHNIxC8YsjGxrO6JTL5
gFiM5aCtey5yAcU6m5mK/tThSGYfzAB989S12bxVHlif3xYeeGrxIvG0j7nGYP+S0BgwMZ+FFL0j
gjByRgSXJzs/hVHAhWFk5gcJ8w9y0iSgRn70mGTU5p8FZM8Wa/D0lC7VfJ8pAafKlvMLxcw9Kav4
QqWMeWJNlmmB1TsmuEbhVi3lx8XgLUv3QJ0+7/6SV1RAHyyClC+kvwPJDGaQX7QIQ7RNRJs4Ot4t
rl0k/8tsGU3UcFRWz7X0TMX79U8yUOEZMW3uV2LV2TVBybTtj3JDOx6SYUjM6RZS8mKs1K/Mxfg8
X94WuYzj4SlI3m/tpYtfvRJ/DqweC+Q8CO/PPVTeOe3dtfmvA9XyaWPPi05EBtT89yiYiRFV0pMb
VqQM2lzmXGUdOm1RY1U1gdxmEex77n3slodANVhjeuGoTLHsTM5rqgXYxFVUI8jhcEcu1lWN8WXE
0MynyTNYphDYVQOSHla8Br8b67KI4o5/+P2cj1xwuTjPn3CgEWZ3WBXWit77dVj8Xt7jhPZM2nTL
clqBNebC86Wu49r6YR8MJEBjKzASicMNKsaXnVjMY8wPe6i4SFNT8CzBzFwLrpW0EVhu5zArxU2e
TORjsN9Wy/v8XimfrhcHdaYuRfX69a9KN5SiTU6BFi1YqrPHXj3A8Rf4tBzrpLW/+pl+bRiSEJk6
8JEEbYH0i8LdYVaxSh5gdtKLPvzcTfwybMN88VUnK9oiugRXzHDywMaQ13f6zkxjK3443ShKV+Sz
L+rw8l+uvxb+k/ra2t/57lOSxEx+AyUh+EWIHNdx42GCLwXr28aSeTLC21zFaMbufGfDYYlGT2ux
yhAst5C6mXz6e693oxTnhPLx2aQoY20Ea68wzlG+PEXUEX7mvx/PdDD6iEjhf72BEVV7ui77cBeD
zKAdADOQXkbyB5OkYse3nFgdZe/eH5tA+2Sr6F6ZNATdBu43xudBNGnnvpFro9H7Hj5eVaFT4/9N
VQILRCy1AMpB5RLM0dSFILZpXkTTbvIqtPrfDtkcCLTzPoAEtNtMKswbUb9riRPQADSLFJJiRNMl
SuZY+v+W+tQb2xJvaHbPSFR3xXrCvlq2b42kFFoHajS+tIbjV21g7QBGUoMVEwHLn/xQMFWASs2P
Mes4Ltkc7Y0+LVb+1yRdK/A4LbIAVOsIWAYr3ztspcakKtqZjhXs6f1kXav/Luan8ErNGx9FvG7x
OtYJQ9Oj6blRxOGGRGr6OK1LOIq5ph7m2iv65mocaD1XTXTPl9O5dSoYPM8hA4uzjQTkXH91c7dl
OnvbD106w5CgZrKWunopifB7Cb9liOadPCmRBWUOxxrJb09R64pJd4KuSUueXuLVfJ/AD1Xcnhj/
Zai6wz7aN8vAaSPy0om6GT63A8hlv9RejLWrZ6UZwpi9EXpWHIwlsBLUKP5wjMEcF9E/AlLUclkA
9KHdEj2LYI8sxohKWsHtutMhVXfojcyDKrgpDMQXx8V+EM7V7cV5HSsnD1GYXeQnaY8EBx7xG6QF
NmvppFYwCVOxigreRtxbO4E5UT572Qy/Nu5l6VLN002J33DlaAQ0krqdoLo93nJ4ejVBXZmeiM2/
x8C81tqYHBv0g0RQr8ugPiNcWg7kFXB27S/PrZtiJXv1pfhj49wAciMz1dGFOeeHvE7+xsij52kW
MH2t7rxrylWu0ZTFmoDPeabg6FVwbxYeF36drAVgikHa0YJLcQg3SkEe1YaEjp4JXR5PnoCfBEEX
zu6AXwehmK4c1+aMCWH4ObDESzidY+m7Nk/sx/obTielRYnEgl4N3kbq/0IT4VN3h6YMOo3hthwu
gD6C3uI4+ELEU6JDstmI4VyMlmntwr3UVdOuBhMdGU2mlRUvrU5/ZbSFlw2xeLKcsVmLHSdBB1GB
JhvJVKJLUTisn0lES8oOpzXQhPqjTmxGupA112tgpYthJ4fcFm6yonJDNnrRKo5vWszcMaOOaac9
y6viVBCZvy/rZG8PE5CnZkUSFnG4yIVqcKJcXo5nULeeQLBvfZTkVv8ahXPC/cL1NRXAOak+t5JX
Eu4TfwUmh8+ZgQE60hZrrnhzpJr3INToJpaua+fqGsnbcx6GaSZ4Q26NH63luy4lYYTZlLFsHgkU
VRawMIFqaHuH3mePlR5R4OnT2CASwgCPUEHA7VCSw1PorFFuqII+TaMHsxDPsSp5OAe1+skbpYbx
sUfchrLnXygJPA7vl3NanlEv6luvkOZl9Gi/+oDVtnzktWjs8+oqMk6N/6d1cdmO4MPPreZJyHg3
jTq8wMhJqNQW1BqTV4Xyds0QMwlkTGRrt9WFbLltz1mHPuZe43ZlFoVZnM99f8JGlYmsVZzrchjX
UNsjltAcO7XCoZZBYfc8vju+SeAxC9MVCKmlB9h6M/gNeZfe9G+yIwwTP0lltq8LB7UYhRq+bL5S
gKw05PTKCvbag7LXd27PIue08m6TmLtisj+WRxtpPsAYgIGbFsGgRd7UlZd2aQmsczPKCc3qi9DJ
TPvGDkaHC/RN9TOv4mH7loo77s+92jSTmGJLsNWc8ARfZs0fvRWCzmSYPz7DS0dfPdeL5RtrIE49
0MZaVA+qqspdfHrrbVGR/105VSHYXZeE+YG4D4nqy+eBD8eya3Znf0YtFawjbxfDFcNHTae5uTiz
YBkMaJnO8Ddb3Hu5YGW0Cx3M0pplS++tFoSGkU1f3euhFaO1rhVXh21DJmB4pNDLOfC7pv+lxiK8
qkqFLxj8om+K4sH1bScd335MvlLw1A2aRmLOmSd8h50QgJBgVVbJKQXIWiRhEXP7rFt6bf+HfNiz
U4UVT8Jn91tUNYiPMgR3n1UXC+9e0OVmobV4il7HHBEBMY/ewdlw3xydZldwHmjEWAMcZ58nstyO
kwT21vg6kBMPcaa4MTKdeGdXYxjq6BhFjlyPV29JMAN5Q1x2G3NIGVu7XeCOZNb0R1Aw45KAZyFo
f56vH3slxoQ+1SyRq7fSWFU3RgNi0q9hfSVr53pn8oRYEHVT5g08vRV1+qRcndzdJAhA6Ihvncpd
zpf9i+PKGnMYPX+wnPlPL9HDZXPYbPbxey1LAYpnaGbUdAOPvTrqhJttFO+xlMfR4gEpEoaLb7dQ
3+VEroqhfTaV2pSlJxBsJjlVt4l1aUGV//psXZG9JCfQHeJsznoxnKL+LBkPhYYFMUHAtMN+ux9W
ahrKZpL13fy4PKxcRBgs0SpicVyFeOC2h1p5nfnIDyBZ3fF4bK1Mj727QGyYSbhKPMR/P+LdXZh+
7Jjmc9Ka2xWVWLqPx/w5ERp38Npj7EGqeUY+VKH3rGVdityE7logen0A1MA4fp1GlR2KT3kLOguU
hrGiMFzYxM4QtEjX+uHr2USYnPc2wpLOtUb1JqE8kw2GA4v0q9rhmZf+rFNczBENumk+s2mgy4J4
Ei3sPGwML+EsJZ/063rbR79AnAgnCwiUx2xmoYhZu4IOAc4rwJBoj3nDetlNXr6nEMQTu46HufnR
MWA0KKET7wMnSQG2Jn/drOe4GuJcS3cTE4Et4CUh8W0uPy3z1B06oi9nL+LJy4VwKaET0Kt0qxfH
/CXBUzftDmHUF3tTPTn9P2tWJazRYHP8CqMNHN4nv2Di6rJ2n4MFwtQLA20sdA+HOLd5rQN+NgqT
A8NZ07dm4tUBRpnBfhXyqN82rwRmOU/glqlcrFc4wSM//lTZ/x4ZsTdqtT7pGzAg7iNzcdcOElj2
roivA1MYRyfhxjBxosZ57j7PotiEDFwDn8ZPoPgK9GzKvOWixvus4ekRGdp3gxtVuXRM7qbygmBu
fic3eHoYTBaM+Uoa+WP74XHpSJP8ZAM26k2qHTrVA41tnaGyc3IluPGC+xyFy2skQ1mgX04a0IIC
8hWw/WQoqyfQIka+DeDzlnA87BzQbPMNyUo2qsIqCue1v6owTQ0wFVKjYukazlwHX0iRSiniEcmE
2IiNrjVVK9iLBu2aRqgOFq6iRY+maun9cInkpUpMsDDWeOejC8HqTJfNpd6VAlRRXldZcH+LRf2l
qXZjJSc6k3bfjpNA5X28g1oZ/Yow+ZxWD8TnjVsoyYqWPZynkMKo60a7fvunlM8QngxFadI3xbjJ
5/CIRldLMGxGL32Tz9PdC7DyZJeEvmSzjNvWKHPK/oFj3+egGu2M+sqmiQXlmKBAPsCPe3GwRtXc
z3Aza8fq/taLwtWgFEQ6OiYfGu93E4kVC/FDHME8LWYloZcYc03VRdoA4PC4+4iVZnS5xNnPtJFB
SxIndzr4LLJtFor2JgErwkboab+opgwI01hQoKlimrJNlMrZfQJQiJmCUt9i4fT1Y2tQEKBMJWS/
WWXm1tC2zOmXgD0/HjBzstYr6vnc8GWNsOC8XbJ4pJC6nmBVwFXfK1tXtSGfjsUTZGaBQxvNpIrP
UMbEB3qofqnsJAtenl1Ccn2JOnLbICkbZtU2JtDtlzcRnSisOwmndZZNl28k5JQo56gzQWh8LUap
iqqF4T9eHLWvvybLqlC0/XuVkI+CUADC7vF1Uh4wCIQgm9xZnwkAmGTTT0iiCekgcVaA7LdI3eTg
XrdYAImgM1YmzrpPzzz0nVIzz1t/nC8FR8PMqk4kzYbWYJ9xNQFProStvOG8n5o/LVFIza8A6Fvg
zXOMLDE1NRLkdPrrzrJu1fe/FUQ5Y7YYgol5r/pTYT23f3I9zcL2IjPYyLw8sRh79tCvabmev+d0
9Rt4t0Gw3aRGyq4uJAkML0wG5ORoMzTVG6tdYhAYqWDnNC4NlWn4/Cc1nbQWHKMvx2HbmOzwpM/0
+LW7M0p2ga0nnlLGtRfJLuoYFX483Ft92ssk4ThgIEs0NF+UsPlV9Kkw4Y7pJ7M5g/a23nM7gLL0
NqM/ABktStRjUOfuT9yBF5KlUHM8ZOiUO3Q8mG7UZzmcxz4mx1UC7+GUu+B/K4U1qcIa3rNLjO3l
VV8xO4OXs6HRQdLXs+8enmihgjW2CZeY4WC526o4OXWLY72DAFwIgD2f84bFyoaJriK3oz1n/RlS
IMqZ/7qws6FRXhB58QeluYi8YzxN5K/mCVC9PGWsf4MhUgfh6N+8Hkx5bQDo0KAZlmSc0C1aeMyB
tZU8V0+tu9jIHbOXAC80UUsJHkU1ZtTAgUvma2EeoZkzTIAa+4zGckx2KpNIyfKEcYYCKVN5uuQy
2Kg1m47TRe6V9/3Up5zmZhjqeUtqJuSLvE8++mEE4bdeRQtbV8mozX0qsBSXkkb5PMqUA7YhxOpk
ytlaKH5zO3MjdinlGfJ3nDjlM/mxi3SsU2pAwyYVS8PLU6PYmOvO0QtaLBKGkRHZdBH3CjlBs5Yr
eLqN3DzEkQWxwsiNiK5/y+OqiWe23tQoXbNWQ0JhhWqnwLyXp3ep7gI9oFtxXh4kIUJ3FKmndx69
8BGtb13LMLATryHDOUfz/LlQ67J6RL084TN0VG/5tCWv2uA0geSme+dztVi1kB6Yiq83z0+UKhpx
g03fLu4lCGT+6Iu/SpEep4cBYN0D/Vdm4v03CaWdwfaVczWYzIt/6gDd5RqH5cky1Q6Za2KGkoy2
adT66iB3XdDoapcNmsynzuwCmJrXpdkW8WDg6dZG5Q3qFTqSgoOWPkNhHCAYWQMu1TGrQyXXiU8D
YCPMHAjIApCDWTOZ2s00JXnM4zlFhanzN070JNYUiYcSWya/lcbe3jZ7zqNMk4fBLsFiYqgVRoPO
1d8WGYuRidHWpGM1DIJTgEnpRntcgn6WJfImuWGloL1MP6L2LWHu+l3qTFmoDx/4wCgSjZK5KqdV
KlkJWb+vrCLC2RDI7i9AUZ6VkBul1T1J+GX6EvibrvSbAKRfXPyjmzwNR1FFxbACY7Yr3vvp0Z5B
O8qH/iKzW0wBM94hTONSSvBWY/J47LrXLZR9KgXPmVX4zrmhfk2zY5ey3XDlSnJQPu9Mwp6MAvIs
hNir5MhfVpzu9G3NEnykOgyl2FMZJ21fxafs0PUU/+kUzKCq+aoNTF5GxvqU6fASq4BJzird1oLX
GOzP7ENtD84TJ34wY2ToCQzTrhW6YzmhOogx5LhGBx4q1ej7Qw9JWrF0lovS5iakfZG1swLuV2/G
AxuahWsHkMBchujBrRqWeu6CEQfzBPkEGulc5sOfI1UvOQRPxEmNi2hPSJU75FARq4cSm1c3ivB2
b40aANF1atsYysxze//wjFD1wTznMbAiiUPhgsq0bfWqgHLYIW7JgLwne/iZBwrY82avAP4bxs33
pl0ZVCYCRWuQi0B+Ga3yJW+SmY/FO4F8DNoMA0FIp2nSqVTh5G+c+N/7NRN04B260aAWXSCQ8kFb
7AwLKU92I+x4Xp652RUkecoj20YHE4uKsA+bwPKMmcu1BpqPb8TtXUrRSHuDy1bmIOIusB3HHslN
ya8xdFCdiFcWSkizcMUdd5Ma4EVnFSidFylMb8a34FV6WJxNT/Hrnsq77YkFLQ0PUwK56B6+9eqN
DwbsmJj1rDHSGV3EOLtCiQBGveiYjruvoi8+oNFDtZTFL5ZQzedqwu/QXqtttNXwAo4KOsDR7+Ge
ywuHG6mCyJU7m8E4w+3R2gBS4ui8AYPCw2Ptuliqt3URgFfO4R0YQ3XRmw0vnmn2/gMucRV8HiCu
RGNFjUzKL/YflrriLiOn2qoKEdTqihmp39ac80FxusBcsncFlXB9UI/uhl9flAZJnsbsKyJq+alF
iSslesDaxF3uwXoa24+Vny2qz2gHJK5FAOzMWQC7JSIXUzCmJ4KZotpM22izJhAXU8KstQxHzybs
RqeXV2RVxS2bosCxwcV1iQdAw1/y0yhjtSIPxuZRa+ajuZXgD2gIHrrh394NMV09KIcEib3p+K9H
XlS1n8aiK7nuGODSugTspTSgZ3L7FYTS+zVc2zx76GDny+uGW/nlwQeptlHiPemqnGMnWQai98vM
T3jN3LPerypEfI98Lh2wqm7O6Bq12IcVXIUCHzUjC7/YwtOyE83a7bvZ7zzeH+n+YY/+gkx/drPC
nmZ1yhdFlVImkiTF50peS6imI4Js246gb1qZAC/ItO2eFJIQNNavFDrYD21oTYlY8HMRWiQL7+fO
7i7cjWKErCSctv5t4HJN1341MA5juS7/papS7sa8Rn917Ud3W6iuWe2iq39h3bZSJ0oTY0j9ax8i
7e0ozizyRVFEHxye7GfXB2VxCdjZZnWwPZUBVXWC7waBDzmnvab65mUcddmAtTGQR696NTT7sk5d
42rOfwa9gGvL1fmAywn21P0KfP42pHWUisW1H2JDeT0lGu8IXWVj1eUCAIYUi7mtPsNlSCO8zZCd
yGqF2bUSZAyi+P61JXJZAThAKLnDvM1rSvUag+tLr3lUA2bPKzsSqdZSXMq75T57GTecxL/8Q9I5
8TnfxJCNE13Xjr49pamr5nFn/YDgbAaVQPa40WcPrqyrn25woPO2nF8Ecz8xA6XflZt9GwZrl8dV
uLO2MyyUGcLYVY1YD09Rel1VbBDPTdBdu5VJexzrZMuVdDe29qWt53BkMY/pDYpJU+ZKOMAxihBR
pLPUm9ms8SBUYquADkJ9blgXr9VU6i439eIKEj1I3aKiYH43s05fVTB4KG1/d+paA9Jn/n6tB6bN
Go5pfxPT0JCpkl7arkGH5vhtgkn8D7i07EVx022pnEiYKLkHCZKJQjxEGAN/jYLYg51qnLi+SRXx
VAQxE7zRkXGHW5YGnwwoLGHtE5gfVJq4llzNDBp4NTLT5TSszzPvLiEdHYe3OzCSgtdD54jhE8H6
INHbxARRgFykKVBtYEwbujf0NffmG/zQ9geX709m0XcSOyKiB7ia/K5HmF+ANgHOjhw3VSi2C2FR
B87vGenKCL3yw+UiaFqXxCSsivMRm70uBQoZFuWXc4Y5egsr0wO9CvRFESkNDDQ+cGzA5Ea3wJyy
ltQAXSpzEhSZSU87Lx9iUq0w8tKkEHIQgNPxoyQKf92l4K1XwA9WUO9shOWF8u9gCLv7/NOhm69T
eYsOXMl6/uTn9ReNsx4gtA7uauV3CLCNqIil2+NdWENraROqYayGUlkUThl0r+fPH+rgusflIrK8
rua+AgiAEGGSU6RJRV7PvYZXCaw/6TEe+PsVFUZIVmoh+X0XbdXXgvFhegD+mFu+J076ACwjMqdX
qFcPCTvDy+RMaiO0Djldx3D6jIMa3bCYWRpVU4HYEpm6Wss8+ZRBBXBRKIAnQtKDlOPP6VxiRE/J
JbNdhh7GoXbrxbJxIhX/d5D52oI8zoxCyM44IeGGMSHXKeQ9Uz8gHTm8fK9/TP0WVuCDZFor1xjp
dxidzXQwRS8e/z/bIzZIunC3n/IYWzlwl7HaNYzIIM2GB7jt+RGdhT+7wcSGuiB/zQUWNPSM7YWp
JnAOe1mCn5JrGD/sMJMSRNYCU1gQAW7n864fboyE/sIIu4a74rXRzDekx5lv35sBKJ6j5mDnJDLD
zwnbE4wjvbHE7vTvPleYVVMlZL7+eJC/wWrFKq41FOzJTi/0cOjwtkRCaMC4siX7EE98X/XYLr2v
VMdPI1WberEXxBZYkQ1+yEagLG8ZhfA1p4C95dBLI/enpsEMPsNf8cg30ax2bsMAlD9BAU0uLzt8
0dCtrZR3/Vub/QAjGgNIVzktra8dBfjxev7aijYE1moOv/j3jDTXmB5k4+gkcSmLXWPC7YFPNHDP
Ic5G83EUjT+AHc1JTOpCoOrOxqzb/HthKZ2shZjyeJdL7jeGgOP8yhpTsbz9Law6pCQDR/FCU3KC
c/bJetdRby+XxTYcDZno2egLbm9FKzVcK7TU/PWhYJvO1kNTJxLsMPjunsJi13H4kd+xK3+vhwLr
XPqh0POQrLVinn+n0RoU9fUYQZo/GCBcaDm7fNU45Qjq9hHm6fOMgiMN0G9RbpjdwlXaxZfenD1i
wTPhSgIPdt69TBsqrOKI7YlIMnYF/Z//ADPUEgFOTnhypP0FL4V3RlkYCSedxbtJk55Pnk1BbMYj
GY6RSPGYNjcLcHD/dKQvQ+fxSPyK3ZfdnGjtiXWk2qM3sFjxh53dU+8oqrKw5s4FlcHB5/aj8Vo6
96F+H2M3T9Vzr/3vHVX32WFmm7IZXTHiqM6Eo57q/xbTVGbndYGT9E+8FiJyEU3T5cfnPrRKxah3
qstUVVn4//g4UgKfi6EQXGg/xptGRRecuD/xs9QyyyZtYSwe6pGvn88ur9LgxbloV/gsLQcHIK88
s6KBW8cLY6UsGr6etxFHCAQdDMCYE7RZO7DtJC+57cLBfqaM9PTs5vI0qA2yNY4ooJ0xkL2QlyTm
BYv+8he6RgBYYk1Vkj/OYiKvclGFrHT0q05sa/Kf9loEDQcdI4lOuXcrr9o4JHsdGscnfhKoODl9
HLkILL8ZV7l25hRAO0ghm3JlGlI5nlrCm7fAMAA/8OVTILoNAHPq6VJhFTEolXwOi9Tc4FtfBAP2
DsYNddLR+YZbShja1D9LEs9h2TSnKJoOke1tKLMPMi5vAmxC1FUrv4R03y9lZz8O6BSSOc0+TaU0
1g7CHFDSTeEgj3GCK/I1Cih/INId8EKalpukYUHtCuizrKZh/M+bHsHwJxpdx+R4sqBISQmZRjtd
QmHSKqme+TF/xdkskEn/p3MI7A55cAHKICal8uKjhM0i5E61PukDRbCRSNSMckOo/pzUlvhzBm6u
E5t1806gBVpF/J2StZWmO5A/DWK1mb7Fxv1VULrBTPj/7fKB6xu28cS69NjtTXS+bwFLK33iT+N6
B1g666eSM+sqmeCPKiRyPlZ0rA/XTSzx9acMcbGuWGcSQPcCVDXq9mZJQzxwhvncScz+oDFhRhI2
tBqmw7FfLSJa8QHtqTDS2FRkj3ylm0kOacGUjXEI4a30Xhcb6RvbcRsw3k0gbLbAsHDXYeBYUV5o
DGGWKlsStKNodUP4UFzmA8uuEF2CHlTuh9icdh4lzsVtgmBM/0IOUqncM6HGh0tRzdHLwmN5WO7S
kXR8JB9YuL7Qk0JOx/zdnTEypc4YW5HbKMl8GZCLlimopNq/Wsj54kAuifdCxHGp9wOMIfNwvNWb
gQLHlIKpzz3rS5lKH9Qm1uxwhd1U43f8vfp04ICse0i6dh5nTYmoxFdUihaMnnRYHdq8EIc6M6CO
AwomTW3DgfLO4d0wQSUVG0R3ZVpPFpVCOr7zQze9jQM+sGh6iEg3XbdlZDUohga6FfBEq6R0ydxF
Gx22Iyt0CUff25/Kq/hpDdveivbYTQ01qKO3Zxc2zoO1ntgp6W4h/0Ff7PxtuYoXnG7SyrjYx85z
i8Ik2LgBIOqqkbg5dq1CsZRbbhGFSBQcXadgawucKHUktzpfboQYIN2wGjT3ZdRYuNS9JbnlZp+e
1p4HaeFw5DSz6z5W51CrEDRw3LB2/EuP6g6yS7XtCfdiLPv/wE6inaL5dEOSpi0dg2Q2L6fhCk0B
UYkFofQLOkCRJMiTFJMm5n5Ykj3qP8u2ajxrrgQQ2tmu0shHuUnDPXAASnrMtEmUom4I0/tq9XUB
d7YHNHZ1MRBV4iGoB/0f1qg7sodwIJEED/bC/rM0MsO9PltDNzte/bDGNyYJ3lqQQhq/0PZ6Ulae
PCB7TZaPkjI12On1WWOzLVTyNBfIyXkToynSSM8X6PjXLx9gs2wuKDSk++/vPb8yYmMT2WrTvm+m
qUOLbtQMzqlzyJj6eyz2FUTBrMeDszccKwnBSZwaOjBKWB/7jMSTfN3fL9cJlcBse2BlNLFoLjlL
yHmDPjRWdHLtXVhSid+Ix2u8SOt584FB8a28MpJd4YwM5H12l4vwaNk1IDSUG9mpCectrUr1Jm0n
87Enpk2/KARyIXfpj4wTTHjp2z2Nk2A4OWMsKZ4SPJk1H/CsU3QdcpamldhYDKcxjNZqkNfLui/m
gUpGqD3Ztnm4WZGBAw9As6tglplc6rwYWhNAQ7bUxLCxfeW2n+gPETcJnduuc5jFy7h0hj99eBoE
RK/IqOXBo3ZyWxQimLMcyttOwvSS+DmcIA/ACorMqfj9gICWICcUPnnPug6CAVI7uAmAcHWGdEVs
GpfBKZaiUmgnzEVi/Pziy5zQIgiQju0ZKenHS6xnU3xIaKDVC9BkWTWjFGpbXwGzTMSzbNs7hoZE
I4//hY2nsO8MzztXyk5zJwTo77uQqLZ1GSRUz3E37+bFO/U0mbSKVPS6GH49FBq1reBEt8obuNML
ip4/VdcA39jAf7gt/AsxnAuQgyJkQg1WtgQHdJaMxYSxFhjZ1acpx1WCD/FmaRuV+4/ZcDbO4ACG
6oz+vDyYcPODPiW6Ne/sNf0y9eAQ64OvMN5iIFKeGhHa0m9qVcKWbxJpQxZ337EzJfnjFvd8uqoj
itfUMR3JFe3I81jA4kWCujplS1JexlOGzSvKaBv2iEtDuG9KvAkK56hWC13IsDbWnhRjKBHcJDy7
mFJFCeBuleJQf1/mOxHblsjoWpMYpqP/2iacBJYcwmjr+3aaXsYpnccJHVZMqVxQPBiNWg1IysAw
A6lCk+YKwdltXjoscfMfwAYm2aNDMopRI9dlmx1aGBgyeLsfPV6Ld4wQOlRn9DAt0BN0K3Grym1l
VpV4Jrk1gv1Zv2FW+B+Wv4fbwBt4oI3Jh+NIbAKpxP+M3Zv3EU2C6EmWRFQ/+yLIMjHjHNIPE1UZ
szRid7dN947XzM0lO4XGIG+Yd6DAMZ/qapfu6mzM0dwEwRAlDrgPKNPUusMVEPi2pgQZltLF+wWS
gWnTHQM4Lyw401ENpFgw7SoNQf8rXDMLWVc+RX0mxMihuQzqiby2H1SLFhaeNaTpA4EbQcSuyD0S
3B1thUD6J+U0N0LjL38C4L6E3OB7EnM5o877GRMPq6EZ29kIsxEs4J0RtBT5dTEW7Kd3w3I4NHpJ
BnrJAEJJdS3TxpO8TynadXLVr8CtxToVNuc6NwvxZTf1cTaPm1aE97fTz6oYBQD1mkWxB/4Q7DUg
jhmBrB8uVbVlVaZCxRvo5PGk2ZFb+uoEmBGJHxHAp91N+rn7TsBPGZXf1iJK1aoQJSpPRKAP231J
m2St+xN8kEJ0ba+iEeOEmaKfWhgSBcO2NIxHeii7loh69NsHDaunLtzXvbdRkA2z/0vXyJBJ0ZMe
D5pNc7ZIZHZfHLnv8YCAbI7uUUi87m19XtGLQkqjiFEFEkKm/aGlDVSpEEL+4+WgelrcLYujm5fr
5rdM6T96fGJj/jCIZLruGvvZJXHp5T3U1sCHVQOt8WhMhdWSH29XE7n+gKENX4siGKRnljIrq6Yi
H0Du+qihSjhQeZKLf7QJ+2YTwxrSFRGw8MoHXPXjEiCFQVlaE03uRmp61SDlK2uOXz654SjF66/a
QF1sSqCdsXImGxIcVanUuMxz/cqIDdHDzf2hvqFjoCnxaPIgazXATDNVAHR2cydmFPHQEaSF7PSK
Kxlw/tg9Lgj5SxoYMAyS+kYuoSasxbj/GXLXMW8dNUbGm4WMuYW9yJdA2Ryz2/8c4xQ2GGcwB2on
mYXM9TSJlJ8UNPGB7BkzEoP6qSG1tMYwStKn+W0TzLFKV2R//jWpflUM4GuWW6YielT4+hkCA9gm
zxQIE25oa3Tcqab7Il3D38r3sW7QqWBXoHma9sxYO1W84MI5nJnBS/tOw0c1zhJQ9rmAtCUueZLb
r44OX3bIDa+1x+io5hrT4u1tcuQkdognsS2DWYzGKFYBTSLauZ/IQ1ewy9FW0Gd03DfZ/YgvWBmw
0XZR5B4vEjzYkT8jG/Nqa+dv+K9ecpAtAWlsyAFUn0WE0gZtQQaTDpB9Bd4bwyCW6OBKTj0IoyjK
UULeMSJuQhlPvfG/YZLMAs9OYPajUDLbMlE9vKxU4UZJfvspnZpY6oPpP9hKG1d0PiDv16knISaw
K0l8E+qBz4JccU4JqeTjqNRODsNsYfoRTgruIVdWwDpiKzA1v08M1uIEayruJdDqx4PqXsgHFglc
WXlrvkPyQQ0v1LPx4TNQiLmJRJn93vXB35fvOTh+/dgVxGkTqbNi+tu4b5kuP3pYErFH9Aicxyek
/qm7z8i3VGOhF33Ruc+vyK8BdhcSVGvBXw8igRYbLnJp5maEy2Ry+/AJQSjEA1UMz8BKM8WpnA/t
GSH+LdCrtW/RGb9V/IFLjmDH9cGyyaxSwToSwEtiMg+kcjdlSzDzsHjwdtL+65SF0u8vKVFwASpy
oL2c7/Id+mQlv5WDDO9KoMSlOdjdebDSu4uyW6SSK+Mg2din9qIhy7OYFncexqx+AC3q/5YxwLg/
Lo/+t5cMaR9ygSbpHPc04YI6H4HrEmenNyKM8u4oWJEXZ7w0ZeRcftthLD/uJqLd0VGdYKLgYoBF
lqnqFvSBtQcFwA4o7bgima5QGRwv1q1rx9cffY8cllgk4VrsIE9nvgLJyp1kp1SZFI2BrleSxLL2
2ObDrCRIjZRc0eSb/1FgCBQapuZaESseLCeBYUyTpdeEVzxLarb3pJQtfnx6OzPOLgNN/dCZmTGx
4MxzjgEsOuWdcpYHHyZzBtf7twqf+Jy8Rx9Rkg/xus9/udIcTWFdXIbu+lAyVHihyNbJh1cv80RS
Ki5F4zGRhaS2iUPLXuGpxa6jxnIyagIOzmdVkPZ5uqwMWSIxGyQQxZJKr7uC82VfeFnPifYz56SP
CpU6r0M5St3N0nIimH3KitxX+bL5tHojCRQXM+MsxwUvw/8bRiEcpylMLte5RNSrRgEDHcnjU5Lt
Iyhg7L7/qu9OTOY2+HjjAJjN4IV3NFHqDPXA9jcNcCk2lDkWq+MlSsQyMv4Yi16P4KcX4ru9pvYr
dpKGUK+BCpzTqhRj5OIHeoyvo+SoLWs629NboneDCvQHTuSLTDgdzPXyndQ0DW1F6CK8kXQ2zkdv
I/k1e1HXw12oY1v67+1Z++VxmKjqC5JN8cskEnXpOd6yf352eypYsyflY60+tsHeO+0AgtF+7rgb
MQN+kSVGLQlkCNLMoT9su6xUUd9NDl0dD/376Q6UbU90pi9aFCXwCPPxhkHcfp6DGRFuAgAAom66
y6p7vP/YOr2WUbdOSt4dvayR24TkqsCxASlDdTYHuu67yZQvLsbYEyBCguVVFys7Z6X6WijU+uGX
myly9pZydX32MgPoFnE/gHsxP0aicHwlkxoRAsbkIELFLlf5Xw0MLppGe55jWGgXIhiqxEOTBRgc
yuVQ0LSgdEV3Qms+NGuoDjNBcfx5fPqi8773DHtNftBDrvo2FgxCkJssHV3OV8kzDJmCnckcm1SX
gsS1ggqK3OJ6sesqufLxxz7U94zHYt6ncOqlT4keuwiVEVsIy815CIXhQE/27mNHk1bOWP3+ntUv
pWvrKyZbCasMKYvZT0JqOq1PrSnVcM67gjoRHxsxldRIvfdz/nzPBo3OQWUN+DRuFaZnFK1fG0BK
Ut6I7NGMGpnf2p4A03gEEx/PV1GrH4OLvfcfLiuul7SSJjqMpeHcllHklhLHPSOU9qWYRg2YJefE
2LUiNJaGzd6cPPM9xOeNXQSIWp0ac/lq0Ap9M2fQI9g0/dsEWv6D1U3HrD6TZz8tXkMCKQdMKAN0
pDwDoB/HbcaeUbudsC7EEzKMzyX5XzjVIk5OsgrTng1qLUABPUoiwDsa0/Sgs+J1bi0V6SCoa/zN
0o1NXOcYhC52z2FDyeVeYg7PPhbZl+e0gFCqMlnNISM/Rk/UJ+d+OyhuW/eiRBUnY6LsQFBByn44
bMXzyE6Kivtqi4NDvSJ8SopSFSZe7O9qX64rwe4yGfmUg2AUlL4kYVDluvX/22sYPL3hw2vMOOw3
UOq46VxwPO+Bn2oqnBLn2uQ0Py+wW4HakG/i2BNxqb057x5a8aPVzXGkVYsS9qDqsVbo7c80fJ4R
UgrA/k3iBw01DhlyYlWPudN4795NMJsLov31bNRCRRkj/2fSK4+ZtlN8Ug5d8nFfsT99GKSsex5j
+Ha6RxeLUuQ4Mb57LxJ+gp1kN6l4/Arh96EsdO9Q0Q1ZW/w1sTo/u5KWUG+5B+5JWVfChF67cBpv
eCXKPuEyfTpKsDKq45Mowy7yHw2CUDjLhlJ3wowHtimwv3oDeYi9103vYxOtzFXsrTjxCQ99P8XD
n0USyb14IpGnXXIMoc1b6teYbgiUYDHurC1ByddnHazbVCNXvktgD6Tehv1oL/i6sfEEMa9iCzYJ
YBt67Y7zkEAllGPYEIN/I0gzMzWTbGIMm3Aa0cJNNFkbKungAhgVomHHEt9uC+wGGU1WVnapXMnZ
XHSRW3G/RhV2QyzzjgmCwmvQJWjnMIQRAEX1xwUhCxOqBoQa9WEKD3GLYaD3HnSTL45m0oxO5e5J
BkqPwl3p3AS4GlmA8iJfCU/m1LNrMCDt/Eyb8rQbKETgmZ+Cj2ISF1BU/q4lWdHIqgBugsyxD/T8
VzoC7zhyWzYj3VK87rb6VU1uthLLxPw4vyCQ77M+yL/4HE7zsu+gZ3l1wgn00b7rgU2daysLsMLX
7MA+9ruvFTHoJ5NKla0kueMzFIkxJ+s5PN5M3V1WWnvxhhOjnIMnPn01clXDtRmV8AiBiNkbxH5d
bpMzjnPGVkfCYh+GJGyanihpVm+uVb3QGBccwscvEUObOU+1iWf1shmxaQokKXyt/ThfATGrgmAI
+2afGcvFGWfThiYnsSF4YYSIxWln4/+rDYge1C6SnF3u1NhY4SbJAKre6wn4hK8OiOKuNXokRq8j
ZM8VpDQj7c9UVZyy7IGUgh8t5qE3AqRTPML61oD3NdCtMszVl11rQtiHbqmYp8hk7VKau9DEjonM
N+w0dBVbBnh/2BGw9OhAB4uWFk9CgmZjSd+JrDyFRgZrLR2zk7iB3F/trTl9vdyRok8wy8gkKaTe
53/JLfikKA2g21ld0JnBiuJyRhcVNsretqH+fZgTtwLXQmz4iT0J6e8BIHjNybKESF5RLAHH1Y2s
fkk8oa1ozb5dftOcxsYvL4gjIXwBiLjVAYpAOcFR+izAneRUv420ZXpF28EBaNX8hPrBkHgU8tCU
xMzdIpg9neiHap61U6QwApnWsitybKfYcnxwDZLbFXCdQhrFlFPjEl8zNSbA0E3YrCxxzi5SdqYq
NGpbecOCGeJBMuB17LYWi+/zKCt0t/AIdjxN0cI5iZn8hsOBCD6mQ7RUoGQ+sG2ThLDCbaPMDqe+
N0OT6r9RJmoARS+2nWrd6aYPI6q2TZMFZzI4z8k7UAO9gquCNUmMSD04z+go1wZ3oqxxTVFXHhib
XYEJ2UgB1pwpriwtiBoSOUDM4YM8kRal9Xls9ce0iv33+y5qwLJV3F2PG0pwFbs8paYbV415QTrZ
1rjFYwHzNclYCgKt3ZHWZVHcQIGTlHmo58wSetoK0011atsNd70jNlABv0aFD1pZqJGXQaGReecg
vs+pMtO+9Eq+i+eiUCW1vzsEI+UZ4jUGzSUUAXlVZtp0MKGcX/KWVEoF4dYC+IfKa96sztKikUOx
hrBrII0rtJRJH22q/fgDLhXHJ6DhaDPTqeTgqkZ46hHhsLh7ra7mZpidxCQZ1VofUr2j/jO9ZdiW
IYPTU+o1AmniVqeidhb9P+luSy/iXtsBe+hP+5IwT8eZPh6urvGm6zMbm3RMzz/3Ra6Fk/BUZry+
g3+R0JU3sj3Pe/5q/9vxNh0G8f9P6HcNDitOlwZGKoT7yhgRvzCQxnKuzWh/aZ5KXrPBzLsW++0O
KI7gjKIj2KoeZ+aZehTe5Sq9MeaVrZCGcJ6p3tk2TZZL+Cf04SJ7xEZZWyXsYBaU6vo0Xl8QOjBl
/NIcn8YutkxFRCE59KMnVwb8tB8h58PMp6C3N1kNwmR7RpPjRa/FbCVLYz+P5VlR/pnxCtxnD4/9
OfaUCDkoJT8PdonjrX1HGr5ODh+UyacOIMfImt63CFwW1YtffclZJC/2dXtwT66xrhv4J4qDbXp+
RmTa4rJ7nv37ijtSrPcI3pIlR/cH9GucYcgFCswkhyVdSw0JdcvwzIr8JjYr2ARGZ+9To4J6w8FL
JNgZMtdp7O39pOZsuOUScLyEyVPTiiIztDgD9sgExnh4uxC3JX1QpBUJljfEUZpV9/zkTEBHOvrz
Mw4yrnUCfAFXTAKJ+lXIxB8spaXRK0Rl2vQFzL/h0X/d1uq3oVy9w8gwMdls1DGqOUkl2LeTkQZ4
AhS57TKAaqtHfho30UShpD2IrGCXavqZruhW9kRHQRK7eRhdTkbl4a09ZmY9u5iEfR9yJ2VWreNo
3fus7KToALwVJ15jqaTG7Y3V60nMGky3MoqCNFygP4mecmFmXzafP6Yd3V/2O/LkSYExI4v+CL3F
+JxjyiDnX6Dj7OxUj1LAlyHnFkIjd0vyXD/IjUg2KxmV6ksFgT/+nWQ9jLaqR+4eTkAfsWa70Yia
EVPPV4lux1qDnCN7mVmfGVD/nJ8QCGLw27GFzYB9q/fddhORMSgoGBp0J2BkabCdIeYiYJvpDccQ
t4RbKKFNurSk0ew+G86d4R2XzTYB9t/6Zi7rrG/QdR/ZYLAFTq6Pg8rL4XULRlvWqMf+CywMpkqL
2yrtZ9NKJiH0A6KKMuiXUen6V5ZLPE6SrlqJ74diy2WNbLt+aFbyoAuW9CywLBvbEHxoWcpvvobC
Hex6w1oGkvbLDlz+EN5JokpT8gfD2bhzHMfZrq9TbondRvuXxrEEtX0P5crnUPWYKGZg11RqgXkb
dStmZRhSVuCQ4A5CTk+TnY60pxyUVIB8iCiv/wXJJP75r7UYG7DYc5/CJ8CrxeWnRWSaiYe38CHA
nucl4+lVayjpPG/i2jANQ3Aif8Hl/MykAWADpPZ8Mm0pP2aMFMQzHsZf54cOGcPZL5fXkcxxGnQw
YraP1yziA+b+m4RVdFh0E94BA7Q7S1HKT209vUiPD/hQ8C2oP0Sql4R+BVxAS4HerIdlmUR4em3j
UOIFepX/JiYoSvhRbG3/WCBYms+1JGgEJAQIPJMWhf/3+gBYZGBq8ZACRQclKu0x6fqEqAUQHSZP
7i24T3gcVOw04XvkV78u3Jmdqk/PH7+4V7m7i/ucFQaeu9PEMvx+WWWtdfvgL3tnBH2OVKOVUNAP
a2li1rzl4QJ2sBS832Zzt9c/s3NG45NCK3HRMdu2jsxCZMiIm7IkIqR6VHJThAl7NxdkKkluNSdT
MhgU8R8kGPnlxrIddZ/Bti4v86X6QC6ythAiUVUXJQC3Z12SVBRd3uPqazpuOMOf1luJyb2HSO33
8ZPX6bib0m03OcSKud1B3CmyDzB3Fkk9r/FVjbMp5gCtDEQLeKPZO6eLZJsu6FrQZxSd4C3YbJIu
89hUUasOA4uDR89nrAlwAM4jm8/9cOjVS2yKZS1p1sNhmYtr+sz0pwpbOAU2ptkokw1vAZr1h+rj
7f/G7Jz8wexNuN+16Atbs5JeR2H2kXHw2KnYU4m2W1LNeoBDTvTLlCE+OJIR5Iq3o5X8gsXw1ug8
BWZekdpgnjVMMuUrBaKTvynz8FxZt0iTKIuG3o6mms/AYW4BicSaANY8ZziB+db34IAxGr2zgHZb
8qlxPVzoQ1KkEayabI7TETQQsSyCbeY67gf5Mq7PjDIMFmU4ItRTGu/1fJerq5GaINUlutrSeDWw
5ma5XITQ31NL1CkPpw/eKwha3MslXcEFDq+D8HqsJBq9EmPc8g21y1T07KnDV9nX7g3r9YJIhT5D
Ef2foNI0c7kfRw4WE5bjmew5Dq82LuaXI+6wGgJsXUGOIxvhjDZPHc7QsVUaz1Y+hoqlrhaAdiXn
Sb5/Tv3VxaE3W5a20r+/cJ8boGZ8c/C9lPafB+2F23dqHnklEssCw823Sx/XjDaMVQ0bYM5X6Oat
66Gt4zrqKU8bMgbfM1UOFfAL/EkowwFstNAJMuk7PA9WxmDqnM2mcPrXyeGGmKpYHpKfwZA1MJOM
DzwwfuswtbxOW0/eWllv5ZXK/lDdsqYxJSqIwLGL0yuYbZVPxKBRpFpgdb7BI/bcXWV5pZSoVqZC
C62ZQOUcZO9yqsM2wWW+4cwrJQSSukVDqcg45wr6gTKaNOsT6tBork2HM5DahOLKtFvF4MCSh/kA
gUUK2hBPbCmYFLzt7fy6ebclsu6+SAOHmt3zGuymtK5kMnkfXn/BJRxuf/jM7iZ+Q/e7AZmlQGVD
GNEu/Zath7XDgF1KzNJ+X2viRLdEBXWT0BE8aHLVF+wU4wBJdw4+bBr2SzUu03x5wYLpNksSYl56
EaiG1l7gI2hqkFK6Emjdg+9TooMlI+2aVTNtaZ/pbortGukCT24+9j00wzvsFOslam9TEDddC3Lw
cvRXgmPKPFzKsmorV4ukdhlQXholteqG8AJR5j8MVpTya92pByIUwiEB7YsTq0iWWuvB0fDv1ZVh
tqMl8yuTS66c4E4kOP/NHTHVztfB1rEaNE3Xrwp0L5ptdtIFSsBBwexoIk0Qdb0bPLYq+kXNvBTq
DCzsI6GNqTcGrHJolh736/z9iFDBNrjZuFj2+/weKk6lzRYM/vB4ZZlzPyGALOFyZFbcIC6Yg7bW
kQrCmNqsg4G0E+3WfkrHEgVN8EuC/TerwEedMzc+1GPrWirnS0L2IVDz20w2C3W7hAvOQu8JsQ6N
sVw9+e/+uDdW/LU3iRoALkr/EeWEjWjhsbSSc3wG0QxMlfDurQECvuLaBPWuSX1tl6C0rK+OIfTT
0tWHMQKv5tfJ9OIDofKLrkJulddjXn8wcxeWcC5B9dzk2zW8WRvGQ/QZg1RllzAK58A66nGftXvH
JWZnuB6ZZMolHq/UXahQDGWBviBSN79f1zHYb1iHEXfiiz4Sj3gQth5cFByFLfa5LtIEtWPZ7zdk
DhtXZYGU13/xevehGyMvrBIpsEqo5KRO+RrA4kft1cLvkF3vbQXdKqnTOUHsLvxrzI/MJzbGtCEw
6t8JT5H6kPuDirNVkqTLyt69d9qtCT2CtTca2tMfaULdZGQsfyhOmvv6tOKCPXjFYV8g/hg/QCcn
QvAWOV5AAYGD2JXo2C1yJFwJ9Fv1EQSuH1x+3fwFrhbbp8cdXkr08uYDwf4ZDzB7B+JsMT0IM8El
eeg7ifYF+pivz98eRP5Sm6bMyPRypvb/k5M2YkXnjk0FJ1sWUOUTcuv57OQQxk9yuHWZbUTB6Jl4
u+wGK33UGfoE58n5zQR/bX1QpLlkMW77ldMdDkV+kudWHuirbR9mfLcGboim/POegwF/XQfpt8Bi
kGyHthst2wOMRoUKh04LMZvrpJaEb7fN1oqBMX5W2Fh2e7Ms5uFaVimifUNmcqMAbtxz8hw66ZXI
i6lA6Dyos5yTXdtAEPepS/XJkDqK7a75G3uwE25gdl+em7j51uEvkmgM8GRNHJFWretWh3ymLBVN
d3ONNrfA7knswQ/Z+eci8OR02rFN9HPQV50a/DpUqmNikANP/1USATbEddGy0kAA8lh/+mQM4Nf4
hfXQigHS3/hh/Djpa5tUwEUltmXcgOVnaB8ulaIXvYmxp9fxKYt24gC1qWBiknyy9nApZBB2m39J
sw9oP88D0fbcUiwcRgs/yk7tHQXrUZ48TTRnhZghctNpHAEfqGgL0VTtISBGZzh6KZRCfRF9M0Eu
r32EFDXqzmGogPlBWkOiGLzstqCKErgGIZY8O0ykPnabJ78t8SUkDXHzst8xW8BTwTwGJpjQ4zgg
dd8e4CZGKL4PJmCQ9UpdhydBoZ10UDn3Dv8eu302gtxuLvBKSO+TABY+O535EqdaXGhK4LwP/W1x
+VTiuq3PyTuMMgBlNIQ0mW/GDeslpDL2CJc6dRmf3lTz+UqJjZDEQC02MqvI4n5nyOnpXAdyqPmu
wk6JJwVFcfGVP563ivRuYO1NkCB5H03gJoJvI2VJxjxX93ZwyF8sQXE7iifK+ltkY3o+9iz7oy3C
Qpub4U5fm4mzwl/SRCy9nKxDskwbYO6uVFS8ApplbObMg+8yQxfv3GGzUEkzw8SHa922VCvU/3o8
9j7jtVy4AuQnRwA84GikXjaeUwe05pueNRNeF0cdnxZDbprGeKwc34iFXSr3XW+RjhbW7tX66ue0
qqAF2D5DtN1t/avThvThKO1D769DGzpd4B+xZ/cUqx8Bfgm0+AXc3BthEct5QZOnG0hQRIyILcYs
s8ajJFW16c7Sve2sSICXuQ5v78pCuLWs24eNBpio7MAjcalA2DUGqliMaFAJ2qOVVEXNKMZHKJQW
dvD3THZrx4179PrjVuGxU/TJoKkKkHPAnmHR8GFjlROxp0QH5w2Ri7wJ9eAGAv/5flYKPhOUvRLB
7IILrgqjaU9iyP3GIMijVggn3kvWVy2tpij9tvxzub/ZFJZyAczcoOIqVhZexKfLwon6OtqqoDzd
I36atZyoXxZiNG2m8bnLLy78LvGSGyvT+oREmGQeD9y6UzQSCJKWT+IIJCMUWdIZD6AaamImooTA
tnF1x+4GHJCK2Bt1sS4MN1j5cJyeuxd5Gu2GowJayvx9Gu7REnGnzrNRKLeXZVs0TNhUzpEnRtKX
9+n+FzJtc3fMygvoKWoYovAD4M+PD87SRT8OU3R6k1W2SVrM2SknMSwuajlh60si9xxwvLLzI+05
2fITQWEshAhwZvvrTOPVYDg4rQ19eu+OzZjCwGszGJmPMBjAXundaqOCMTmJInuluePAHydzkfJP
/uNuvCA9Mcl33Ga5pvyuizf/09h/wlLIBnn7QI/693keKCsyR6IJVZwgdGpht9j/dKLEBnpqKzdK
vHkQ4MrFyjXXpqXtpd2obTLN+gklxbLG6jtQkQtw3Y3i/GfJh2fXncjjRN+L89zKj12JEKqpw4vI
5iG6RLCZJDldNyoVahq2t8ynJMfLzXA81rgxQKWok3fJwxN4+ENVWfuJoRTieWZriuz6HhmpKS2Z
qTupk0cbTeuxTGt8/RhAl+oGtzIOKUv8qgaSBGXJxnL9BGnyhmgB1oT0VoZbXlGOwLUmpCf+HND5
gGRmTnsm1gRFrX2onVszcu832y4HP7zxZ3JtnH3J/D0BGkmORybfQz5Pt1qzAO9pqYzY6pxjdfpr
VM6lkhd9avjm2Qqyfd9+NRMwuxRdU8ghRcxAljWCu88GDdikbN/6Jq+8rIZelkVGDSbuE9WfwvQX
eCzqYzY/yWr2vnzU5R96tGpk+rPepZwg/Yki6Gdp85p+kvTSot2ph2gVAtTo2tXDBPaJp145rIRs
8IBLIL9aCmSXQeMxZeuGJpws2b6IT+pj8mOM78UuIKZtD6s6K0N7PFlai515dltOo3co+Su9zD1g
9CFfDiHYXx3lk8G+vrSb5iIW+Dh63E2jmdReTdhaWEyY7paFbhi85SHQTD+SphPH4of9te+nRnss
I9+4MBs6gZU38feJSEJyZCrnlhwvL6EUhiSnSmtFVS4boTP6uPW4iFDmU+FIFMyM94qBJXtNA/CZ
Kx1ahNf0OmUyd5GF0HW6n1n3f/Hzig63OHOy4AYeDZwpNQSlaue3VdG+T5Mr2mjSNf83p2E979TW
lHCWInyCvWILmZq+yl2ikcEX7eIM/RI2dEiZy8Qx8jzx+2nzPLob76Kb4vBWGHvOkRPcz9I0M5FS
ryEeg2fGXSdp+oPPEaf6uHIiuckZ5pVc9uZYPV7Sof0BNRIkBb2KKm66EV/rDv8hYaDc0AJsxRKI
rLJ9RQQseHt4yBV5Fhw6Bmr2prZbOlt3yCnFlCD80F7jwgIsxL2FOIWk8rTIbMtI6/xbNSqhPj+I
hrdmVdYfKnvG7+5oybeMqZvXoiH9RjgRtPJGA3Nkk12YCRsb6qXSQVEUlKCVZalNRkaH2ABFrCXn
R0bi0FjgE0+lh3ETOMgyagrVf/3TVdoYwqepf3AmGw2M+aQIknmRlUAHlKy+JM3AbpKUe/+Mn7Nu
eajITShWIpy0tm1LnVzKErcwbUNX954l5jqitGdPb5wokwpSXzvvNpNGX4GPT+cwT61E4Lh4TDL6
UDKZmRjfS+mncCe50urHUUXW4RwPq+VQsQkhTL3aTJe8L6Z5crcNh4OVr2uvhCOECPA56rKhKjqb
xLeyew+v0WFxENVsvM+77Uwd4RDqovoSI3lVTO9jkTpGoyPncyzWR9jLSkz9U5+rUbEE31QHS0eP
nkYA1TiDg0A+CynLqWNOcJ507zfDH9mi+gdZ0ReRSvCZofyyb2HO4TN66qK2YENB5IdEyaLid7wt
4ShLP6Q17GOQGjvjYfnt0Zs8WSbibSUMfTtDdL1MfVo2+gpxXSCgoRONHK6JnjhjX/MdI2bgBzQ9
xJLGH4yzVvRaDgSL6ambNWBfd4T7HxI01d1Kk/1VG9YiGbkpoVQY5jG760EpcHjG+2suu6+CeK3Q
BZ6//ks5DnluR6quubPx0zHTWLJEe6fCYYpJpY4sbximK/votKNo4ivnhFTbm7JjCYA3DcCZFpVa
eHVL2rXAAKgfD0Th+CvF/heixJEnxg2bjB2DuJjzH/F6kMcJGKyy3c4x3JDbsR3lN3LmsfiXvcZ5
vSPVJ8Cpxf4FjnSoBRKRbB3gFopXJ6eVJuobEMxQdAD2XFatzjNdVBwnEdXe5SdBWX4dJBAekD1w
CYb89ae5t/2p+4dL0fuPeVUQnZgy3gI6/OGd5pWGFXfzB2OFqVWY5AStTKbQQtzxktPpt2V9QdPF
5EMHA/QDFaBeX2tayIrR0gB+icqhWIWhjRJFlvmM3Th88SHd6+Ym40GbSrp77KoNbgBGKg/fKvAr
AFBILhy65eroWONYo0/j68p61al96YFBnmS1OC8w/L3+uafhadon2xdShG0bAEXDndA4wV7ghrUb
pf4dLXatTwGzNsLOTd5T4a8QD9iAPzxLZ05oc8qkQ0F+ix0n9vgFspgU9lMzbDqzu+juI36sZ79T
+/BXWXpfc5iFCqRLV0bmxtBNrUzWDAIRqI1c7zYUaK+OcScEHy670ACXnK3wuukCF7L0Y493xcLn
mEVmbMIsE63FO+G9VOdvMj0LMTa/atpNoFh+KSY780J/HOVAgsdWddAnhgmBOmNocWp6acL/QfHa
iRl81f8dF1g6QCz11DhWAEEaksXGXD9tVgAEZ6/V7km+D8wkIpWSm/IzPrpChihHkAiycY9kHUmi
DHkrtKlJlvZSSiU1bgbTZLiQ4kPKP9/d43IUxuVJxtdXeHcbA4TjZqVK5eV3//Vna+57+lbl8DYc
izaXQUwaF5klruAPMS/daCM/7Sdmz0Bhbbo94sgOt4wuPSmi+sGLUlxtrL8ceJCOjtaI2Dd6ZIaF
esqxv0/GMR4sDuLiinZ3uuzAAoLVZPRDLCkP+oRYI07Xm3e2P2KdhN13rCNbB/Q+SE2gXPxzFjfZ
9Qig0K489sMHluCqG1C/Sj3mxUTColOB8gLHDp14oda8iqUgZZcPdJfW0jE7zx8+qg6+MXFxd4tP
S24Kz2nCYuiExTGy5kYggBPbK6AdzTi5ajxiUufAdXWuN6SG0f7DFKqfGMX6wuh3TZx3OkiVheQC
orG37xjx1BW9NDWRuywr6+OB7oOwTErb26x30nnqQkxTG2kwMJdgkEjJDX6fqXYOY+fsKR4sNqRD
bfuDg0O3DC2g1dFfuJzOHUVX367AMHSDfjGI5eQsb753rLPKV3uYbFyzR2zAvBDSoHZRp4bBwwyw
juA0u1c/MEXQ5lIdHcTbz+ry5oqjCax9LEriQDf8z24ea9wE4uL+3dLO3aYIx0B7NKAwnAwSHXHR
aJyIu0L/DggyXmqUCiGWiLlstW9tk/MAlJf6gt7kXqr/pnulU6dF31bmxjDZ2Or4fduBiPRWDmYl
b+0hQ2bi54oViXaOI6669o9ea3i+u6Z52gZEwX2vIHJH8vc3GTxHd0CoYMUzD1eurxsnIvq7q7Ba
wruwLuSWSiBnMk6oh3krvc5RB31Lbk0RYuHe1+Xhn7yuLyXxRrwdLR62ZvF99RyRoF0Mu6Gh7jIT
hlkKyq+S1HkNHMO2wrnsGpHW5g0/G7kWCD1oz/kHZn3dKUo92KXH9QfHtRVEisUhgSXWzgaRZ6In
r1wpMJxMUkkMIYaDdzZXSOp11pmIWkvC6AQdcCjyDg0cfu0GFEUmz+T2o5sfQLz+FwtagevCIWYg
rRhE1+wfSXfUFug2+cfdfAKw6Gf2jfC/HaS4GFc6z/mdOKPud6DSuoJQkVWqGmkbww4djZS7pUi3
bVyroFu1aWe7G8YJGtcx9e5aY6vSKSYbnGwYBdFPf5ZPJlXNNHQ1cU9YiuR7i+Ui2XcIZH6NZCnr
FofB2GR3eCxGd/HKApneUNqZxdSNzRi7Sf/BhbXNQYoqYDUIo9vIiDiRBDJynT63JU1Vifs3FuAn
ddIUPvZ9PVhp5GnNOCt+FYH0IFJMS2UZFtvsxWKjRbeoqtu1fIeAVqTAHEAnv3wh0pFpr6wa2Jfy
ZHrIdxtX1nguyXX+2uVMh0YYQlg11vzy56vkJb1KZRY8dAq+RsNIDVXf4FiRw/bJ6S7Isb679XUy
ZQUOuQg3/bvga2GXf/qUoDj5pIQfLcg0xFu2MgbufG1lJQY+iGjOG7ReRLKLjAcauNl887JrjOn5
gJJXBgpWPFxTTflYUl5W65XyA7zHAzQgumpJYsDUq3zuorqfzn/Tm+b2p0sP6Uq0kI1fLRUWyVNw
2FN8PSnBEJluHlOU8v4kVqDR+bVuF31tQoy2j1dj8yakxbLatb/tclsWb6YU3mWMApuCE93ymK2E
hii+GYQA2f8RDAobH66IuIyoiwSwL51LbnJZVDyzXEDbs6+2g8qnUPLRlOILt05kMkEegnmczYEb
s362kkwh+9UcJwIqttyCo4RfJ149u11r4Bi53AK0Ek0aUKKazcm+3dIX0lHpicvhAT/b3jKBZcQk
eQ7n+QGS/AbqrAnc7yukKgtLfRHQdSwtgt0NDwEoiTZsxKFMYBgdhu9RaNcxbLZB8fuO4BPvKwh6
WjA+f1qamLkyC2odcrDv01uYfKy2UxJcSGDZtkSn8WZeuhlnFi4oxHWlV+smRY8ReLpZWeQDLKFV
gHxaiU/YfZjqQCKKU02vU6jXeabx0hnz3TSejEsonJXTElx/Fgzb+dNbx2eNs+vn8k4SBZnGhOof
LfCzMauymFfazE6tUV34FdPPj8sMurEbN35n4kNPs8Rn0gIVNm1sPm/ViHZHw8vzczX4pMgy/Bw8
QcODu/lVE3hTda89FT7SAMq8OQyWoU5zZCKQFgqhrqNl/8z84Nnb0whqKyfGtwh2mBnrQF2XILLx
YxB+hTT6A+phUwJyVc1Rwru5KSwgXQnsoBncLyXARgQgHwIvIzpOC6GXYSkNdtHOSEYLzStQ2Zx7
odcfuIVpFA7LOYENs0h1jDSQ1LkyZiuaYtnaee0iFiuTlnhn2FW3iM++NVLQYVvNddOygj4pm+hO
zsI4ydm0OkDSIe9yU+AMehPd5mP/LedRGG48WLtJ96NsQkGMzzp5wfumDAiruc5WSVg0Zvr62+oH
c0Su5kUDZq9DJvqiWTqpSEMCPCT5yztbqcVJcGTHC+BZUAvduy10QIMQSd28kOZSChuyDiquDus7
AC5ie/lJegqvdB7m3AlrkZnDCnsv5D61Z4lcd+5c5cPrJVoxMp6YPgZ54Oo3MJ5YwmoVBr78siq5
qi/a5O0Dd7VujT8fI+XAB0VTYZDY8ei8onByIfgDrpouB0pInYZt9vzsCCKAw1GEqw8HkamaaLkn
3z2FepuY/Ur65cHJhYHOtG7gs0vEICK6FKKvBqDmwd7JvwtLOIMPgQmDI3f3vR+O5cZ0a8huY6d9
pButFaFJkqVA6tjxo1bMg0AEBAnOrMGhvkjETlj1D8ytxAkopTqx90yOckmiMpy3H5cpB9YID4Eu
275BaFSxrIspjfsqjt7E+TJgSktGZEEUMd7YCWgPSNtxv67qwdJOZ3wh/HE47RerM6YAzFM6mpfF
quKEAiMgxtJ3ehoXHO66irq8aE5CFrOPgj1+fiNmPQl52uxeNSNBGWai7zhEAC43SjK2xzXJ3Rk9
t4NZzw00rHLD20RkQGvQmUu2SwM3ynNArPhq8CXD/7flTmdkqK6aYaY1ythHd/lBrNPQfg59Az5E
epdR8gsaUWUqUjAgsVofVwptMU3pBy8J2OfHaLIDr7DMC0NCAMyYQMCRB4pSpw7Mi1GE1SDCd9UX
VvOjOYfF1SBILM3lrh5YHp0bhbiODvsz8hGVfxs5jyKoPKdPVBnk++rFTvVW9wkRK1w1hR8ATbnx
TCBpdUl9S7YlYWozdZ8eRYR/JET1W207iydAjNmNKVQnQhWZkJZRfDqmtxwMXnvvO7Z7qX+KflKP
7BAq5zPSXsYvbGTcHlisEs62v6nZKH2SdNCU1ISLALVSL4dFBNOFZmIGDYDkrR1cIspGYFPWj1Xl
IAtVhFOss3p2mjEwEwWCmQMa0AaAxaNkuHzzWdz5c5hd4PV80HyViwQbiQu1HYNLxWat8NrUSmWp
j+n3xXog4qDkEcaL+DnqBAh02FD0tPl70vqprSyXdu5P68UHbuJCOtKG+jQ8ZWrgBKxDQEY58VVJ
auor/Vk3E9LHatMAn6JTcdHcbvR8LAAxqwAxTgqiLRR7pAL/joYs3fTmWXDFHgVp2auEI4GKfJU7
yv+843NDbTW6xTKfghpHuIOihUTwhr5u6pIxP1ut8zC6rcEU/I9mK5lwXiTAQZUSuow/2Dbbv+57
UwfL2Y5wfMeciFyb10//qbBm6CZ3gTO42qpDNqXIhUS4r7wBQr4EKNYhbJJ8JyfIWl8arMJiffHw
RO75ua9xOjFPKS6xYnnRDpQ2f6Y4EylgQFHjybGXFfWakuPjpx1DLrKkwX1+tRHnOWMXti5v7WTu
j0XCIOHJoobBQJrSD1GqeQ5ZshYxxS7K9IEsR7rM+HYdLHbEzKYjKGeV2grr4WOJUTuXrx6h/IYm
XlYgJJGoIFA0fs1zdugGnCKJbQy66gSMQBCmYY+5UoFXORaI8f51sg+VrD26foWu9XrscUXAqhSw
r+/Ss1yxXqvg6si7RKIwFt9C5lEPv5EKH0mZFOMOSP9Sn//a+mlWhHC7qZp0byQB9HK1By8tuyb5
ZmWUn7sHHyXK5cxoM29V6OZvaqQqkwymIyNUz4YIOkgpSJVU+5m0RW0Pnqfk1rjJoUpmdQTYGeVB
RA0DDu698i8QMyPOzGJ96wcbGO/SuHhZFAYfkyhDXJq3ZVXYTFaQKPY/DZ4NLdSKvoWk7BUL/+I9
6B6EvupEWTde4nQCQAcSX/wIzTdIBblrSjQxPv61voWYzEE3s5Rqay9PxxpsqKGU11LcX2D+I8rV
5un4yFdmPYJRMdvEOMPNpROGlolMjXil7F0REQl69ONivn/1FIVM0oPVqmwHS6bh8XtdUmBYXaqg
PaXMfz4pFaU0F3RcnTE0CcstD5DNX3legnEF+DZWBlMyCTrfyoB1jZVP7peNO1swPZ4Ydztnz9vL
syMV3jP1+g98UDUKkdedIn/8EAvGQjQkkLTWMMxznBJvDEaQJQfkCOUj3C6apEUtbIip0wEn52u0
2CLxKC2p5S1tn9n21yGdj7O5xcCYfc9snBa6eccXyvK3mKWP1RRb13Y8kkjJvOXXeLSO/mwj4Wy3
9BdiBdu03/fI0PpJJ+KV8OIeGIXmZ7ACqETQ4uplW+wXDmKEMmkVMdsiwYqoFtq+vHjBVRdoA33W
QLd2I/1rOXG1QreCm8fbKi/UKpYsdzsxMXr0voU0sXSVNK2xExEm0iOEXJhrMJ1IK0rdUVYKK5wD
uOOGYvKqKZJqDbzbaKZRG+aX2njB+zbGpsr4sNMyGyLjuT/K6PLwNsArGCUj97qBvwFPC/T3aLQM
UgyswuacBWNrlF98XXonmX4YY8Cjf0Z+uiUnbrlPikICqRcp53rzbWKVQVQbgikhV0i55ejTX9FC
nzO5cYrNTDVzXCwGij4/Oxb3D8CatwcsZjQ/2iLx+ad8HMxWNCDI38BrOHD3a3zogS+Obt1/319t
f0BC9xj6zRcqPPSXRJtljztTDMppSz60Z3KmhH+ZWslIXnpWxsJPBHYji4ObphtsbBQ58DjHOf3Q
mLnS+NfJ6IX2DKBUuD3K9NxA+yJjykken81rgcLlcTYz0x+qcRrmJVeHxenOGg+1j3wnliZ+Orzc
ZJ6DpDKhklg0hyA0CSolq5ihuqAMBqKRSJzuCcLuPPw5wEkDllIhkh79lSJ85nW4tjlvdnFgwIZF
qWZC3uLxFmiUOT/LVU51RIw/9VSaCgXwybHeaUIhhSrNpF2C/v4ZC/DHq3sqZOGFLSLnS51HhCMn
kVD0BeOYE5pc7tLd16eKkySUtwIOMhybd22dkW/o6gEFmcqPbmARas+Rtr9dt+nXP3tTOAAZwhgP
gtuAh9keWcZZV4Lp0DnIUCkgpI4sBlcQYDy4aYwzvZVdAaQMJOxFbRGzHbsljYddA9P7x/ta6ddL
v6owCQmSk72cxvbOBw1IrfT3na9ut5jZ8IKJz149mQJPc7qeMKrIT5VkMkQ8N5urKhlRoxhaZ+WJ
TBVDzQLI6mmNCZplqYHyKR7e6eV6KEinbF2zSRiiPmmiAH2uj+zBC5YksHt6SML1GkGpni9k+bbv
9Uxr4emy+KbCcbTEp3AQpJ7l3MCdfN5XOmlv7f5KonOmqoTKyr9HL1hpSQCbYLneIHa+4dOJ+8M2
RWDZ69f57xAOSoQJg9tBeac75du3DzW5a8DnttuJBjLOsw37nqwfO2x9rhDMf0T/xSqBJ9Vi42xJ
UFszBvQwtx7atWG0I2byZsHA9SS9omkYAEh4bWDr51CWRVPA9h6gIFQuUIodryKuJbdyZAZU7Uvd
WaPRfIjnbchN858hjwwlySsu4NeakQi/Uj4AuYrcnVb/8yQkRZjB4EnPeTRiJwVGLYal9OpBLn4V
cTDeQYBVqoKATpqPuswJzywhd+ZRKiIJT5KhYzBeIoIyMzIBr5KBq/uycKzqNyFOpNk4X+rPPKeR
7RYYegNDRRS1MSliz6WvmdSQCmxEm8VQ/QnlbXK+emh2RGMr8fNOt2Siyb6dD3l54CsRvyF3CBKx
k+bhNVphB7HES7JREn+stwCxmzJbhh/GKG7Y2jVf91iaIEWbXUhfVOfwd2bCi08GAsCHe6pJwBJb
MtBV72wVXa7LZ4Odn3T0C41E+brOZCl4+chy0NnThb1OdUWu1fNImVAPXm5kBarkD5uqWhiDZ40O
hmkXTRciIQ42gIH4Kc2aZk2FMhrWqY26Hl0cMgJSl+JJ91BlQFtHwul7zg0rp7fnJP70miD2AMj2
D2ICfBJxMTgUZZ8t4RERlbqLbnt4afXA738u7MQiu0c4iOU1C3ILeevdR42pyme1E39/eDv8Hmpr
rvRneap4tY55UFCSL2q0UF4QedRXnONhjTv8ctL1LBYkTM8/NbKRCOg9OzlGzmeSuIvfTPEGQ390
avuLIPhpclTMtt3o7g1piFw+DFLclqoJFFO1ZWnLOg14IoDx01C7d3/kyVXJaCAvuT9cqsVWNnpn
PVHSZFXbbpMSK/lMLM8QFxxTXT6vGyv/gxuS8/jdM/1mIp/A/mSbicE+9v6bWsVu0VW6b7pzkpoz
FQosCkvw1E26h+7UiwPoc47/6fp7dJn5QFhvPJYRPyZxBvzCC/bYSO+xNhkcg05JLsVGmJUZSKJs
P2jUGDXzC+8MDxLe3OB1IXLZouTXxnwEbzlf2Y7IOafsUFyLtou/ZsbA3rr3/BkJyCi/u12ahS/G
yxJsd760ExwPKq9hufk7Ig8QfI0f8DC6du5KWSC6nsKdzyQHq/yTFXqHu7ilP+gqkqGZ5G7COmA0
jCjir3yGHzdk8IAyFDNVZt1Hyj+WD7kMbGRXHc2i8thrRYLQaeZGClx9tLqsT9CUC6Vs9kv+8OM7
gDGJ7iI+i5U970D0vF8kN1t5V2E/tZZ9a+UrWRCE/MH+MQolo+/hKw5/NQMDIR8SjOKypGHb73PI
d9kVXpRizFvf2DcGHQR/OLwGAWETwgMuQBB5G2JZovbnaW3WAu8Jzn/yjbOtpB+ipHD9ax3kvaNd
xqP0pknbU12uQb5C7tsX3ucGGyziA5LXU31PmKWTHDBKGBSTQoTfQGk67ibW69kWDT37U3rfVKq2
IuBHb/LVwkNrwGEGvDnFmv59ZNGGPlCdNgAulDSuLTAARDk+ASCwbhG7/ylFPJ4OGWeipw3imiWb
N9X16HkZLN0hOZkEUhEWsOXGqiYiqDv+zqzgVksivjUyeSFH3l+cV8HZ33r5ZHJbGQYrMdoVt74q
uC/+qrOfX7AeFX7JJhO9UuhgsDoQ5xnwHerKpF+IOI9RxJafumtVwY/VFRir9ZB0Jm5Kz5fdrbdh
1TpChi01rFogcbLl56uNGnXhKiCFQbW0MxnJjauXz9SDhSUaRv2QaYZ0rjtIRtdvEmuCE+VfLv3w
Xx4z9V5QN7Yt9zXR+pwsW+STivrintBIk1b9QUi2NbchaiMP/GL3NfXfiawpKtMIG+O02PWvhONc
lpEyGOdOOn9QxRDKhcVyKIRj4010MO7VQJ6UOk892gZX+CBSaI4uqcFgU9eHGkghXsFBD0EUOClp
95dl5KmafNiXrii3cR7jB+Ppems5xbC1WXIJAb7wVM0k+K/WKnpyoiWudKBTMhgZMPQMOqbX1Sn2
iRHrWgMODNlX+abIsxxdreWPY4rtVcSEU7qdkDufC+XdoBmp/N7rJ3sbumfGLUeKXFkkqw6Cki8X
2Qj6Yr9jGitGWKR000FSvmaGq1cVGXLMn5m8/WKDS2DFK5cj1lbHPFRIRvzhWFDTyKQsWRvYWTsF
sIhjkERX2MqPFY+PLkAQuXnw6KALT/dbr3Jgewn0Ybckd5TCqE6rr+q0XyyUv75WYDl7DzDP9+k1
4oYJVbbXnf8SRLTEhM61Nf7whFkOr5+dPEK9t/5X1e/ntQ4BfiOJzXaue3wT7we2vazZwnHcgZFn
LAy7fIE6gllTVSPq1nAwvgc9/rIUoZiIln6JtuBtHnbUv9RdTClzQZK93visUi56e/bKwjvBdhzE
WpDvuIQt4zoaCNqHyxLYMs1bks9jE9e/KVm/cZB/1dH2CApS+ZHaqQQqvoB3MFLGXFkVGsmuvCjz
x3zkW5NM8RrAyxR6goc4kwohtvPZyocn99ULg+MGFu/KfHKJSLK6mG7/UBwLG66Y6QtMhd/rlIgG
VSV+PTQZnzYtjqwem5LSf5oa9mbroy+0EslnW6cewMJDpxWiQU8UPdhqGOAFBiOdSJXovszm/IwN
D/eHNxuFRlVsJpMSiOLPbb5bpVeBga0qZ5Wu/ZLVy89Cimbgn1yZPAtBs9dnykKO8O2l+STUtpCi
Az3GW1mK39t4iKARXL40/6zqLXuzQHT/ZAjuWr0m5MiJfvGxmo3TTrc8eMvLZa45W6WmJ/+XPk7P
ra4Ow9BmicOgxrZZZUY9gxYVPq1yTk0pY54J6NSVa97PSCYUrobqRqdA8TEiIo9D3sC12XikpYw4
jHND2UGCkj5ccndpyykx/JDqQMF3OCQ3kDI+xc/0iBGNxpcfJ3mc9gHyCHZFW2jsn53uj1WrZwSc
qpFezrrwK5W/SAfzcVPKRQ5izTKkcMCIwdfXHX27Cym8s5RNPGY1AO6dG4/xYgzKvP6IhcgnYeaw
q9u3ifOCz17fyLRFqWPTBtN+r4v+7VSCc4VGIXDgPh5JZNH4+3bjTkIVGVZPtybF1kVbWZOr0kRV
a/Ozn7RIAUjOfgoee65SL4ZAOhqTxUWgDRZhqCXT3WVIexAq2HgGh4MQGhTwTryXxunll9u2ulBD
gQcv5nUbitHOrTBANlDfQF3907CLAyS5lRM55A+4pgxDcE79efMeBKAuAAsaZ7sjIjbOnVb7yzJj
XeTXy8oQrxDhMgRYKtL6p5uQFNF0BFdAwmaT+09QDNyxl2rtNRjJY5jGk7ldtw1TDLoAx0tUVY/S
4sIKePRuZwZQnhS7EIvslicP2vQF96y/puu3TNayAdPdyEEkkYzXWkcgkF3+yX3NONkToqbEmm4X
0SbbNM02erQDiJ6O8De23icwnyHnu1H8qSRKtqmdiPQ+JY502eod3rMf3SJjkrieyjrgW39U1Ag/
51Di9oou89D/Uz5U2oqTjcEiEqxcNOdYyFyKo0cXsSqHjRayIPdYSuW4NOwpxpZha0IPFFTsV3tQ
JZUBO5VK0O6vgUMgvdgWxgY+ehpHN+Ay1yVBnoXdemArkkFhcnRFxSjntbykEvwNMrulsDUBmeWm
PlRR1ikBymXxifskNkRd2zFPeC7F2tXoYKKSbZJ3C3p6Twdx9n9oa81IACh/LZ+KGMpcRsFSVgFq
LBObcNsw52K/XEyhwkusoEr6rlKWd/Lqq++eh9A3XvBVywI0uK3ATn2Ig7oa/G0LhjEVMkYSFL48
/P0GZZJEeR2OTLBu/+VlNXZcyxNmzpaJWoJuuiTmvGnWVyOs4lAFgBEge74IcA2+0j7oNMVituB4
ms0YRquz4hCNKQYeoOaq/dzBpKnjh+JIzI28aMrge9xgrl+pzcrL18ZLZd9kzx4+jOQpFkCehAxC
U+hSdKbMkFRms3wYjiFY5ICTtOGfvKV7OtJCQ1J3KtDsDVfqf3QVsHBs2vZoEiE3KxhsTNllt1Ea
O+mMI6l+4Huf7Sl3j+oHoVAE+2dDLwg13+4Pe/oXHfknDayHkRmNq3ai2ABG0k3Vwrtj0sBbYUrt
zg/U2CFUIfeCEweqTEOuq+Nm6I02BvYtmwKNYkQNTTtamw968Pq3hYwAnX4opJMyBEzNGEV8DWeP
1igYZxMbTP82Zge7eL6mDMKpOVlGByJx+gYZYaFqaPwcEWUqo/b+Uk+VHskFiXB70JPpPS3f3suu
idhsgM+cGbWzpZoFWzxXNGg4azTb4Zu90EMr+BW2qeFKqV2sD+OGctxRO9xgELeGVXZcgPTbft/0
57Kerhf6gsVz5H0ao0DShboAui9th/A8xmmYqIsUlRQQMZUdKfSBjvRJfah6er2+kFBuiOyw+YAH
Q4gdmqnv4SKtU5dijX0VqCFJ3z2ZD8SOylXL2hS2vOf3kh+FHwh5sEZLLICIJhLukor6QeAS+UIU
VFriJbyHC3f/PCQN1AsyVUiBc5nVobuySMJpo7bI1yIC7ASK9ZgG69i3giCDa00vV5l63DDLQg20
VEzzD5GUppVjV9o1bb9yvbJvwyxpDZ42jrtNxjkMNzRB9SFm636JVg5QNHp3EjHlWFBAKEF/TEuQ
5CZkMqor9baY3TmLEo1wtREpP0ilPr/zQf7hVRHAY/KHLqwACZLsdz3w2nUxqcVD9ZXKt3Lro19r
CrM2dTd0izCVIa1CV0yIvukWdz9QqPlU93rzQ2gzLJX+utEDsv+J8N4ho5G3QHh9L2fPAhfALVme
7RcgA7PkgG6WsyB/TWQuWgo6D9F/sjhKf41vcaRkKPXayzrijBA/SaIXKTGCY25szSwkzWtfOYGs
Ht5KKwDcAXLLeS4bXy7GooSdGaKwIQEqPvIcTnhhC7gDGhapZPrL/OV7/++JEMHf+qjlnTYQkY+Q
zhYFRweqlJpqkb7UCxG/gz3ax+a2Ebjgz0Fnk3vo3xdHzZpeagq48FAGxR9bNL67EGsCAsBF0qWi
My6eVgy3fDrZSOz+VbskN6py+OE3MJMHTPnh/E2vDCVUcqNQ0bKlAQGyTIKZrf+NkGlTAfKeXpRS
BS7VdWSOEUTx4V2DhHPHt82QVFGj7t7gibu9bwzjOpDogfp/L2PX2iAjRjv1Jz/W0/RleDcKZ67Q
XoIFFR6fT5wiNyTiAM7XCwXNmh2nTrDOC4h3GhM7JU0gKRUSrZRmSkKL+QJGTuNE2UQCeLUULHXh
dzhgKDyQteYh+RPTHfAOIr+8NGnk55OJrSZ6dLHh2sciD9LcN3dLZ3HN7jpRsUhAfQPhm339sW1s
C7hfHCZsfrEu9KV4BCNxeaWoR2NX5Xt+N4vJDSjrnsr364ztDYbxigkyIzV4ZnM2ZRd/bJlAqKP1
MwGjySS8Wmo7Atk8AyjcmbTOzDMxlWRu3lmV97D3AdFR+yLFhVnEqbHWbPiBiLYVAOOyq0Kz/+oF
zh1s7iAlDGG0fVC5HuRp0ZOj36caHoGp0szyb0O08nDt6yGymo2YG9QkwPi3ocTOX+XLHTRqRFNy
dxPypYaSp8LndZ18Gf3cKxt9U65ypovDV4bpxjZWxesgKZEPK0sbpCtkUklSzqCJKBa+Q//NXXlY
v9Uu3ai24/0S1IR0IPGW59LwafTlGAyVBtjkulLDLtdfCguoJyijy34IkgHyDLdMHxYujNq21hb2
1wooeue34Mka5vYNTsQ1ExTESp7SEgil94Q3FDhTw/r+w2qhV5o5nLjTPaPCpBEBOeLXsmFdHt3n
F3ZFGeKvu0rwRaCfBxZIZ5yXrvMGXqC6O2aAeQAgWDLDDqF9oEadjw42ErfGP0WgOAASfTHf+2MA
rod1WEZsXn1ZvqrkPKGVervUdANZuN7wdYBsNEKkNKMdR993dESSbz8OFZSwxc+dReoamMIiOyqZ
5zJEU2NB8Gp1jPEGjbwoXkMq+X5IlCNGJ9nYebeJVGplRJgzmFl1zzGXmEY3yA5ikwZ2kN0vwura
C+UDICnX4SAgrAO0cSm8w3tcrRQG7Zz35LxK/V3xDQjT5dOfhxX689mM65bQKsO7m+iTFBWPMYfl
rohj2DblmHb3+OwmeN/f62XVGC6khcXSdJwy/PCAaph9QCgrRdOjbD6Be4yg/g+Ejzm9fhbAcp2+
nMJrv7Ww/dkfqEnoVW6Zk5MJQ/9FEqjSsEs/8vgo3ueyOnRfnWL9aoX4TyH8/6uofKGQBJxEWqGv
gTmsLuOy3QeJXcgA6jhYcThSo/OgnLgABXy/q0Cprpzlv3RRz+NnDZ9w+byqRTvv4Ry446oLq4GC
c987BTb1DSRT2WBxOeqlzmVlMtI3p5GzhzSiK2tUJGvVnlDTayfsNMBjOwxpbz914ze/EVMPotRm
V3z4FZ8tO6l4wVeRRlgRlvbRlDdXef0aJk37rtKfXHMIjBBoWVBuamwgcLTMWcYu9bKdVETM2rjg
aoGN9GgwQ1aDoEJaVUILP+V6WvXjMO8eD/zXX0cGtCfHTw2LwgEEceRpNuW1riRCKCRRH7o1HWml
WO5n8xpw5AB75sAW37KcFWfSxQwRir9+A6zZryokpuummPpnTwdg+aYXVHqRSAwooFt5dGVwRZEr
rxP0vzxMUXdrxUlvJ/RLa5/osPqIsPIsWflEon9QsGEfGsom/O+BeQWdCfHNhFKPIBT9tMQ+RJq3
fUm6pKBNOw0DEnhJy3Mcn19Wbfuo29pmA8mIhMfUGcDidiQbgjfRFTyyQEBsba3xfVoPtWAkkLEf
D/XnPElDjvSaI9AYGcSEM9OP0ePPvPfVRbW64YMgVVstkCzFJCHn4Y5SgSbSJzQN7rFOCm21qEdP
lLx7hB1NXvVUTOJPWhmgBSCZoJBbGj5efWlPOzQR5MNlXSGVihjlblt5HhimE7fO040TxH8OLF2b
oiXuNQW0Mi9+k0CRgKBgiu97cdfdF5Py3lq/tizv+RcAswBJQ/a0jkophNqSFmTp+nsiytdZ4VRP
DxJbkj0LMKZV7AfpL2AaP5R0p+2JhMFBzlYP5prEz7qdgxRMEXpdLvFInCgaJyCCVryjlAGC+Zpu
0azNFiqbUU+f8+PLFUjTaOrpipZE8JXEP0O1qAoaaEWlPW9TIFPV+Xa/k2rRE2tvavNqXPAjQtrw
JBLM2v7UzxXvP18ordHrJ3BW4dMj2d2BKByvm1O1QhUkPL75A+CVS66ue+Or5fbFgo/i2DkeiWpN
m/md3c2OAUsA7hE7xvi9ac7cykVqGPfpmaq6OSaRiH8q1Ny7TueasDebHSwudrUZqjieAgd+epVm
9Vhfnt4C5qTZOwOgg3pnz8u5+3WmJGzV6AqZ2BRWdIn8M1TGL53B4sFaY6COH+0Ij/Gn/+qQohad
mdh62CQOm2aBcQKwa1jIi42DiZIx0FfVeRwYYI/N015pihczqGHQUu1cc/DoLbjrSDVc6AZbNfE1
7FlA/7+PsYCViRdD7VSkiDLjLcCyKbkdLqDF9Ouu94vTEgd8YKHKm9mfvsO8eRPa4FCyhful32Hp
z2/l3K1jQeN3KT6upybyvU+i0u10izy3uKpJqDXZZaMymBsGKLOC2RgqYBs2cSdUaTw7rGHv7oK+
pUax9lmoIjoDMvB7Ad5tPyIDc7DktkGjDtFaRVWqnIQHsE0qAaGde9yVcyrOCq8QR8a/jzNtJVgm
0xTfGbs/eGXJjq4Wg0qEN+xoOQKpJJoLUrAWfy/4Z/PnqJdW95OFQfHLONvEacdp+27w7PlNl5yH
ZFUjaedwWQ09YJWAh2SZwmo3aQDzwHRLGcKBEtTe7fxEQ4btZuX1HlHphXapwne18BELKroZaxIW
cT83LD3bu3YS274wrOsd8IIAKozkmm7HGlnnSXKPhhMzOqn/cRn7c1kTqSdFse6RLyLY4vGkBaXI
/Wo2soAfPP3dU6Ee7vwjJKW2PFEDluizqeVt08jqy8u1ki88ssVAkSbt4K09xbjMRyWsMSUDzvAZ
hLgOtEaF1YSCZXFNtS3BGM5cSZ60vAGA2Y+iLqee/zZ1w5j+Z7HVRsDkesNNczhCQ2Rq2mV0ZX8N
vfNjq0mhKfRY3+MxUJdcZDsC8OQraYjBSE1aAmiFB1fWt+Txp8t9o1ZkROi0/aZfChC3wCTg2hgT
qUg4k39o7YUj/j227R8J9LiuMK3nlaAqLDud/CSduFidP1FOjQYGjlwkXA9Pn58z9FZ+B/GA5twh
k6C4sG+RU3MCaXbDAEi8coUZwF+8vWWaaKhflEux4sTjuhwJYxyxntwLxhuR95FwBjjh/w0xxRM/
8v7dBBfJAfehCZ8JSIGw2uHm+3vssh8zsbtcxyVBRN6TkpW5ox/3oU8Sx9tvnzLB3BiqTxdgrwcU
389YGELJLVybtxwEgXsEYs4Gj4IQ+RwO5iQxC6XpkKGleiT0RYM2FWlADJtsn8MDrZ2ixf2P91wc
vqfeUKy7CG66kIJhim3S2gSNaCXEkiEhiyVu6rLedrNmSWbXlLtZ3PeLouvUZu+CVDLoAsYx0Url
6X9haKHsOLvSLvt4G5kIlwrn8QDapPfESmJ1y41y+lp5xusr7PbtRK6VeMEbqZUIDMmKBrSWwLvB
8lYNnhB+M03RRiW9YEYCYNj7YVGhJdQI+rcGq41SAoe2QSzMhy1VuHH4muN7yS0wjqPAj7EhHeTj
Gl7XY6mVM88aXa7YKQovbmcm2W+q2lzRXjwDmfFn4Mgl5VzhZOlcsD3NMJprbrgFTu6PtgRmzMSl
3ayKKeZXcgh7reD4halkOGgWc0FfxQgr77Qri7jl3zb7npWQLcZ4Slat+4blqdASgSs43Af3fTRZ
tqsIWVkdDUPesnUI8ZFAeHR+pZ+am3HqPHFhehEKEjy3Y/w4lcO2aaDFAP3Y/CeWalxpx3So9sPY
iuv8Ik7Hn7qVSv2uwt3mVSSR8NcBM908Rt/jIpNwMaGqtYGFcDXY5bGVebogd32m+pes3Bty59si
hhTJ1KCxKLNjf8d0dxpn4y44sGIZoyNbCbp6ALIj1/qJmyZaCNlxk6SIue1P9p0SzYS/40zssxpJ
CgK7y8yxmk/lXczorDvKm6beDtkV2k+fXazFa2CCY51xFQB/+Jt4X7c7XWJjnY5GBc3R8amW/VJQ
b3Qcx7IiM90sPtjxfeyJqxQ6bkhdVUEPTT+fkmb8egYMFLi19Hd0Jwx7ftO3eIG8eGIqUMDDrfIE
DIGKaKJaHuzxOeZFE0NHzrxqEB9N6kicfpefdf0tNYqGkz+6PHr7t++3kFIa+x58wPzCxp07fT14
Iu4MLQcvVX9YDJGYq+Aqk+skcOKc6l3Q7270NDCxc/xYDRJX3FANNSrvaZHSlRNBt2QwYdrCXpt3
2JI0Ml18q+b0gQNsdyzQXpKxxYwaQMlEqrxHjXsa9+1l2YHCGqdpbRcbvGYcTHGmDkCq1SJMHOZg
wegJqsJ/1PXuPZJW7Lgy7vQUYn9yNISLlLmYcr5/jtuswb/d7tGenbjxJe9Q5hT/sP3CAwPhdBI3
zwMNGtj9R+VpMat5xCZmvIPfhq1TD2v9CNeHH3VIdNvWda+6gdWVLv/DfZ+N6y9lgedonJd86rRE
HuvDnueVWFF6DhxaXWutGIdOpCgZiwMzINCI/c1PpIEwdY8Sayi3dYO7ibx+WUvR7nBAC6udFFWt
mnKmIX08OoglFW3heGkd9zRBeKIkZQfn5e3Jk4/DtFRI7TJsggo1rPI9/zyqMhfP6/Fst0oXOETP
D/HAHqzfnppeKr+KpNcKSIKRYSHCxI01hR9NBh1YLANPlP7ZBuL8kcfFfUWaxw4RUzvm6DoiSqGH
LREoOhDOH81L/RjBrj6/KD6cnzMjgL5PGX5f6EodEpZgELKPaCKFZfOrTR1SxM2pt/vcYAkJzv0L
NTwdPAuYgtc30RBhvhAvNgCQfHR4mw7Y2u19oorNka+p1PSdVsgWNh/P1aSuNOin9hS45FrHXaXr
fycIFFKQwp70scoBlvJGLxZzYdEYMmCAHMi5/ub0nn4L0rj7caoSbKCMdf/0J+BczbkrhI/7rG+B
62tNHrieCYgWtv7P7RP7zALW63dhFAyu1RbTfPR3C3N7OrnHoWgULB27xLQL83ID1CTDXawZPN7R
YQDgWZRJ3quFkmDOqqx6TFg+E8nLDmH8Jd/P/4IpfqT92WOkme1DnVvNReO98De1tpyZH+pCNfSx
9p6SoPxm2KkmxbtfJgdC3+cVd8XY/d0uWD/6dpGUDkhbMa56KgN8mEtCJfEKvsMBClwzn4WA8YVh
2TbgPBhSSRyaShOwx0OGDxWNv3kC6HL8j/TB3csMyngWqYBrROPhal/gvifY6EPvtnVIp2Om4vBT
d1cJx3KngYKoXoYl9rn5ZZOM9SjE34j2g3D8FY2eUmYv3rZcdL1bHrgOKO62E7zk7+um7i7jEos4
bo78w6xhpdcFYhlmZLFiL12H6F/mrq2gQBa2K75/gl32nny+DtTkTAakgpuqayxU6IQFPQLZiuRU
9XJYFufy6omC7XPkDCKjPjz2mygDB1USD6iJFd5nHQptdYvUL+YdWDOG4n78rbG9M8eepeBPM0VL
soWcYqy8qODqHrXYizUvEwlaxWT8t4TrflXgZbr79Us1BlYWjgqUFo15q9JDXG0wn6Bv5xvOtCnV
LYFh28gZBqAA43G31/aIcrWAq8nQEHjx/dfId013u1wk8oosWkn70WDzMa7B9OfS8249fkB/g30G
wyvSzFa44zV7gKEQmeQYOkAhMLfB+8tCVYysoM8iByRL6Vsvl4zOx1bwvAfoSonMXHjT06UO4fRh
Y5uY3McDOym1/cb53f3s/DQwc+pVTHlTRyzb+V9yk7/zhfXJFg1ZdYMkEzyaLIbZAVdWyK3YjTeE
gCvopIV1CwiuDfS1wr3BuLMEROTyiDUWasB85E/Ngjbz9uoT8j+AyvJpAuAnk/bVXLVw7vHZi4eR
z5Wi20NfhYdfOY53s0EIbpfo+PRga5uovi4hSb3xgmvdFp8FVn5z06DkP0qNBTZZJ44UYHvbL/zb
yFFbZj8MtREW5r/QGH8KuBU9RkGJDLw59PTNgrnppRctmpUPt9+2FktTrCMYrjDEjml64e8NngY+
gMlF7V3MUrxcesodS5Ti46HUlcnU+vMpRbsHbi0ktk9NZDQj3PDA0fznt/hPeuqr/G/it1O9cV9F
Qo3+ZpwgMmEfe/4E8p8hTrXlUP4Dx+yRd80n/eqyjsf/y3OgPSX7S5I4Zte97zvp5sh+MO8CoFdS
etLFGSqtjcrAo0Ju2UEWkPEPx+Tsi3Xme7dDahggK5Yg3Van2EqvswjRgTH9vD9V0vi1sUH5F+fw
mE3oGKjZ+Qfl2sq7BxUn7Xe4hJTsI+bFF+GtUUvTm7hmiZHQLdqxE49cRb61MB6sCKlR/TyEb9AW
O7Hp51OG9erykmv389waLWvMaXgm+UkY6BttpsFzrNOpd3MZUoI/o9frSimPmyyIGdVovxbZN6A9
CdDozOKNzWCoj6vUAthB8qtm+15OrlTjMAEUoJGAHuF0EmZEj1tEv2FNiIrSMQ0LaOAGER5uRA2u
e41RQqmBEFi1oCeXO06AJaGzladtbKwPARPgAFR+tRbfDFjhkhIFeJOdQsZQ9C+4kuDs7a06zNqJ
MGm65x9LGTvVN3iWwTv7WQTI2Sl+mGAUwEJuYgGJSurOIEXJ4nxssFTnwyxZfPd9XzlZSiUe7PMp
cbksuyKtRtJikXTa/hjCDTW8aTtAA48UJfJ3AdjEkkhPAGhyETHLHG5b0LPV0pg9EyAGNKrsmDwh
lGahS1bvzzfyHQLHnVpV/VM49ZXnhr70SDOTxLxK31GhnEyIIgaR2gaBRxl35fxjv8Q3nadqCmsb
oOkmBSCdZmTgXIp26oXsuCuHZoxALJ2qOgxjmPimS8EhQWJ+chOJUpRlA5bgQmZwSwHdiheUUn77
Lh2S7nsngqs0JmAYc4J3aJg5m+rCjb5oLIpXjxDEdfBC1gRpQ94Xx8DOFs8VepMO0DE8IACePsIs
QFW/qQ9PzZ1STNEU3t/vwnGYuFJ7IpJ8BYoUet2susmc5LYjMGU0iioTbW06GmLeR04c13S8vOzs
l7G8PUjWZBvQk0AcqSwInxXg13xXtNkxJJWWV7ac9erV9538OPeZ9/jroovdH2THMsrDIavsNcbC
J7IEJwyYOlEwnQJEK1mGYFMjUi3AM3dqGLcnbKxmihB8SwlTKoKB59mKyMIaQGCDb9rbreSoiwbn
aBVXX96AFYd8GMti+pFLYpOfhalwGz1rPoVQKMVbGmJ5rNdP+3lVFgOagSWClZOsB5h1yGfgvaJh
M8eqY2VTNQ9JTGFOZ2h5yAPCJ1DJNeRNSIZbwpIQ5wFH1ni9eULHUJhzM+JiIGpBnXtRK2IhRP0W
+q6E3zmuVBPGSyn3Bg+usPY0Gh8qhzxpbGKzCYEeOcT4jBhcs/PoEOowVqzDpJ4vVKu3GZg1qOrb
0VsULY2Kyz1RqT6e2eANFmYaH0pCdzIGSpQTYKFcKLHfLDFgFC0zaZHHXm7yewXTC7nEgO+6j5Hh
hatQ8OTD5B605zy97mIPZS7JR1lpRlKXSJqjfGhtFC5TKFdj+KMmGmJJiF/sO1X5KxHKg1khwUzz
n8zGFJbLmxfZ81CYneorgNht8y736FGIrLXoyc/tATIBzFS6RerLUvKOXrolqWPnn9yhi9BfO4Yg
ZuzHMVIlrQ6BXLlo+vfeQCG689rnFYCcRtJ7t4ev74wqXV7IpMg0xpbc2467abX9yrWy/3jC/QbP
Q6B62C0+xA8P2rq2ZC6X4bvUY7InmXuBcaFMZzVs9vWnFugatCy9RSsnsRwHE4npWi1iJkiu0S9w
/vcB5WRt+jcvPfwJhW3AoLXQbU2wIJVio76fjI1X7/LVRcAfv0ngcjkQEyDRdyAGjED33ItK/08E
1vsZG1ZEOrG6s3BDWk78UKhaIqi4DPrdLhmTGoIQBCX/HEVLOtU8As65OxbduXCq53SOgfgDSEFU
HKLmQqWM9d1dq8ZKz3/ppOUOnfvM0/5MfKCCcOP/QPWxBVKaNT6GjVaIhuH+T3FVotcDPboq2OG/
lHj1jjBn0eONio4w3AsKqzk6TeBEyCb3RMWh6PULo9WY+W/EHu+kki6FQqTvOffNWQi8wmRJzhNP
7gBF2KRogPDV3Y2ioz0JZItBYW3tCaQ0r3oH9JI59CV/2Z1zwyBhnS5r31h2ZbhkHSaIE2jZX5rD
of2VlfApwe1Cdsb6oFRnFI4VDUXYQpk8eNiLnrcghhxdVVEdUfWokt2XaZx+2jMsADp6Fx82CiI2
lj/Z0NFXxiTV5EOyd8QTIFKHlmFgr1HInbukF1L4Hidd5va4zGBXM+x+gkxHals6mXOBxkEo0Adm
nqqvQP4sxRW138T7lWADJUndFZVVM/yb8pn7HxVb7dRWLQq577exsnEAiGNJ849zXOFKlUn67Stm
d+/c8iI+a7cmVejKvcc6ZW2dNDuCpefPSUQHk4+0Yasqg2PXgtNep5NSm0fJXbi7i1ptqa3gkyU7
EFdpMJedKXDIHrnDfh8qFaObDEr62hdD8VC7CRO8xBYC93ZalTEXrIccAI871I0cD/SCigCjMicw
TggYl9Ya6AHhkp1JJfa0SKjTZYfOWcvjEPueqspDVqt/icg13oPr8ShTxEEXJWVq3H5eljE3hVBx
q/ZTj+Vl6hWpMwZmK8ATssI1eVvB/7WaMDu5jJz41ucdLBu4aO5MH0iTkTr871p7X3N+L1a6ythZ
fGRnneoQ6T+Rl3p4JwUB11Lzmsjk7KQDjf9v1AQAcFk8BfID0uugwKvcTbuuRFZE7efiugNz7nUw
dyposuLqk7Hp/n/eF0Fsuu33eBFwcqbLqoLZLmItUGTPHEpUzTsAaBRB0+NcwxEJ6jb5YaxhuO/6
tkxOwTu/113GvoGkPA6xj8bhgY3PaibwUx/L3KkLJbfTeHiaX7e7qAhFMcme37VXOCypw17CZKr9
z4JrM73i58z5Syem1S7w7lD/7vCBcVh6qocEDCh7LgddN9PLW0Cw5ddUO5E+Upx0/lHpGp6Rf7sR
wNExE+yxd6HDybx284h/6N17qG3dGK03JWB5wDDhyBHLWJGERO9mP0L4bG5ocAPCzBohTl0cI6ja
PRIAnzqW6e7wczA8cGccK+rglWFFSE7AAWG4db9hWFLxGUCABqcPbCiOCFN2fYoj/Dxwf6+x62fn
UCxY3C3hs9nXIlGzFIy+Dti4gkc5xmllm/aOHqUFED81/xObVXGWr72mEX8NQnYOqQlNhqvdWeHs
X61EtSTTbwvQ4g5yMvQNDxE84E2j5WYQvvDTKbRz23IJTwMDJceUMaqPH8PjjooeQ1T2XlFahHmW
Iu3AnBPLlnLlacR4sNhkRFG1uhmd00o2ClGrUry+QqhXfSPVeLXUgEmFc45q4i++acRdfTh2MNXo
SC/E/WtZJNGIq+/hI967zywTmMqxNIKglP4tzN3is+jwfxyW0NVkygwHglM2LltAyzwHRVgy049Q
nFjEEbxA01Tfi/eVkMAAWYE6JpywicZxa95yE3OtjUw/ZfqL+ZOYRngZKbQ/iwwwinUdJX7y1tRw
VwJyrEqpy4jv5VEnTI4zT2oEKW5EIqhDrLqRHHoiaoW270yXlk63SWZhHVAcnTh82FBlPhXmjTwN
vc7/pZ94NvuZEWPZF8mlCBkVQhTPllVgUgkQSYvNr9PLC4TvTY1iFjGeLDwYn6YNFTAegZk+IF1R
AMZPU7JDVZEpzQnmRjK7KvnJ/wCg6fqKhphuLTeHoKzUF6mwONyihCPqdPR6V3oWQwGmmZT9Jihj
gjYaut+8c6W7KgQtaRnD1GDpmohryXkvZuvYHAJrX70g3qid/NPjcgfewIQj8uzLt+RlHLAhK8yQ
kCO0TdPcKyYjDzqdqnZn+SUaZ4jZJhP3keOwgIDzX7mWMLq5QS0fZ93fNc5GIR90Qt7mtahav1Hj
JrZJCQC/P5zvM4GVacsL9BHxaDLKbU+8RKbes0Y6V31SWStJ0zRLoTd0huLkyuA/0afDHcZ4Nylg
juviDC06HGlf82eFUFG/Z7e2UXewWh9jmulG7N9MVhafomYeTezDsxIqOSVB3YCOMkWPNfCJ5ErX
kU0X+xHV+KsRbIfBHYz7FIoVrBG9Fs0v5BzSljcSqrDQxAgr0kAy1bTIev1H8Lsp40LpIZztz39o
H3wLBx3SAFYCVxZ06STPwxX2Y2zwFwZh9UMOfDuIZwIS25ETjNmEAVC9TJlWP9i3MHM3EkgYS/Ae
BifyZkP5Lwb6R4y15pWgOvL3ocUwIjKg2oEmneJf0A4oqWtbqf/LChcnEPGVC4Kgd6am5vU8Xf5S
v9LkqwF9D5la6/IT5Xy16va5U7Q5UCZFkI7hsvhiGK7vO+qk3G2Oa3Q4gQ2jVBYHMWpue+utdIo9
SWh9jgDXh0O13K1Fg8jL+naPJNxaa18Vwm+Xlf9JpM1APdIylwryeckC+FcgbS2QMACk05I0koW8
NaGA34u0N6HIeLyNTHz1r2ZxogvJwIZRuwc+knuPePufX1uuAW9lOhw0AnWJ48eb7YoozXXLeo4q
mU00f4m/X51LxrhvymowUAruFiG0IUzy+BPhiLQFpPQVjO97X7kLOBTvhvdYiAnGRxMNHU6irlrh
OIGemEjEWk8dI1ZWQAj8shk/zkaP2om/c9BKJ1WFYYsmg463D6CrkdbWUgIeZefVYX+AyncLKjFb
KCazXP//Hgaa+EtOvGm+K168RwTF/NXkyld7Vlg4mbriZExsOXZj40yOa/ZlU9BL3uDWsw6DDf/G
A9G6DJ5dQ0gg+xiM/2xx/iE4f9/8nDqAqroAlHzBZT8BOPMvRfjvkcCPffMEoVZkWbUC2Db+8TTY
UR9QPv83vHDWdrzFdiqWi+1E2VdX4sq5pZ7EhpzbJdlLn6zKB8lZrB6Z2334kD23jYuKaLDDVevP
0jXInDOe0Si64h2NIakIyns4Z0/UlQLO59y49Mj49OHKUR0RolqCl00NOMfgBJYrNfKZE8Ppwhkp
XLPxBtv5Vo7heq1BigR9Mq9P8zU6wqTRITnbzGnFVgP+byk1KJxBRQYuE0yGgyqyVSYj/TZt4cXT
vmWRyAIw3gMJIa/ol2k5kgnxhXeZs0FAu0DblWUElyLmYH8vIHymGe7Q/fUVZG/2qYC+TjuHRS/s
QVN9k5LwuXZFS9ny8/jgaPwQvSzgYUZ85zQoycyBLOQwu32H55LyDFWz4/3xX+m7zN2SaWaygglX
tEoUupACRYuY03j9UfRgy9JA+VSU+Hj3GiL0rpRjT9NIk24mbOIJDcthEg2VLTdk5Q43pwf/BH3Y
TFtAq6pFDkFuz5UhsGjO5/38gtlpjT6/CmLd9mDpa7FOsZI8sC129lPXLbqL8G3ntN0tr1YfwJ9Z
rD51j9KQuUQ2o/Hr0WyvnpJ54P9/NVHki+O+iANHNSZFGa910iZ6c3Vj/oyDEOw9HAkApM7BFHVS
3Z4vqGQMCPKu0HAHZU7YxBD8shxACQVzEL4lQmK8Y1bEH57nLoUIvmI1CLObXhilncWNlh3c71Cl
jlfP945JOVC2BDPIBebcVlFY2/YAvOVrLIdSoAB5QMeiw2YU9gkqTFGsAS4I3GKxBa3U0gfY8iSo
B/Sqre10dsOKXarvI0tqOI8TDIQK+AGzawh5wKg+n7MqfCTnYsOcIxbgFhRek4TkIBz6EV2Usgaj
cAnwvi6wwFuR/WH0dSb+TndoiyVqyDW9KIMJiE6arx88kVCx36gqSYUZOghqrq7EhjzAEJds746w
loEBbPnTU2J0gSyV3u01FLrweo/u7d9sLYLaslsG4CWkt5zJ73ZQx8n4EeuqWBE1YCsYFmN+TjXX
dCGe7QL2uyVMDr1lVC5hiWPyVD3Vwbj0y5gwPN6e1+Guc2mzSaV9ED1J0+CEWLn1Rvok/NyeieUm
T4rmzI+5CWP9Vq72czHjNSuR0PL/4wHQeWdFVRv7zM8dGDPvkRYHD7wFeWU8ic5qtd3KMFy/i/hC
qvbVGuOpJs8enFMS3iQqVHu3lOESXyy5IxwqOu56OGKgZiM/T8fWANwDu9rA5BzZfccVhWjqjTaC
NZr2kOlyJ3921KPvxqinH8PhvVLAyeJPaYuZpJe+FmY+7z9NVYVdhbUYD278HAj6PUWi32hNHkTx
/9Z9hbuZxaNgzamLbssu8q8RZSIaxXPBncmxxD4S6Z0UYmnqpLs1kwJzS3jFNP8hsWsAMMjm/P9S
ym/r41gsqsRXfRwEsE/oXtx/YSD4g2ST16cPxPLoUpJH27eFBQItTg4MSsJNiG5br5JNRudh9ZbE
Ts6QUryb/GUpsXIR1QjYAS/A0m3KENmhR9xX/IeqWpn9iqR2kFaguo/GcZ+FEXoxSdZsriTtmVxu
6wJi76l45Nhzv96RkrMUgKQlPN80r0fBxwflXHVVsp+4zXHPRRQvVtFs1JH4cyeghV5dRGE5CWSN
F6zbYGgHCmuweYElVdzxxlRhnJmvOz78BzOk+3ESZHrpO0U1XCEY8taj5vP3Oh2u+j4Mr4PZoKnq
B96HqbF6E6PG7QFbj+EgItXfgbmqv4Q4lZYTlLAy3LIoMYMWACwcyR/Va/gzaKIn89I6mx2lYsXn
ZKldaFtoGGiu+K4XgE880lt49Slbf3/oW2mikRYujSCv9g/nTOQdzLR5skUsk6hVnnWryf2vu1Jq
lwwQJQRXIUHMePxDfdglY373q7ag9Jh8moAl03KPkHIy2i+XfRv7Gy33AbEAmaWMN9T7yKpObT55
LU1AB5doDtYQ9VfOPmi0JGfJ+/Ci046BXJPEN8Hh3JxNLidKNvfrA1AQ+ps9TQpPFfCqtPDyG3iS
+13howuodhaeKmar8+fX0oDf01SBt+qAD71niYMo7fU02X+3X6ifzX2Cz/03kl+oghGCYMNdOrxy
NsKY++9lK6sGDxzq5INSlVxvsySfCxEGZLs4HsHOmKM6YCtWHvhbDjwhI7Cqvy36uS/z+69CNrr4
tXDksbgGtgyWwzfqIqw7bgOsNo2Zhl02c91305ZHSQ3GA9BFilDfnOpYlWc1Xv3wg8zUe0osCwkI
aZxEASMSqtZkbfWrdrhcDF0EnSOAKBqdwgU8877ssmC1l3BMFTUdLLhRiProg9H7YKgyATdvihLi
GTn6oJfUzfYU3EhHPKQlecxLu6nNum61S4uoxGjtJiI0OHFTMkI2qFtBa55YqNDyOz55wZmww8Rn
LvDxLSYT7FUhXAWSmYBOf8a1fCAmg5sf+cXJrsoyCwnZRDT17UW32OMP05c0O97mOgFnuNoTIyPx
uRFy194s5BVTuV3FZwdgcAzcwQsrBTqH8+Fogo9LtFY9j2ocNRqWnTYjTc5FiDIQ0rQ+LO7gBOnn
jEzLv7QyB9ZTU/v5XeA2Ijg+b6jCon4Aj/JKZkPUKr/H78SBk/liTEYCm0piVnAS00d+DFjXMnCp
BqCiCt5beVvCrIYP102WM+07GUrQA+4l02pL1IflKY+PKtVXL5jHEC5MBLGfdl7D69JxMW2v4hgd
NVvL5qIXkzjfMXOmHMGWsqleoLVE2T/+Eb0CAuDbQrffMOBjk/wCnvdIG/BiZGTpv2N7Yd0VRkhj
/vToSNtMdl5Y8DXiU+jtqth9CM9q3M+8AIwADXSKZMNmtk0SyK9rWqbSlcZkooyzj9WUfZR5RzHJ
5ViZ0dxowtimukYGRm6UghScQVIoGWc6bdB6LGefC6xP94+pMYjdhcTiNABqJMoMhY4uHRpoRqbw
opLVk6xwyF/pnxdd3vMFFGN+xB57cTeQZ6QBm7osv8yc65Ef3KS+ggH5JQ9yjPEJ8DpdF6LTHm1h
nijZP8RhUi6wIMCLWJ8XT1/ZoDvlDamX2l7GXQEMFQPwk2rrvF/n6AA3ppIn9s8t5uM8IZ0JUzMJ
78F1j6Rtzso+OfN0oX0A0vytk1AYYCVSXmHtB/PiuMqtVwsNkUFlw/PEbiKl4vRpVV9PdlwIlNbL
XTqDTs2Bybq4scOOZQ1D7Zal6ScHIRUZ0cLN+TrzjosqTypIKxK3lsdg+AeWSMZolrn0k2UiF6e8
MamM9v7el9LQe/n7XWw2in3JC5zhwXGar+VQv1SKoSxBtCnZhIR1fJC3vEDgfVIuBcaoFjAoh10L
QgANLfP5kFnBRc2Xs2JZgw3j5pNOMqtf1Q0aw1TiTxTkgOuLCWhLJR5k1uA7JYbZjtXnvo6vDPzL
pNazN+ZZqMPBxDtiQCPTVYT7V3UrmreEPI1ZWIiIcaF595oEOQj0ltk0doKYyqCAcg1IWTgkKkXi
lkoHk1Qx2nlwjwT9wRxoadcXuI++5cVCNnidcEamIn9Y+Dta+XCMCe7BUpg/obj42+plUAj6n9qG
g2hWnvM6alohZ7vtMxmRCzDx8PlEyzBeczWkxQm6dO5KHiAAxwDLl3jQW+bfDzdmI5Kw0ETr7xkH
R1+NjZmAS5LL1qlOUnBCC0kLwG7iSFBGrSKBBTh3AbwBAEmtryRxEOYOy2yJZFXaCMKpcnxMSKXI
EavCSvXv7VPOLMpIM25eITvCKYvQI6WaS0utggbaLKB4E2hoDsf2/VvqOLdPfSJG0Bj+j7seSWFa
PacGJjtQ867PqofV2rNwbCGZb87T+rmh3Di9bK9GDGqi4MOOEa1SZw55vozdNUd0SDflWKM/MwWK
88xAptbG/Eu7/BDeZUM0LbESKB9F1eKvGiCpLqCXZV0jTunnqRNcvfTF91WJ8Qw8HWO7a2DIIpvf
BCDbU+OEbqu/hKZFD+s7VVm2a+mJ5UYs72jxADJmoDmm9XcaY+ttQdxYkDSKH+3dLrRbNt00HxW2
Cc7TzrUnKoCldJwF0+CGaIJYltURwRwgw7vlOQxmWo/hxcXeOqEm3+rw7AHzou22/c61aLTxcs+k
0y73a4pzDvOCADTKiQiISznY3u2hvauayHynZkR9r8N4r1wBzqGxd6tc8VTDzHUVz79ttkL4WHDp
vOH2QqOF3SHwsnb66fdT0edrvxrRL5WPOAOv3coITaU0QeQcw4UduwOQq93Kt1MULN5ABvmGrq0P
C1WTFRUttJ26aZKlN/nTrplAoP8pREprM333C6VRwj6Y4qKvrbWb24pRv1J8Yu+3uRNABMc4DP1O
bOiwBEYlpAaIVUtA6X+aCJo8MFCOEZBuTI2YuqaXNqxi0c6LeJrifiLWCsnG5M0L2tB9mYJDC+cP
yxa4Lw+wX5G8FdlrMlcOWadKDLKCVqKiwiKxgckqGJuUNOZgiq1byxqNlIilDzZBqqpSPcPBLC8b
7afnMexkwHz5G80xJoRMKDkCsxZeSsp7v3hRNQBtIb8TLY+5E3RBAJ7RmETgMe8Q94LOGQTMz22f
OnyRy8QYHsfxLm1ehpqD0iTotNy2htaBgUS9nRLSTt3oVqyoUZ0LxHNFMSUOexu92YeRhUzhjiZ2
tFUsjT+TANmCgSbYg4xAG5WJO7mmoyFtUcfeObBJTQyh231puIGdtHXbt101s+W+x4VCgEiMIzKw
5vdbM1Nqay1s1IlVYD5JfFnYbpXy4GTrl5MurqxUseU6RQ5uEg+hlBtR/Q2/lJH8a4blMSM7hb7r
aFOztko8e9a0n0+TY6osOzM4nG813xc9Nm7m59dF7+6OL5KGl0HNNTepb3q8QV57NbZ2pvi2zPfx
kPTMY4cS+hCBs1QM/ofuq+oyTLKy9uQuWzyoXEVyB67mgUI4pMnXqd4pGSi4FADUNzH5xbTAas6s
LeYkFa38E72DZyjHHUp9nI33uckj76MCIE02ibBw6QPo/CNnzPAZeexlLKb4fphmGmjZeKT+b2vS
FS2t8XXH7UNRBdmgV5bFXUr26ja4PhqdXWJtqJpygWJuHVbzc5ftqU/sqM6zq117D+ZuXxIuQxBX
AVDj2tGvwO3eb3ygeAR7FCKzstL7+G/mwAWfe27PmcZsVHxQizXszDRsETbjaBnGcOq53jG15DFZ
qGdFKgXy/PfK9mZ/sQHKbo09sQwZomaoNe8fYanqMG+Zv/0cYQ1AOWYAEmhLdAoK8vJnZBxKjs2M
EWe/62k1aPdRKy2CurZ6JPY1Jurvp1HYh7L+HIwP5YyBm8GYsOCFr1TU3H4XFiBFBY91FFU8aTsI
+GaoxN6dSjWAzQ4vECto/E4NVG5O8BlBppLfEJt6N+M9zGQPUmQ+i042u2qpizFgKN+9jksXcSX+
A4NQVHSXmqBgdo6jusNoAYbUJ2EYz35PPx2yXuC+PzZE3eXdXKiqrT46XsCWD7SjpueIUqR+vXxA
6piXPI/p53CvaQsRosuH9HXhS1RrQZ/zDV7wZjuTgcNQGuvt4JPWm2GIz47zUA5zrQ7TgpcBOLpk
FEnii48dIhgySCirPP95oQMAVwcVOA1Z1lq6jvnGA8wsxp61dHwO+AK/EsMLvW0gnRqzXnUYKE16
5iVdQiwPaMbjm23HmRIkLAGGUqRixyyfVi94YJkzXcEWbsasYcuq3agqWv4wZT6avlr/Hndmefb2
NiAVYeJ4jw1P7/V7XeUx1azqRByf/gcKn0TP2tPzWejMGWDlnOv4WETUYNE+UbIHQd71WEK3pXGv
CfjHzWJjWrbkMnO7teWWuKM6n1lZE5OnSzPE5a2lNdLRAWGowYAhBWWaVZFZEF+GLf/q8ZwQeInf
bexxMdrHQ9TnfSCUsJLd436wxG/N1JFqEPWOWe4WpX9HD3cc1ai0KZ1ryWin77V02qdhOv51qftf
M5pmvzAyZA6PMPa3OW0Sd/ilveMAV5VThrOS9PMLVXjSS0IxkS4sy7m0weXiXQXqJihqOQC22iLW
KTWrGO0HrYFzsGSJ6t10Gy8Vc5KlBUr8ZElwjQmPhkoysxAbHIH006G2V5SuT/LpiBAobc7wdnc7
ZHu9Yj8KFRIolSE6YWUFa42eZoFjt3s7CjTD9VMQr7jwvXCCO4FfijzcH4xeggy6Wk+dB073Qs5T
I37LEnqY2LrSLXdYFHiyQH7MXFjNaODLsHKLyK0h+XupeVcy4dVuC3CqUU50um8yrzT+M3Y4A7iW
9Y3d+U+xO0QkkEg99zZG6vIOpb7T7c4fh+7GQBAp1elQMoj0Fbf0DZtLRKQSgLaJBMlQ7AEAGRGi
f0Tt9wGusUmjInMtPzqkPg9+tdRaN1yxGcz/48MJ+qPruAoGwf3li+is5dgX4hQ7P59RsBIvJjvG
mNwpUc/CHy1QWr5xHk/rSGrU1vp123vNrW2/D+rAMvWRwEu0nYO4j3ridshAPaqWKZKglPCH76/B
FZJ5P3Q+Lt2JD6B2eWHUgWeF48S3wZpFT+ALQqlo8u7Y2fHlaqpDolOVigAinKX4tpOoFbsNPQrh
ofpIs0jssTDjL+aSU/yFNXFTq3lgvbYTT/XV8zvy2jkwM4zUjYpOMcSojDJgF9IaFauwIxcNKNLT
RpawQz5bJu9EgtEc7DGl4zz2Avdyhft9AxzQ2V0REtwdsItyOvb0Ay4jF83XwDhc0/G9LZqxrpow
wP3EZRRDvWzM07BKfeq+PyHaSktfgiDb6J+aAisMp1hZ3yBcd3F01NpO8VcFmDE8lJuuXs5ODOxx
Vk5oOci7oks5E737ytDdBY9+YX0eQUjMOthB/EDNWngJN7Z4SD4shD7sexq/q09tCWsNc3O3jxij
2goSZdcmymbxIhYtxkDvC63Wy7wzqj3Gqne6Yt4n3xqfVOGNuu7gh2J2dCusARSuXPotOvj8gbUJ
UHbzv56af680DO07vX7zgH7811Qlqnj0zrMvxQ522fNgtvDnRVGV0KQpzIWSxT63AWYyMSdilqem
OwL83GG0GGbscH0z14gMQ6zeIVmJawsHOc+uleeW/Yx18T6KOqZyNEMcafmpjNRrlxZlb5Y3PhMo
PxwsnqqXvomXLFwa7Dw7ztqGgyH6N7rx0asz8cqETKXHPqYYD5QDNWZ7hxoz6pQG6KDH7SH3nocK
ZuGC/8KW5KeQWiyPWyNEDT4G0vFCyx1p0pP5ax1vn2itWBjuJl+D6DoIGnqUHjzrOIondhm6tYi9
U3YX5ZyYdKY6NqlBgexRLzLEa2XsYAsnq4YvD4h9vfqnCw7MPx+o8nSSiXFFYnXBDz75368YKAH6
0L5+hPaIdcW+JiN182KXeU5Dcoefga/FdkirW88TECUdSFar19d/eZsZelyWsrlK5+1EqAx9XjyH
UYjiRy9nKeZqhYyeUmPeJwXo5tOniXJtNUqX5VN4XCCNJEvCwr0P+daTnUk1UM7nWG/aKY97ztzv
yhTNSrpJfZ8t69dAjZ9Q0fxV1ajxU7JSPfwN1jKa20gamIQxBcKHkF3xuYlXloUhB152mFvmnu5r
G1t+mujaN+R6aID7CahzA58EhE5mT3xf33mIdoE8lnEEZb+jhvDu7gPTs85YAXuQdp5jFUEoqDVR
c+SVlkyMjg/4DanjlSxhMrk5CxVqrHss8c9l61M40TuDF1BfDsDs7iuS7vzABYyAIwdUh+E5St6X
QW/seAr3++K3ZePYJNzbK/biWqTSZOsYKEXotkYGrIyQKpUpQ61HP2jb4vcypdFuNq9aYC9CeOGt
jWVLS53UmUnKJYbEwNvRNjRcni6fzUoAawaZqDL1qT3J0Z/6BBlLGRIeulPED3d5WIM5oVczZ5D5
Rc4R6QEXiWBm6q1T+Gti8Tc/SD0Xe1T7CrGzNEiOo8JtExt/NonnbtIo+R2oH7yeZwtJNPgz+Aly
zIi25hZ5jnRF6QFOhztc/H/omvdtlE2JqteewBzHv/cVnE7Pdl5c7J7iCMEKDsDFWvQL2cYBVx9/
XOSWhYLXXFNxN3VUmArcAJ2IGODQTbmGKLDuajDyCjlPp6+ijJ8rsLcmHpXWYXDg8YLSzP3pbNb5
RljtVmzkvgD0dcgxtW5XPYsoMS0tJsEHGosD14RRTACCwYY9TIbk6USysys1yuDm9grPHhSF2DHq
CjpcL+lWlp//ZlZ4IGecoBaOwun54h3iclO7SJCks4wYKulDjgh7ZF9NVinSwFVDDgr2VqgQ/Cai
C8qKXALgdljJ8jKetBrFubRTK/VFlo3asOKtEzEFLcW3X2TrvZLQw8+veju3bW2oGFAuS/CVykOh
8qWxrnjUyazD31Ig+52UfcyfuHYgUVmOf78YfgDd2RHsIRo6vPgq11BXfu2IxvyrrgwgFum9UGfu
fnYzGPE67Up+1AlIRN2jKAYL3K0SmxRhB3/1pLVZvHjXGMfTigLzGmSf40grtQ/2u/xk/2Ylylo1
Vmm6FQrEoASLGdPK+3qLsyQnWJTmB2txyF3A/uyPIjo3C3V7hGK73rfCCyu7Ek2F4jDASI1LdjAI
+I1iMHVJtwuxes4jNXwpFLXAzqvyD1kPPSlMrSo90OafpRKCzYpjyE7DN10h3nMqn/q1w8lQQp6R
O09A9WadSTHrDFv3sFlQJaeQdbFJ81IFvFYVaZynuULVK0PI+E8I39akkrag/jWwfT5Gge2rIeQv
ipcZg6ZkkekCxdKK89U1X0klThT68HgmiOzhslgbiJ3B2KvToQcJzl3svEnlKMU14jiLljY3v+tL
5M4VTJWhBta/w4nA+3TPa+kNbPFKCGjRJaxQzN1zbjYvPCV+uAcNmsy26UrTumBasrw+TTC+31pt
dmxzrI05s5AkV7qfzbWE02FldMEO0K3jdJwSTnuwavgL+nNU3KN2+IAcPmbgJCf+qCjA9iQ8Ds6z
Bc7vqkqYvgmt0B6NDv0AB5/exxZ6d72Hk4zvmGOpfeyqo0Z4BcICwd0ufOObALfAJ6swuQAOfMIT
IlOpYvsKB4Vx3yY6UXfLAhIgc9o5BX9XGtIi3hEZWpstj0drtnNMxA31c5/NLLeX60wnlWeHd68T
oZR9f5+h6fipCNGwiJK98IfQ7d+kA6MLDjVAXxeqZ40DQnN3jfIcx+52mLWKMxiTtFNqz6eM90gF
OehKjInNj/+id03MbItKx9FpiFnVqaaa0hANOcYg6HLaL30YIehH7UFMh2ZbV1O3UpdMXdYpFMzJ
R8MMj3OsTVsFDuySo7LkrQjubM/oO7SCtTIJvNij9JvkcItkaOP4jbpISK3mIDMr/6g84cSk9AF4
64oixeVRPIhtGSovcVoVlhj/45HkigzOaR0eff/vPvVHJD+BheCqr9pQRJhRcbRu7ELfWiRx79pF
E8ICBjvsWrcZ6+MnTaXSKl63IhUXGipamaCXTU+9pSTjNwzZdLvWMOtEp2Zct6TlJ8bpSL0URrFn
JGM2UiJvSQCgsd8IFk0lebWUk0+07WS4Jwjv6BbT+EGv4o30S6c/+GigeAV7nkJCPzJSZ/xWQYCg
02woD1c8T/6CWoH7jtLnAeCY1yyZx/kQFrUXFSwEnaLfMAHaNR9GtEeDBE6H/8g+doaYXUg09eW3
1P7+43ZIr5vXkrG3gI79v3BeBua4AuEHRWvxe+fjaDOcAh5O9CPHfbIoIyahfwnzn2klahYjccmx
4ngSUaO7FGqQOyOv3D6eDjFeE0ftfaI8CIXu5ieLK7fJbot2V2ROwr0oCyOYuvAih37xup4T7Nsl
JvNigKgImWRE3w0Hj+xrk1LhB+TqDDd7I2sGUzOta/PeAz93Z76IeuhBaOa9xA4p6QqzDQEscNk/
FtQaQp+k1LtCnHKsUc+/nTyAzt1Jk04i3MNF6ydKoSuNvSLStPT9+EhEi7BuNSzUKkkHXmbCjmCd
AACtMLFYXdrKJ4iCxXDG7nyUKvlw+oa8FMmwhuUdLZseygRjGALOji5vBjNwFDPPMo4mk6f+LiZK
Epa/vHCbML852WONUeqN891Ct2Ld+NWTnC0SayKicKwZiSMxCVSt+Fx2x3B46pjBsrTy6ptTS0cP
H3vZe1a+mMCwKyrNYxXM4rnZkCWOe6E3eCS7ZphfmxEdUgdzjB10J8C4BENVxYZnC8BIvL6UbPsR
VJSeN56VcNgvAO9O17PIiy7CTMho0iOMzhMEczxqj3J89cSUGkgpH3dxyBg817wOaIufQbxdyshV
+AiJEdsWT3v/6kqF4XRpQNuuoPaB9+r9/S/Io2976RDio6nq5D1Ibogov6yx/zsP9WgDnwnq2fX7
BEkU8sJbByZcyS/zZh06K3lqxmGdDunCHOoQs6lQx/MV7fCF5Q1JOxyluLU8Pchk8KkiJRMAYFVR
3HvTIlett2Rye1gr6n6uxovAxz+VxGe4HjKqScaK7A+avB/za+T88y255p8GVYrTu8vld5XeyDU2
iCU/ICim6ZsuHNm5QbUKoy0NMVy1T01usIolcQLxxLzWAaWAF18GC9j45ZP7a/ghV7b0j6qwb+Sp
1MNpSM7444hk8xCJ9i0zkhaFuR+XV0VJpZdKHhLon/KUTaTX6cI80aCLNRyZ3vlMCjfpZ4+Je2Eu
lNa+isy35WZZLokomzVqWGzFjhDFAdthFHl/wi+GsGHU67xuNg5dvJmcNHAXT0PpGxQzjZE4KvwR
9mmIKLI12UcN1GknTMsNlOHiIrp52c16jpgrfnlGStrtmqLl53AQZMzNCkNuvdOIzdNt5krSEG/4
1sG8HGN/N68gLQE9YnDCQ5YrE9WeCQCsA31+3mQcX2qvypJZuwJ59dsh36XOtznjdDNG/OoAzS1z
FLtVQyFPr9nllWDLJbMCf2ZjSPAoMrjA+hD91xQ/dOocyt4Ccb8Mv4sD3SYDFxGljYlvcA9zU/CD
m+oitH3sg4PWjdj7AFk/ZxOeekLMYYbDBnHqHWjkhmn/vc+lpXAEiN/y9VXS2TQTzsl5KLz8g834
Jiu8a8NNAzx3XdAS84XxalnJxISx1ra7dIsUfYOw4b+5iGRoY/oO0ACwLK5/d1JHTlb86/xEBt4R
R9RHvKO3GAWmA4wC9HfklPRNhjARqK61Gq3vp4kig7C7S/BpSw/8JF4jYlbiQ+uAXp1TZV3HjAo5
x4Zm7TEmRdtEBLtrT+G61yn5e5IyeL5jbNl9UjoOeQmwkN08jhtaSQlEOCghD+LUuSiQsQwRwbaV
mfnTvcSBbKBucY/RY3viQ3lohxXLTXyTH5unT/Yzfa0snoBsXDAIPW4rfKmyshRxDhY/UblxonqU
B+1Zn+DN7dqSvz5XBVK7X841offZDTJeNKsEHewBOoD5K5WITSmb/74gknocFjFZr9Vn306cZfwl
YU1NJDKFRbfRo2hx8JhzPbKapci9yA5u47k6M5F3GtM2Kr6pMjYrkNGVXEAiMoYjS6bH8n3lCFAR
qjd/RGURBX9vSP3eJcftaUsY9UYZbDPpPDpg22xhn0OWimJajtMe10b3R+COisMLAgr+rRqimoMM
FT4Fhg4H6S3Za89HscIZypo0kwL0WQHSdq3ODsO32EmYk7b2ub3yLsjIQr6sIlXkVljfhQW9td+u
jF7rmvTjGElGJF4pKS5N+Piagw/lvSOpySk+Vgc7M1ULJd/MJQptGqrc7eyyHI4FD0JEpIHKjv/+
OwAthbrLUAmE9wXmSASn9ggF8RHZHzJJZN6MkN93Rpbrrk9By2tZ4bGubY2P5AJkZpNiV8yoxmw3
ojg4MgFZjp3u63kpBBBVtJ3VK41O5Fh2Cc89BqJdYTBVTp3bw8yPX3EiCzkOeUhpXiN37h985dZ3
m52pBFALg7njAe7jrMVIbH2DAawvYlTyqUpHh2pChlrASjoqdZ6ivDdffBDaLWKq8Wfg+/zcDnEP
iCM0C5HeM5lYhH7w1k1Zi/o+I4i01vm1G6WDsnDgMSYWE8SHd/xOS814JOeKlidYEXQH8Q2Sr6nh
41QmbenWn4RdG3m2Pqgad2KUCHhSAlmb30/LZagzHhO6MQReBI98XZUwV8+nRxzUhJx4Jj/bpQ6T
FQXWNBAoWqC4ZMUvSdJNzzRHDo2ikmDVc5onAn5W9RRd6+pNKGQrodLmvVWIXhst7/A5nqLq4VYK
pnG0PgLqoFuyzub6/pNoSgatHdWHw4MHg2mCRh2pGk58+TzEQa7pCtpBF5iWOX22a/TXN2S2NwwH
sY31aiap3lM0SkJ2fQDwXWtaYAiRtdpyT7VmMFjEndpCfC6pOUVWTZUqgg5QzgrBt1+DiBKyQs3U
v9Hj/iD+QnwWWnZ2Vv9f4Be+3qhe5ZRqrTxa2K8GPBqgHaBwCCf7gZV0/a3bWzKcgqNQqlRFW+9M
sRNe9ulmfXBDVKldel7mAYTxA9INHSzBb5hEpYAdeYsFcjCMXoxtj/eOtgvGa+xIZ796h6jOTIWK
C9lnT68pM9pY9EK1DSEGGhDi5Z9nZ4to3TFHCyEMgfUgUPB/qg85ebBoq/a0kGoaHeVmNTTGzlRJ
bL0sk7xyIrv6E/Zcss0Au002xBzDKRUuFH2UhRZ/XSELy78uMubPkzb26R2S2d5D+pmNuVy64dzv
vXETGNX41m8uc+2WeSvh1P+RnDDmzQdG23Rz+gGpb26ZHxZ3J80MInxqCCTQCfj28An8PWdoCTMj
DTIBsGedox8QcX1kneYgbVYDsH2B1hYm6w0zYDgRTgdgocZDf83yyPNMeTOStIXXsdMyt3hiMESb
3KQlDuHg8m9AlxXgLjdtDpA4vXGYACBjzX4jUtCExP6ynq7QJKhfd5/vY4I0bTqFGvRarkRwV4Bl
Fmv842gYDVXvny1LlUQHW3X5TXS6PkQbd5z/vPh3psAFn8OutVdZojLV8+qZ61Ezo8pLCHrRTF+C
nfEEEoH5RBNZ7/4mvgLWm/w1fRXJoWmuZxOL0mUF5U6cz7c7sXhoHoYyrYmzy366OdwdI9yn2o5T
J5sQGh/lxQX5xLVXboy2Wc0OY4ibYVlgyK3RacDmhuCc6XCnUlgTJKQUyOXH2rekDMvLr85egrLo
AJpkq9xZ34FuuQSZNE02lQzjdmYDizUEwX4ZTQLhoyEsKO726iXcITX6tVTcGvl9PBk1q7z7rjjg
795AyBNhJZcI8BxTAx1RaxSkuLwwFu8XnTHhS2BeOoxjz+jOCe+yv6/ab2lwyCSWSIUqLQrQXqsp
D0H9+IAgwrHCP248ZnObEA2JNi2k3/kDnlR78VydjR/T/fF6z1T9rVGDi/lxkXxUEgVE1qoFn9g9
Loz68B25/0IP5DgU9uSIp8m3l+WA+QSx0vS05m0WJbyzmQhZWME91gmDaYtfx0DRcRHgiULYCftu
o9rQfw0QJqZUbVwRNf3qZLZ8wiymcuw6MSpZV3La3gPtYJqFW3DbrfPHOMXGG6Ee/3cfcFoBAuNx
boUqV72RAMiHGjtIDw5Qe1lJ2bnK6m3UUxZSjLC0Ur7XbqCUb7zzP3QWpN97DiUzzz3f02rECGV1
p/kZrT7oekqha++K4fkbWTbME4im87+x5P3q9qUSBqh3I1btoocqJHyMSW7vy1LNRsT9tAqniCB4
PNqEUPYdXLISjYjeDR8xd+Tdt+6SW10Ho2J3SB6Ot8lXRQVgaFMBl9er0CT6mcrSgRjCi+Ybq5+b
99/4SJRC2B+VUy7OMSFGVbPHBgv4tfRcMC+Cz1ddw19l70+UcM0NpbA8mbgBz1vnc4J8vIcIk0Y7
Ci4LRIrxK/RaTy/PO0Ta1vOk8UQYERNUQzMvgC2JPE56ETTHkFM7RLUXZ7dXRmyaxlGXljStgQIL
yBKu+te48y2mQAlKTs5709W64DDV7ArgfamDNhvQi1miegfxIgL7bhJLlWQJmG6oSZBMMsLM6aHI
q/3fK08SGxTLTjGTuEX64nYjyMsY4bX5w4v2DIRe0eVOIGk7rApaVCf0130hkzxwpFl61MjwsN1u
PEYjGe+TfT9Lu2cKqmJu+KRoW6kQ1XteJLEJkHvpQCJxFgfhMB0xc3Hs3burVCVsyBKQyzl0x6fQ
FbjMJMsWGlbc1ZfiUUMCyL618rBEk79B69ACzKJvb8x7RffpNUnswuv+0bD7hiA/KqsLf0Yetuvd
ENrRnQjKjgoMsLi1zXmK2wqAUKBdHljZ8MiICqZvWd7Rsh8tBUOKJRKxHDIyvKrB3zJWZMvXMMoV
pMsFM4mgXP7dniwvRytL0adt2jJ/B0sx+tugfzzSZBs4ICi09qdHmlWmtdk0fgEOROqhiHOIWpq9
5NyZdbc1SXkKCIyGG6xyxBzVNDPi46+OotkDCuqqIpIf2Vh6z44XKWi3P9FExOKLTbv+Z0lg7MaL
ZUM3rZ2/ew8VhNkm6guUKkAul0rksloSN1PQyAw3eMff1BS/6VTkDPdvQuVN4fRgvJvGEBIa6lEk
DR3h+E9fu8zD7exGqtSysCZkBBYUbw1P+fxMUMsH76nWzf6NB9nXciF/ntqAqkvp7vyUAyy6v3Qj
3G74Y8zIwo1vtJr9RaNqe4Z1pnkWCIKuOv3bX4WlIhHLl08AnBfNL9cZk5BIa5/rIIyEVSOFRfcI
NncXfowZkL8yAVTdaPOwZU8sYBpe1oLtnvAKh5ub9idf9rjZ29rotCUcPot6W/EqFXM0Np6YfYvg
b7CLPkH+0xjnEnfrgRCM7Ff8sc5pxawzZpOzbCuel5qi73+cZD5bxMIFv1aJbKCYE9HR9VQLxe3+
Qbrx5QTeZlGOVu8C5LbR5uu88+G6V/71u3EIhxDWt2G4YRNrv3lTp9hqCOZxKcZsicBBqElyDg8M
jNq5v6ccX4cFcnato7oWAxN3+erD8enk1yn3OWNDXaBhFZQVoPgbioGk1zBmm2YLl02Lbg8DcIET
MUD1SD5motMjIAieWVqvgWBvl0Cw4zZ2sx90EzoWn4lL4wnn/ovJCYDFBghdJ60TirJuIbocYfwl
u2uMDmUhp27XV0TpGbEdZRBBCHH2zaxtP2zlowbw1LMrROAboZMyU3PXXE2zBF4NWKYAm/6tqMzq
eVTQzTfkTU2DBZpFk64dBQ5X2QGG77WTJLguDrpVShQV7EpVBadbOqctUUSSqX703tD0H09rmoe1
n57L9K1J7J7nQ7cyC8uHQMBvlwcAvDNujBH8bk31BsQb4UTHl7OpDtkX4/9p7Dt1d2njAoyxafXX
Rj99iZzJdkjQlm0YUKi8/o9659PsYRj5WYawW9yZUwcXo/r12dwmoFlx5W4GccW9f39JoMO6g5na
31WHZRP6Wj+au9FXZrghrMUawf56aERsTRMwNEbVZkQyDFIy2X+ikpQYkV+MJMNRovvmynZLiHeQ
bcGLTeARjheTRYzMf7neFAIbFkfH5vJzfxjcwzr2pb/r/p9q/HP34X4PFOBSNRsRky1MfCMgVnM5
r0Rk6gFs4M67XlB/jwR9lFTwmF1EfBAg64FAVNmZ42geDlJwKNsy04qbWFdHmSbM4wSFmRL/zVCY
1SDSd8pp74PQN4gi1fC/CXhAxZ+3SkIVIv4QgdToNpGrUYeCaIGAnJRCj7zeiyl+GGb9heha9sbu
h/vc+xF85rZApEi3WndKe6diZH0n2SqOZQRVONTVlEQ/KV3A06dx5gGxg4ObeAYgFvWR3q5yMcLy
gXaR9t/EG2Eq3dYjrSrZIExKxprNqYIudCstvCl2TN2OUvMyIoJ8vHCxdbuFWf3+0Sn8i8XEpVIU
MLRZ//I2dpztIgmC7XQrJFza1nleY/8fsGEobq1gNaLbKuQ88DP2t/TXZ4vJglN1DZ+lGl54ggVl
xG4HqXtiCS4IDs6GorN8rbGE7vHR4j1oLG7Rrnw/K5wpckM7Md3HiHKPs5iXJMTtqcg5eHdAa6nz
8Q+MwXVuO34TxzabGAQ6dCbUTugcch6aihOdufTKzo341pHZbaK9S1rE5w1+eDS6biv2JpTIL3pt
K5Zx+qotzXJOxJrkWg41cHOcNAaG7x/jjoy3iIsx+lOfYxAvw3vjlM6YwOPN0nuN6KSP8c66F87T
W5vc6pQjXCkXQTJ3bzZTJKlwAxkiAyG2TNaB3CQWQJylO992MR8GsiipMDAKQ6PICTHnzUJrrnW6
eytSp00ewV9f1ZOu0J01fTiSfT/mxtTNlD58beDnD++ewfYdhzaGobgum0xrAeGHyhLpCePwU+3j
NewRpjvPCzPWa1uiOGUNPd2v4Jf6YfQr1JEDMwOMODxCT9muHQ/z85g4RHLtspg6Hly4Q6wNC6Ou
IoOxJ3EnAK4PALvcGmsa8LhrUuXWvdLZRi6Ech7hduRQCd3T0nJIbPgY8n1XNl8xizjX3vtpjUV+
cvtamEpFNX8j148NRrVRM846iEDT7ABgT1Md9Lo+oeha+LKPBCIbeiqsG0e2P+JUu70H/s6OMm/z
AN71Qah0WWGpmC8FzkQ3PP3/HoYasgGoKIPILzkInK0Zdbn4ak6cWxig1YYqeq8oSmRsaV77SYZP
ff1j96q/CHKdKeR0UPCwheT4rGBOnMk2Ox2dHkvM2RIsBRSPQiOBjg+jSD+IqjZ6aKx8V+wvICtq
U5MC3SUYpSCu4RFCduC/OkQng/3LV6b3ivDZ5ev5U48utz0P3w8ni8Kl4Vgx13V3FbzLFwMzZsZs
b8nAKX58Dqp6cGjtd9qYhr8TSymD1fIH46x6y/wfuKUeKlIhckWDHiERblYafSI+3zQsEQOFmb8Y
Wy3KJXV/IaYL/A6g4fTeZMEcJUcuQwEWSqUKTeWv5tQCCIj/BAFfsiUvT954LlR1IQhHS+Njw8XK
s9dJyQrEllOetJ9WqgLKg0BpnCfikLXUPyfnOuk11Z2j0qIzN1uXe/aMJFUXAl+m0s2rq03xqFIl
yl5v6MRE/Mn+g5jhjLewyZSz7jMp3RtRabfMqBNb6g9Cvf4P+TN6NaNY+GNBwOvldB9T39IUsGQt
DXQvlXql47p8Z7z5tZF/G0Td0EfZoZ3c43cWfdg8VgKHXDfw22L0bIX2epklj7GqKk7NWugSC9VJ
ZM21WMw6DIYVzp4qOBkVPFHVn4uGYdOF2Qqr6RQC/5WcnS6RZmAIFLl3j/+nXPi97G4nE461Y7Wt
OeGTKYsTwzO+ijJ+DLtFEHHPaA8HC521XneYuKIL9h2BshHKMnUbzGeThwmhY+BTDNv3EE+sfw2v
iSFaEcDh1HY4/4TFdXLTwNQQCB2gTr0L55uktB1WaLE5hMNk/vyQVU/rNSRvxCmIVLml+69+sFsR
rbYQHToKSicrKFNDzsf1WwVcvBmw/rlu6LejIlqnUYDyzsbRpQINdtdEy1Le5Cq66ZN9VoSvrakz
PIFvamQkKeRF1R8cY3jwS2mswCRERO2DW6nonnE4b8pkEiH/kLEOwDP0+kitn6D6+Jc35ItDSyX/
VRyQMrRQw37uF1wdEAPQiRHEvPyBoRbJkQjWOKMvSVvrz6WFIizC5goEkpV9o8nHuOjb8JohTDLO
zEz0nHfL9wlravTNTsvLdmgLGOQ1Tc47jVuSGMqNKcJUn2VZK+al0tv/OMggKqs+xBARk8/VCk9y
26JHVrJMxFeGHxjHQnR0bmrP4iz8UBs10Osi3knakIQz2u6xqpue+NhkCbxnZSTQRMnmE+k987Gz
+6J1ToRHrtNlQV+M0Kir5cXvvBJ7QwUwSkqDCcJcy9V+F3fu4MltU5cl8RtiRjwbNLVbugb9S7Vv
5avz/snGLJO+yliu438fujnTsUnPCjZsEkDlyT46Lrw0YnfuRMiJfrl1UWuyq9YO6yoDYk+zKEMu
66eUWHKxU+Wg4trfzsfzoVpBH609J4+wGw28fsHhvAEAZoWlbzOvGH+DlohEYRW34QcBh34+shMJ
S2yZIll1nhWm2hqpmJo71I94FU7INxptb4leP1K03hL+GFBSqoFNzo9QPpA3gygrJs3veOLdkFXn
tNZLPYAqw5AH0dCjEMgI7DDAylAeucQeomuBu2Js9xZbl53JA/ILrJI1DNFcEHbSHwPwRMzWwXb1
KPqnFRP17usk0s3BBTzvCVsSAM8E2Lbk1YxT2nW8deLhAkk/rITZErn3GQ4qWHwyskk3Y8PMUUdm
Dvq9FyL6ld/RGq0uT1SfI+aDBkeESBRMt8CzBxBww4UVFxnVrNyRtGApIn51DL6WCtOCjuznR1S0
mPUjbJ/yYB1qiveu630SWTTLuRhU2kJH1dGg6oVIrLCd3boP68ucYr4/Im5vCjLCJAd7Yb9Ow9PU
FBsCd82VCYo8yzsum5vF60HZS9dwq//6WjghCzQSBvv4GKUDVcnWqSx6/bYNTlNCt8XJOMI85wMK
IYdO49eh4pVVp2ZBOFmOJvqX9YxQ/ppK6Wc+giWaxKuFomIECtoPtSPpsWocNqSQIV8X5dSjrZiJ
YF/QWqFbjwA1DYRmvZp4WlwGXCy/VNmg7aiiG75UtbhHa01IKrRdvvxCN+jVw9IlQR/1+5jxbRnu
2LE3e5pj+9O+jIiruyTYW3Q8PJM0SGYTeDbZFy4A5pgLFd8Ok8ln1GRJogN4kx/imCcc8XOI6xlu
tYrN/jwDcfFz2KfrjWzdRFwHZOcLTtAK49iTaRKjeSIpac+6y4Q8HU5pewT9SwCvDknjNroPRT2P
6FfZrlHtnV2+TDOBoNAzGdQcGgMBB9jpIGBXcA2IRHp2oDQN8XiM8sbEGvy1qz6bzVPFNERr3QKr
+ONq4iz1yUcCoEfSM9fnfVt4WzL/hxzkQxYVrUpbK36TxhiZ0Oa+f/I/bAi4z6GWuHHfcPxH8kRu
vzl8oZ3mLq6vjH05qpLNgg/+AnRBulr+z7MWkuJ4M9+Dd00BW9jFZKH50y8NyI+EEeqoB7Apiyc4
0e+Jw05yR6nd4J1aRVvJ4qQWBcQI7SZNxsRbGqHjg56DMSHBbRtBnMZ3PKrr70Dc/ghlagBjUs8f
5NNbBz5hc0mUc/sXRYmVTwvd/SfsV/74QzQlOtx+MomhcSRrryyhycK/YzeyXc8+isPDxUJfl0Bn
2d29J4OoPq4pGD5340D7xgzXzuEJCQHvvthdTR1HJ0J1nAjTOnET9O7En8+yBMyn9QhjkJbpKGsq
EraY7baI5dJTCEs4TqkNOO7cZE6edc0TQTZCufqodTYhifV3uTO9h8zp37qgBtDX7YDxo/Dqj/YS
otejj4kaGNfng1J/hQGaJNzqYL+sVoMxYx14wJJ3MV4+Y7ZcvO5CQDEk7alEXwZpIWKFJOF7lVsw
vvqpxaqRjAe+1Djl+hdkVaNE0ZBT8rrZaS8vdAug0DVj1n0Dz+Dg2fSIY6jaM5aX28kB/N0yw4fC
a6yVUYedVUakyHZ5YsQUFdZUk+LIPfhArIAgXO9/hjqf4RVwe3PTFceTPxUU/F1ZG+Y5CcxTcRoo
GuH/p73KlcJUDQmgZean4UBkAJwwWtt4WuwcMUBpIrUsBXbyTkUuBwHQkzy5bWP6HO1ICyJ3odsc
mpt8Jw0c7rBp6L+dvGr1Ck1PDl2+RVYb2RGQO6Atk953zuygQQcCVplDE0DP71rMAby5sjE3oApX
jRlH3yKkXGLXOg4WI4bss8c3beiBL8B+U0u9OYz1fGKKjGS/OnHJ38QAmlq9hJ+12RWC50/Jdo99
ocILEl1uY35YHwnej8QY3yiq1AotYO51viIRJHw4bPdQAN7AhKBmMq2ls8ov0R0rxgaBUTpwkeJb
VLV/yK8jp6pTARnh+J5Iy3rzbZhqkUP6Z2wdcAVzGlibt+cuDo8kK7iwcibRvX/WvQ4nIjh9xZ1k
J3wbjvt94+vh1+BfTeAbeDc6Hz/YBi+HECVdXRFvE8tsJ2AaJs1NriSgG/U2IIipDkojQ6BZcpHE
+W5zRVvL/YwI1eZfgRVZJd0u93vL2kRtmBBkyY1YcAvuvRhJgYynWaRz+DST0OrN6emhV6Vc75gq
vFj/V2/u7IeDY+eARtwEy6xELrBGDNPfelj0AXcy7E8BUcNy6pEcfeg28aY+DZO90Xzt5xMbIp/Q
G5oO2JS57mW+QxOlyWCJzhi5CcezFXD6+K6pZ1yxi5G2ZCCEXoXF/vG47gbxRC0CFQQzC+C4SVWd
/Xk3djo+//bYzo1AhFtwKHXAn40DM+DTLSAXfn+esFrOKb8ZdygRtI6v1AJdC8UzwWJmVFHOekmF
MfrBAiFUcwM+SmERVNCoywodBidc89vHUIqCL2pdpvJ82eJhBzRNj+fd2STASm5OVZPhVrMDYCO8
4Q0ofgas6UpDYugLDMYhkBeIexLmia2SHEeFrSx4pbpxzDDyVLD8ftLbjFCOOzecaKUACr+D7a3o
CsXHYdX5jKAI9bRz+Mr7MSjbQ8hVWj2twQkuDJiARQvERfKnbbgyvDXxXTLu1mSeDr7PXH2q/3q2
XFJlDmXxco1I6aH178xyP9ljS9T6W0fp89lZokkd9Yig54PlZ4OPmi4/WrTTC/Ms8aKv+RwKmx8R
cS8vIANdrT/qnURJyohmT47PxVtDEqMrvWq7VGOpCMmAbbn0kBKtUXOfp4xB/kfuw1NzaXSd9nO7
6yClFO2G6g9JAfI0Hpu+fzj9GDLVeouXeCQ2JG/+Ca1x0ciSw3YgGM1r1ML9MaLVvF9ghbggf6Hl
wzSKTIKuZemFX7Ke7sqpRMTSa7BU/S8CWS53GWW8SG/NfO/GdT6h/jaPDXfJzpKMXmol5Rp+hLS3
XbV+rIzX7EVo0msyMH2mxjoEWkPsHi9dub3Wo4vpczwKG0BfN2BrqCN8itmuxoTjPvwMDO/ftGPu
FSpyzE19cIUCPlMwvdi0Gb3pK0vw8tsvOdh3MjWXu+vs38ikd5nPaAluH58KmgXqCmmtJMlFP8Sc
1MO+NOKo98uqjuqgdpuzxtsLS42kn1WnG3fnG0Hv+FvK3U5O4lvLGM73NZFD3BCR89QYM08jYHUD
iJIsf3p5NsmOAtQdtals9CS0uIlkgdbjNBXMdsr/9px4rPiqcXV/1O9TrFLzNAQzDz6iE0+vLEF+
BJ0/MackK3kU5vuD2WpQt35qyQBowoTXfOT3kh5hLb7oehj2T0iSeIUGycFS6bTNV+0CpdrTMzct
bQSlmPTPpAzvL4fZRtN3uHfma4w9WCvZzYTkHbLPlMLnHWg5BYHIH51hmKGrOs5hkvjRzHY6EiqZ
TxaIDCECT4ILUbL7Pq7PTyoPNrXP8MfEt6M7PP2364JBnm24LPNmeRCGZCC4B69UuTH74NoT8tYz
moL17BDbjxLHjrh04/n/kYV74zf5E2SwauXkKDlrqwxVM5PQc/q5D8jDxb4J2qIK5x4s4kK3S0mf
N9E4P0FDZKkyyjN7UIccUzd6N+0auJXQm9luJsJ9Qu/Q3cSKB4TPmTd7bYJeMTyj7oV8e2VIxrwe
5MK/EFxhFgDsP1QVZxnoe9GPIX6p7Pg01ULXiZ8+2/JzkJ7pAjtWv3zBVQcnrS2WxI9IVK5AAXjK
lNbZx5xPsi+I3tyYLKQIMSvEkK19uVMnaCDxQf9VCfKf8fBXW8p2nt/+p9nOjuGhOFwY7EPviy1A
u93orSY+s93ZaPjlxxNEXOLYZ9hqJF+lODaDfwQPkBgQMfGg5LIJcN7wGNiR77Fk9qo9FliH0faX
q6C0PqeMPYagK8F6GCwlZY87ZpLSpTU9fu9IUmZ8gw+FEUJzDGDbpd74hoMSq0+lRY3E9X4//Qnw
8SP+PdNetxhQFN+weGbJHdhgMEcdw0KAHPDVciEji3wHvuo44B5Z+4O4bIYxswwYkmWvqoXdbeZb
3XKrixLa/wn3TS9bQsAyA4y4IllJYlq5UiZZ1BAls5oWqnaxnLJkOMc6+wmf/AGp4eAKvu7J7h9U
+ZmgJ9LpkI2gv2yDzFJB1rz9qFzIFBmVxMmVtJX71UQvIP2FpZ9ctjJesCbasU6xiTwDAp3o0gGR
kUxlbt0+RQnAC/Oe3aTOkvtrEnFUAbZPXsXF91vygwiRb4p+JSrTFXe7+KKyOFnAdM8MCSmDALIc
LJXOB9/CAwBmWm4cNk4LYgCnNkW30ZbNqnBknK8NUB5MiFIlsKGD5d08Rm5SE4JHAo10tJB6uCo1
X2wdmZwBtaOIZZ3FEvhzavhK47rEifohbAfYXn+tJtkqVxbTQL/EpzL61Jm+mOzoCLCKVnr3BQif
A3fKT3eoZjGAkd516teNPbH6Qql9Lo1EvCBJyr0nRpffTY9VjP2Jb1tQmwhSGmKrDXlfR9VzSh9x
08yxLtvqe1Gm72mPuwaB9j68KYpTjrOLR8XzBkTEzA/u+xhJZaXUkxvcXf2ukZkaskNqMU6oevmi
MDEBxTSaj432wikihNGs71bX95gczj6rRpLECuFDW/REkP5JtUKd/6a83DQ8o86Z+tMALzeMtbiS
oaYyFUetzDZ0uKYhUKBmbl6u5GEpsA+ZfXMFFkVs9w9rWXWVhoWwUI734lKnTuesoeZwSL3c3Fi6
Bca3r4XvYNQesK+RIIEKudF7Z9GGpjqzvrV5FcyZWUgMNqM2AY4Odn5KSvl/0lX4G0dMr5Z4wX1g
lKpEenisw0CuBQXCRkwU08d28btkByCUJoSRXRGGnqBc5R25Ur5THXzcZgg8MgHIbx1k8WpdTCWl
WoGVhKSPk+Oqi9lysN0vacxP8j/rqsW9Llg2VHNrl6SkuyxgB5mNkKKOlJ1IaqNLgIZkKnEaHmCt
1KJlhmnQnyiQ7xdgXipSE9VumNlWHJwzsa9qvunfrrID9HrWFbLidOCp8ubTnspjiVpDNhPzjPNC
sdXx3XUdqAxp3qqzXbsLhU69W76n5SugkPn6vb7n88HUfJFnPdu7Ic3zqMvtiXxgVYO1qwIYPqyT
ozWrIlvbtaWB1ZQmMsGwUFAsQl72SQbJVdr52nSFlFbetofQKL6CKK5eUz/iRiJ7aJziZaRH7VZb
z8nq08WuIF0F1M6znnDYOnYwlCTEnjT+qievDwfOotauenLkOIhdkDohWmnZ5chQJVQChWzShk1B
f1SPwdoFbA29ifkJlvS1srzxPPUxVbThKXpp42VrTlinTERMN5jM0VeFK1xETPH/O7pvooxxF+F6
/NFmJ/06y5L6MRZul+fO3e9cr/PFnLTnUleE10XCfLm4lQ2nX5lOSceKdQTfzFdOVy+pxiCrhcQn
DhCmgIrwzZ0cBe60Xfl8mJHH0svIw08DmzNDj8U1zbgWgcokRw3FlmqyQGedqSyG4wyORAEUCwLE
GOo0nwA4yTPGKLbK3q4wc1F94YVORFGWz2kRsXwfgKFbagXQs54obfcXuPmcHh6jfYjjuv36LxHJ
9dmc/gUkDIKBPUyJGK8b7eKYs6ca2oJvjtWiErwH/h6brqBIWD8nRk5YLEKggohVejN+QxbRKHku
18Mb8nKjyMUCNCyBKxo7mTIyEP8+HEpFWbijlmkEIn0SOwfHc4u558PuzpAh2PMsSAR8QbFFBgRQ
HN7jWJ9GdKmwcv8gLGpPadsdtGcwiR0POmIIO+EUq90tZgOQp+2UMMCuuD23N9Ch0x3p0l+v843e
nx7199kvYKcEZwdmcRr9lxQ5Z7+0gl4Pkeu2JKXekG8K0oxoeYSmtfHKHRj3gQtxC4prbqv9yVI0
+8EzD5DdwBFKjz9i4ibkkObpZdBSp8ckCACk/+fC4rIvI8621+KQe8OoOFPFpFdGhRGxC4AOP4Yl
xv2KrosK4Gzxmu3zNlbk+PZvQeoXD8nwyaicIqGdy2icN78dPSTaYKXoOHKvl6J2mL4LbSbJUlNT
QWguk6bFDQoZTubfEU9TaFUYzflAwcZS0rmu4KmjU5zJBURWdDelZ6Awrb+gRoeSEyqDRwWm8Zng
SZe6um+SnO2fy/dtEU4uivrJ+92N80pu14xJprHZ0WVRAQ0Km43Z4Dokkcytykz3qlHPmMs4m9ZC
0SgwfZQGyradzyel+tJOtD/ADHCT9gxbaLnbwqsADoYaz7a4ySlDgSciGP6nvKWflegCzFARo8zD
4rOgc/4Eht/0qjQG5ugqMa2rSYI9QxvQD2a5U1qS5Prl40q6sRNX6Cm7RYTyA3XMZ9BpsRioqcDv
e20SR5RHptDpmZ8DlHgn1B1LlwTkU27A22lN67hF/X2YmfvZRIzXBkx7MDOqIzFRU5qOiS4jfyak
SzfL8A2uRpijzcTWD3+UioHmll8VXNd82S5+Yu3YgqR/i36lM2+ulzebzTXVHoulTogPhIL0YVkl
UT3OX8/V/EbMOMVwpFM/03xnXIvliuExh2WVPf2ljyToKMe26m+6dVJ/rBAoXyeBqLGEpNbrFhBD
OrcsXI5T4Ll/dm1gSX4lVee6FQTEunwxvI3a8jG22qIWgeZ3axabFoBgn7jrQGgeu46OadFA8WfB
FmeH5lYVPlG3DIAL73OVAdHXGdVrgZqTOradjkIt+7H9Y4/i4ka/l3UPWL4M+CuPZbdLx7pQ7qS2
+5Pry4bWrLlynpoFFevE0gZbKTGT/wowsez+TjozsIGCwz3hrJ7odX0A5KLPKg/Qo3uuhaA9b643
k35+i+qQkLkUoWXKeMbCfzI/WNAUZFgLb1b0yJwxp1KiAPkgwnJ92aC4BIfUQIWuH7HFktiTqlSg
GuwuuE8R7lp6siFQmFx/55ahiPj3UKkvHkhJeJVzIqlXUGWWmG3Q1YshF5OMqu6NuR1yZAvkV7V8
fht2reu/npW1xboQ+/FlOnAfspwYrUWKL51LwuWnnUXgl/Oapg3ik/tOH5CjAzNUbmsUF6z248EH
Ipx0OamFw9fNVgazNxFMZ+vR2Cf+dUD99mX3fCkCKBlJF/HUzlgOGTVl8kvxo3DeSdLZBKI4pXHj
U6hIyBOWydzx+35xTeaqWgaAg3VQnUtD4UVA/pgS9Gq541Oi3uTb3efqASSwJ8tRcaeg6+ETMsFt
1+ArJHzhy6hUyFtYYDfgjAIzSOABOqWxGihBhZkmKlSzdHUF3h3Q1g27HbbPGmsbyIgLZdKEMp3y
BTJH3hYYboo6suFTANSfOriceqp0i94GIgijU4xEkoNrGd2qJ1BTHcc2RL/6WssIg0u32O65gF04
TTT4951xDZvn+SZms4yRF1vGRyIsNsIQH/YdT+UC+AZfjoemazBbY1QVQtgQZWmmVBN7EYi6jknv
0Vv//oFN4pz4qn+uDn5snumNAyZsWA2DFj2DO+hcUVAk5CynOrZgegNP/u55+vRBDJFw/nk6VnS2
2JODYBeTsXoNQ7ALoiJGStW9Gv0paaSlgqcbqf5AqI6Di2ejw6+rfihhD37F845XEObnm8ZtObDz
K6iklPqQy9q5iTJ9XY2COfcKl8ov9EmCKRwI3IByry+koXrw9vuHo8wExvKi3Qw0lFw60cvq+lEX
1q+RIG7Yjje8vf5hK3ZIA45IqDbBqOnwE3oZ7ronwDGrraoqHLxKZMy7Xa5pJOeUABvnCw+KBc7q
FmFbiSrQUV8GQ0dU8MFvS5IGmNZyrUvpRzL8pB88++A11MgHTR+WIelgST21vzhWkZmaJuJWHt6O
PvvMHu5uSXVXh0YcBAoAirHg/YB64dlby1FXy2/4jdvO5GQQSc5QqiR6QRz2n4dWvqmITdE/TNH/
s3hVI2qgDHfIXMOdLUW/hUtGd3XJr5Etr5hOynA5/ScX5vixev6KDS9YflOvRwx+YRSLxgNSV78F
HDmdfRnxthMQwbXrhPjc71FAZiUBiSNUBDL6sDv5D+KSiV0QKMDBKPbOoXaGjto6QyxIrkYkyzoi
S+IvYG4ae5a5r4XE9FUBL13J6fNUx40PXysfLCP9Q3P8ZM288ctyIZN/qp1R8hsTzAkwO/pinnha
6TZ1XFXzU8byt0mA9n8zZLGh1Qw+cfetDnjsj3BY0oOx2tyDE0nMMzBI8AhNYRiVQfuQ0OdLavpo
0gs91kjnVAzank13BaulN1QCQppcBbjZymrHhbsQT3o3fnjuczqI9wuf1UASAcTi6GLN3bP6g+Vg
FX/ejJycRzME9Wi6+M5yQavh99UTMQ+2OfgvQxRpZjqaMF817BRYZol5oLwuBHGUBP6EdsQeLjNj
zmXWOdOPkO0XmyczAo2JYgshFMeFkjj+YVN4ZUsx3spjze5DfxdEcHLbmjD9CCHJwuyqC6i8GFvc
Ldv0fiLYL7g46kN9bE9+ECmxHoUSiPTqMd8GO+HydxrPCox+9v3VxZFU/Afe14uk/U8OGzu4PYeX
ED6UP/3aTM9Af45ow/TKbog0oX9QWlFy344j3HsTi6JoxT56ZxVOwLpWDW8fd6EmVmNK1uOc+83Y
CH/e5Tx2uGGL7DCN/7VieLqid1FJrIVXEehoKTHyxOI80GbxUTqYiiqOt38yYwc8mz8PY57jTP8W
RuJqgYnTqShsrlpig1RzuZzhiKdftljOFSOcbyKEH5KYb7KGf4fppCV2hAc1sczuENGBehQFH9oq
0WQrh3e/l9Ps8uLQrT6kTHjWosFgxzfVt6wXJvor9ISEkjfD60zFxjYDBBsUUUaAfalsCxM/ruym
3buMLgIhbyPSe4qRdi7iPqWbZ0DHoggFaB+TS2wi7kV8Roa2cFrVL7OLZPddcz2h9T6Ll8DmTHOc
y99hjn7NqwjNh7LKhSOxOQ/C9wdMOCWuKy5S3GdZArKFvfZDreywUN491YA25jq8lFTvXZXmwyRy
AtHdPARNvUVAbTFJ6fZU/VPhNzTDsOeUIn8+eoVFWEqNsdbHjWVBbR/7QGPyylaBQpmYYycHpP7U
t/yCLIFnfNMlUiSJzEmKEfmLSuv0OZt1z2cBP6vNf/XnH9XeaAOsaHtOTe+CwcViphzepe3XilND
OjvfUddn491YPOkRGcXNZCmG6C+Fn70z9jlq/4vsU3walVL2TF2DdoYpbuLleTZtci22+1KJut8B
9X6oXoBf3Qu1PmVij/EYk6jwnw9WcgtiYwOgtoifyMhJOyb5nTdEYKFJaTxGhC5iMhnnlvoK8c4x
pShNmb5x1vPAYyZZddYJhkhOHM8rMykfLhhqb+zL+17qKZrI9f01at4ejQNgcAm+fflPqP9oOyE4
zrPWc78czDUCRKfkcLHwydKISJWxd91tED8ytzgc5CbDFbZ6LdzmPcPWFrIK/W0qR64/0RRYrSLA
4RHFkNK0z3RTfkWpOmVK2PxobW6UTBQHlE3coxU/yoQCU7Lmf5SAg5C3Aud+RMljdrxD8x6fYWB0
dF/srSkGSF401ATQFfu+iCGjhje9lOD+SSlDmWi+TksiCThxmOMot2Qr9vEK6CkuUhYe0hottJs7
8BsJ51yzX9ipu5Zl3JHg+Gn0Qv8fvgvbl2CyGFF092OgmLtJSqtJ8A9tjvmKipdhhXOTrn6XIldn
UUp9SBT+gvxILLV2vN1h0MWB+0Yzu73NYfnJky6tTX6XTh8ScD8/e5pl2usdNFJpXa1UOF1LzN9+
LRSxScTuLtC2fOgtcxY/T+rTn/1PJcL4AgViqgfRIAJ/RIBUUQmWjm86BVqwn+GfyfD3oGqQr/Lo
P6OBxMSyHsfbsThEC/gZQ1/mq94zhOWJciEPR+soypconMVNyBFKgHvlB0CiyBokQmcvPJuBuf1d
oLKVHizrQ6wRLO1j6xvExP/RQvsS/gCOz5UHza0T6bmsfkhd/7GsP6y8XA0wGTgWEwj57lSPwuTY
6ZIQvtC3GEBJkmYJV8mUT6SiOfI2pHOGd7mNqSt8PiLaU/1cswo3Up1GWA6VrJgbsrjAWWsf0K+o
JufJVRMJ9YHYDRjs41kwu7ALs0eBT0v7hIJUu6OLfB5+65A9r5TAC9vtQ2D8vD33dXO5ZXMcrirv
wKIVy+SACUDX1P0AcgSfh492Hdlg6GPQ42/rC4Hl2xWgdxNnpB+JW2MvN7Sw6NG+lHzdttdxDsed
onWYMn3DRhSr3aABSnsxoM0zdfZcpWYx6nDciqOLnrdMbNGxL2a0oORqKh0M91qs2eZityGyKTOI
pn4Z61h9nLAC/W68sg7uPB5k4oX3MDKhiSHt8ei+Wdg6P88AMp0WILpdfY7xEXCmC2Tuw42SzGhs
tZ/Mg9v4AxtbZ60MpdSmohYELmq6YhqQ0J9qrk3smAHZiSPZyVSFE2wDhubUI8x54L+qIQLt40xd
bgLhh7ZsQuqffqvcDNv+KqYEd3sgamEfR77o4VM5akP2WgTIuUUQJiNnH6+O5N071bO1nVMgvpx3
5V/he6US82NpYpyr50T7RJscWlwNMiXP7xHbjMdbsQT9Q2XqiOKIvLbhMru9YpRAM2GmNZmNNRpe
FiMOat0Aadc521jxZGkinGkyJVQhPFv+tpOaiBUXhhs0DzMB6pWlvOF+LDUGh/5IBMoGCF0w28Nw
pQoZpFBJB/ZALioe3R96K8PBMoDAP9h3TjFtwpM86LN/oF3sQt7cama/tGPJHkKKPqyho1Z8I57l
Ecib0Ej+p9RsE634CU93TLLSGZN6zou9tfvfEyNcmidYCeGpI91jGn17E2YoACI9VtNHAiRyd9vj
Bx5PBh0nG8fSpzIAXiHeFIGcYV+YjTuSME0sdh/qbAzmHVm10Tc0dW5nklPnOnOEV8ONaR9a4JXj
hVlrSiRzg7z/GNe+mrgjFLthvODn3ILKryL++x/4ZNVY5YeGMHZvsstKaHqR0gmyqf2f+95ehaTv
cIDP88NeWqspKCAoWWKydEpxg1D9U7Ur5jYlkas3n4KW7HZbUUEJjvGf6rKGAhJo43fBqNjx0f5s
AeJSl5eIYk1K6EepbkSdPr4HHf032TDGVBbepKSUsOColCnHx34Ehx1h4A8gw7X2urNT9h9LXQwX
323dqVLYiVO5wbRon1W2mf03+rNq0WP1olI+zL0DCoL0H2TcO7dXCM2mRHkRCKsMPtldPFOUxdXn
7hM828U6Rn76SnRcaVA6Y05qo+fD4hHkY36ldZhca0YZhoRHqzpdtTexgzEdAjAYCdVGLL48rnjM
UgcGuTr7WnW/T7gfk3XwZ2zS9nfXgQ8Ag//QJzKWpSyuGSqUTs7nVjle2X8t0bgCtuMfXhqAwepz
5rIGYyd1Y7u8ZsK4xC+eUadDQpV/y3NRZRt2JEhPFUvEK1LybiDRmUidSB9864Q3OXrYIoLz4KN5
WLSDLJjNTOey7ZHobAtcZ371MSL/cpztMszLgs2VydbmcYepC9/e4d51QWA0HGjv8KqgwwWu8mEq
DA/Gw+mDwlKpPl0agnptQdEwIFtQravOGmYchcQfREkDzUHP4wSRUBxG+S6qxi+aSfeMbtVW7SUO
n2NoKnHAsdNToNQ3r3+iwzCKwloT2xq//BtclIGpEJ4FX9p8fo3L3nllYt1a9KKje9t8hI2iBlni
TbkY+w2oFGhMCgJiomIT1rDJSenf3p/QdEWDNXSsXEe7fdKNLO5ipXUPcjlpkWqJjKD/g1BOaUJ/
OVuhlksaO8Ek9mtrObcLOlyJ3lRP2FR0RhB29L8joanMZaX2Knd+ML2A+lEu0ocheBsvwIq3n75H
xSGwnQ/Nq1L1Lu3iqyo8m/i1Nc70R220ACOYda/xag7Ye3yEc7mHezrGCuPZXKJzX7///HRJXjAo
9P1MrowwuIJqe1SYSOjuifnylcmEDIoursBTjWslYjPptuSsccUj4a7IE0NZdeWonI3vHtxaEzRz
RsO+d9Mk5rhTfRw6o7ehLmnn+QmngcF/ybvi5fC2bhh7HN0AUKUGl/i8ZRA1cZtpeSZiQuOssoBX
ViBVuJbE6VPbMF3mTGRjGwwheeg7Wq4ynpcgeBuuLz9MJbNd3IQ/DkEizzxNj1Ff++O6qYQBvt9v
UdGNGSsK9Ep3SywcvGHI5ntwFHmFxxqK3lnITZ64ItXkG10BNg7wWqdi/XxTSC4FJBt0wLdvI0ZX
zudmloYJUTXQ6pF6wjGBSUYuJZUr2vfP14GNLpVZcBhAuU62RQ3AoglZ6W3Wd72PiqcZChYlkODA
1yKSgphqMTbTFYbguUOHRNt0oPTGJhJhNh+fkCW+dlDCeYvPxhh1OFzEy/VcT8cAdJSe5TbPrbJs
SHbJdRcx0bo+GlHfgVH6DPgwiZ0X4328TKVDeQiQv7Sjh6EvEsRH4CV+ZzZtPNYPFCL9c4gMM4qc
b6jcRu6viPRhdv+oCWFk0EqzD453KBbqgbT113lACte+LuGccS4Q9HBT9PlZUvwpPSUHR5dOOkU4
nVMXgQ+5ACugm8oh1tWmiLKuUhQ0/hT/3qYZa0AaJc3fnB6KxKsBjCita443j+h3BEHmD67daW8S
cy2bVTFpbwDGcROoRIDW1UCCGniAJ5SyzS6gMrB4dz9dgyWaJwGqE7KUA07SOYhs8K9G+BCn1KGH
IKlPLwUco1UYy8XpLT7DzCV1jSA1dezEcROmOP9Jd/Dvknt4IS2uMJrYVQr8Ujq9UFEDsKZ0OVh9
m/QjCULlnR7PbxFMGz0QdUlP/x6VCY/8/ga7nSk/oCXhBosEVXWHg/ydLWcEXjbQBr5bDILe7zM4
mcaV+QVyleGIm1UyjQMX9rfVNXdiL15eN4X6eXMf075ncqHoeAvkRguluhU8zj/3pcWFGGT/jBe1
UqRwIudBJhkSES4b4v2VYGLuKsuOxsYdMdCsFQ06LKHpsLis85UmGRerWiwnAc8xWVFPvx6ntPt2
QqfZ5uRpqhvdSrAS7psSNR7h6C/N2fD8hMJWZ782f0R7NDEbJ+Ez4p7U+fgEsNruOVdtvJ0tjnH/
Oo9PmY7DLn67X19vkigr4nAQlNX+u1cP7pRUCja9TvUB8aoDikJ8zxTgikyH2raFb3zLbQZ0M2zX
+9uAlj0K+MlIGSVCOy3Otz4cVfyZ+puYAd8oPwiZ7XNHlUvCiHzWBgXukNmo7u4KKmmqwOtV9inG
YMdILWrAG5j+YLKuuaENVLFycAmNqrw7Vn1pyc1F5xy+qHxioL6gC2f7FP4L26UYy6IKmo7eJp/W
IoLpI1vn1yHP0reuSG7jON2c71lbiajVkMv17cBLVFGaWH+KvxQeJmvlffofpVzaLNqjbu9VvSkU
Arrn6lXTHbXCQXD+93g/oosnHpuVksaAe6tg5n3aFPATWyM0eUI0hjjSdJWCj8NrqhWAFuu6D8cm
FZ+RvphVUv2JB/ZMeX21dTAOHggTWsChbY/X7kIg3xhjRSLDOeWldLNvYWHT64aNsZwtkBJBJKfT
qZb34xfuzO1VAtuikHqNNXuzVkcjOzmFmYHs4/rnaY8yn3x22PaDM6NHDAjUoYKzu/qdvUh7bc2B
9YVR9dr1l1pFplRyFDaAjWDQfUKDSigy4ekQi5HHn8rHPfnwAU5E51EqIyBVNgZQs/7ZIrpVh/XN
/4eja9eawGiePFmteWJ5sSo0JDZg+Cm1d5Bl5xWLkeL2mCC8rYeGDCA30ZIZXbry2hkKpiJ/OyXc
IweQt7j1LhfSl7nACvK09poKNBoVcFbj5Wsud308lXMFir/iATKgiKmP7IUhTO2tnZqQxNbP5TYl
2YNtPT8krcr3d3GKGlA+IXbjsPdihIOZ9Hsf0IdsHJVVuNzkQkhsix3231Pmn9qQpMhOw0fJrrev
ApNbaay8hQ8T4i6hJ4mLhWzWfo9Ej3jlecWRnkETXMLfzV6NCxatkdQ96UU/XACD65Dhw2OUk4JK
OdOhaqswva9tWhgCZ4nLIO2zttwIF4Ja2g167vQAEEBk2Zz3zTSzk/PtuUQtfO1gDwGDs11iywOH
MOOIbHWzmc8oukGgeYXXsGnfe37Ka+YodEW00Cd4NAdqz8MzVGxhqcdMD+NNrLRtRv4PQKiLjXU9
fIuxwGzlzzyL/AZC5aTLWeP57lD2OTzoxl8D4UROojWQaKC63kHWDpvDMhu3GCYRKPniJnaMm20j
Z6WvoWnqv0yt9z0+memWL2x2QE+PgNyEF41ehxnv6fGp2yYA9lF4eS/GNP8ck2zU8pkYgGfvopty
AfApP7XutOPUiq/9w0eccFOw373Woo6tNJbA+GDnM3pvkQ7k689KttOZqQf/0TNImITG+U7elYP/
VzOW3X29EaBx/I1qpXn3usJTSm/gQXKzrGBGHKJTzHlR0FUM/1e/adWJq1hMokwEgmAvA+YzOUPf
wsP2ldGeMxrVlhXMRyvO8XIys2RJQm2lolOkMTSOqaFxpCFwIY8TAy0wOJn9/50YNC5iIElTni6N
PyOvKI0CHiilOXNf/wiTMG0Gv9/2vZWgpNFHCOh3iSKgjiW7slgLZkobFUSIDlJLP5ejZ6iHz//W
pAfDbYfr0EF8tal2KMaz9KtrmHjOZ6vsCNpYaeCeQaLSpAOxA2rZJjK0rngSJPKAencUhxc56ogX
ZBwnE1AnEJCe6i4nDIk2OQfjRVNZrhADFF0q7bqW4fHwJV/Lt3G9YUQoLdqPGnJy6r1VWST0twdc
9mtwTrokpsSdGDabTITmm8mE0wKBRh++tOe96iHIubEyPRRIWcSJuvUswXLfh9dqvANsC98W34+q
8JaaklArAjCdO1T2rlXfS+sXrbkeEUALAG+3pD6Qursv8T8CMeEZ0YNW733ylbauGSKIsqHWdByq
4yZdxU5WN8w3CFkanG/drEouLL4K8latP5qA9vLHTl4TfIbl64ixPLO6/SFhuvVd8BbbLsOcKzg0
36jFt4vDInF7wwTXXCAewm5OsB+jPpJd4OF/5R9gbYAZhHRF1480sooRMlaQnejIDrr2Bi6BcP4I
V24uQ6No1eZv2sZjBeQGfS/aEaz2Atz1A+pxAFCTWFTqcfgViCMPytU2HGFx5hYS2DuE2kSdlVE9
kFBidT4ISfziSuiD866xnSCAfO6xygFKg8x5Rj4Mm7V7eqmz54r4K5tH8Iqrqonu/qRITZsz2dUC
tJ43eXAbcFkc1QaoHwpOeJJ0TvuJhenWxuh1/RtiCns+KpfPX8jwoPEFpF2xkJ/IzWLemqHJB/DS
mbEbPqsYAEVb1mASUgxALZ0xQ/BxvgOwoWJxbGw0zoD8H1AdGpwo+VCV7STQKmwsPoUptvbSppdk
5+p+HwqPsdmrv92tUtSwb6ipvluHzFmeuhvQY7Ycue8UUNQs7/UZeXy+Wa+0QXNw/lrk/Bs/vZQ6
KsI3EqSJevuznRbSzO7J5W9UwySsR+5Hy6JYE7l6EVIkvTvQy1rkL5tVyl8018UlhzevrHWn6Afo
HQRq0QQa6f8IVCgReK1nanOSxiVid3nw7tZzag1LkbYP2SoZR8p1nh42iw1e+qCF8zglPf7rBde7
0/IpHRI3L+XeTR4bduz7jyM/XKPraJAevqx8LTrsoqh3uN75mogMA848SwWFms+WPXQJ8JE2IDtr
wGfw6SB9YznZUZNpMmfx+kTVgENYpgC5B3hr4H+ZeTm5trvMz5O+llzR3eeMHNc4t1mTB05LpKEb
rBgIGblJclKAgeAMVVQO8Nt2RqT6YA+zPEoD3a7b2hoIbszW7A4CZgj79T4smFXZEDw1GU8FTBPl
vzfVAb26wKhiGzF1rg7I0YZrZrVuBoEyqBudLgqlRRPPF+gk+jI2LahgqMJxxgHHtSqmjec9kVJR
EU9Xk16FSY9tkAfuVJSeYRAAkwgYp5vikeJsinEtfXjsdXsRohPSB8WSd3qV9TkeWrdEcZHuKaOG
IdEe3Eb41jBZXLS1+ik3QjDmEhEzwoopo5Bg+xX6HExqc8Qb4gfHBHXhfTUwdJDpeJ6VEWOYdTII
epmmlt3do1DAhz/dkwfzq3qkT9Tybp34jq/ku+o52VB6Zv0FntrOuNPh5h/cg/dQuNG/SJnSnLAN
GcoTAZfzVYdhnu+n5QnKIVh2MEOOtGm2Zc/HGKsVXfvqgexphaOAAd9szW6biwJgPTMNc7VjzoFl
i2t9SIJB7pGhxnWQUuG7yuTo75GgPyCD076cGH+S7wecqNhNxv8iwpxwHzyN16khjPg6figdF0fZ
bbUEHvKRHNRBgjMyWj8LaIjY0l+VEc1ed/3Bh7hCC1TFDG4681ElJ7h1u0m9Gj1rNWf7fMuBZGuq
DXIkCd5nkvN5qrQEkmFh
`protect end_protected

