

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kv0N+ODrJQAnD45jVEsSEPytnysm3pvAbJ05V2JaqTdEQNJrijqrY29nJXOyqQOIioMFCyAehxdh
SS8dEy2RvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wl26nrMFXa6fm7UAkMFkRbwMiWczBO907OqYX8JeRapSfb54ShwQXeaNsbVvqp4GNYQWgD8fiWsc
Rg1ZH/ALNgmzzsXH1hqu9qf40O6LpbgjO9M5gvRZkEo/Tsa2oqZnRuXHxvGdfSUWwgm16QfnXWFD
HONMKYo+TnX1BbyoHuA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cF9G3LQheZJrMO7arGfYkxyoON6brspPywtxFKpTvNhoNGqsA1QaxZgfesvqKSR6jIrBuWrdpeSm
PoQl517JxEpEF310dys+9f254GuonHdyipWsWNgWjbTCuw6rYLvLG1y7lYwgHlSqKUNrBaGYERTL
bx0Arf8JZijWzxoSQ9FVJxjXj/PfvGzrh6e0n/oHLpafMxMPZcDI+yx5HuAhNXSr705mAXB8bgRf
GS+N50n6SUyWqcyUqw3kHjqQ2U4vJW+j5ZC3mQaQb3xJkZgzHfCaBKMstoXIjqY6XkB5Su6aeqKF
tsdYwq2h1uyBfljsOFo3IsRsUpNIiryBaM1j5w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fN4hvSzwAQXVTyvBcSPI9qSFGq1b0QWYvne9odu5QkpUwhn44DFKeJSRI90o/blLQLnT5fdJ1IVC
mwqzRlL7DmT25nQgDxB1mM1knf9aPQaDbovHFOWTzAPBPJqGcsU8B7iu5g++kkRlIJA/0D9NUZP/
zdeXDuR/f3RpGDQ9X3WIBcSwde7JdAaZPxu8gycDj+eAg//eJ+Ch+IApwl6KjZF7Lov59CHOoVNR
udrlY4+R4MFUEO48SwDCDlqVGTYZykUVxSqzXifsrNKc0qKvKF4GbqbVHDidoVCoh7f7Jnj0snvM
x3DFGPDnokqNpDBX7xF9L6+GYPELuxQwMV3Yog==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MECPOWJAU4w/UvBGQeSeElgdlWQuUK1on5QTAzUF7zMKC1Dzhpw/yWAmwgERdTOHF4jFwSXDGCYX
dcq7yoSgrYHNe1Z9FD7/4uOTgF7lUDYslV5k/HR/cVW9QWbwl5jLUaoa4U/BsWl+xPk3gCXBhT1o
1qrFxMGkr18FyvER+gYFNuGtJOdwhkp3EWSeT0uUZpww9gD8GQxRUyHQJxyLO7OrJ+p6c8iZL8us
t83ykRj64BZ4A7H8a4gi13wX2JOPHaLBMG6QaY9NxFK4P+cAlJ5tz1UR5CiOSua4Nbo8RZAnEv5U
qSe9Ctk2cb+fZHyT1Jbe89K38c/68dSDrW+q0Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JGQumRp5idVwKA3zzoqht/27epSOGyhvfg4tXP+tPHgo6OfP/FU3H6/X1Nd4Y66ilN9i+iugj0ng
ehLY04ISDe8fLdY/NaZ+qOkmAGDYirT/RxSo79rIeXhylLKnHv9FphaO49Z/wGAPNVJcMj7acDAt
BmSxt3Wb7gOV2zsovZM=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FGXHNsFzSGXjbxp7bvoF47vhF8reHgBm6BrifhO2QcSTwMmIfvC72GA44UQ8v8jHIWHgPlay/nGH
qq6loQoHzagZ/voRdMzWla+HchA2la644cxBm8f8Fq9WGjAfrRKdp+ka7tSEmDbdQiKs1i43XT8z
Q9z55GPf5g5GdS4wXPj3ZM9TkEPcyM6MWas1txHsPj+r/l+N/OJNLRx9g9A23yQcrqoY/ibZoyFW
/7no0S9W9Nh+BPh8OXy4CwqtsvPd0/Zl0/JDLnm5d0hcEAn+3TkTvrZq0NgpjAEEOfrxtp+HqvpD
SE2gPjJVpUBZWou1zkZKYyakXZCQodq+NDtzNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
C4mKPLq8pHcljMM5huzuumEh8R7Hl0dc0eQegMmOn88bgFywGeEM5qtH1sYvheV09lJm17HaI4Fp
WosNHgryKEWekPQz8+67ZRkXdyA6BkQlP8vU6XQ/NJaGXL0+MBINW5oCmqMPvZ2jI6dexpFKD28o
dXnsqs7XAQji03wQu10Ise0FOBPiOpE7n+vIWIQhhbZ7nMYYQxGbMuQhbM65j/74WWsX3XH/fYUS
yxlKpKP1JmIywrnpewHUCU8WALBzvtK0f02TdyPC2egNr+jvhbS85iAVrR0DZju7fAnYGSdKLn7G
EHxyh+ZFn6C14QozG1LJ/wjw7RneRWc0s5JJktgiOWv04zlf0eEELHGdOcP/c3C6RLxfKIYioDY+
zh4lJzVWb7iT79D55p4DHjCxWdgoIwmpNWHjNUkpxRcqGsPAS3jjMK4kTes/anqI+RyMrgSh5JKF
bI/3Wnc7L6aAsR3nDekNU186WrAXbYFIKzHDVLfLpcTE9Imv3APVdGLBTggijSqGu7I8kfTeyFaK
WK+P1xgh7tiJSr9zc4EYFDi5WuSGFb0lD7G5rVOpOBVhr8vkU3ezg7u5ymrjZnBs7XOS2QGKrUad
f1OKp8rVbQg5vtKwCX/Vyo0D+F61krIGAhjti6DrHgBjLXShadsuTMl/eQSrehoQ/wDOuZFgqsXz
V63E561xelaG7P2dpKLMKpTzpqleTYnLYT9xm4b5cvvVI6AKmNvEpQWkItcNua6WNGhrDhNbkDNl
r6rNvISi/yqSC+pt8L7ralfBpOhm3VAZT/dvoziIavVmlEqkW1dheXTeQZNOze+ZrJnId/EqHrZF
6qmmOb3TRJbK2mv0Aqr0Y5DuRe350ORfQOhHGbem22WW8tAqUMMAvvlKiJXpMY2NpjtcxehzvLfc
FZfhussThsT04FJBTiOko+kK06rrj4ROk/RyRj5dsdEHxzY1ZrzJCNu6ixD8fMKjKWxLHQH+skEj
/HWkQPwK0pnoXdRH4W9mOqI2I1lmnLvlKNn8PgNXZNDlOSGt5QCULeO+AGL3bjT8UqY2JiXUfncf
0hK4ZM+ErVJOtXqF6cfBTV80K7vGVLkYvLat0f/M0HhC/J0Ap5On/TZLIAGX2ToSzOsOR5tp6f9X
Sisb9VC9hW5Oh0EEqsmzwhGXrm7LVWvlY+IiQmLTrNCKLMomBbZ2+5J94PDRV7hCP03JB6HZOUsz
e6WVO6DipypU4ykdlLN8F/miGKF95CgV+PeY3blOlXgpAlXrtF9FMKfZ0E2stdVLM6TV5D02B7bB
ns4WTXDZeHj0jIl+UrPhi/HsWUxeT06dqU2KrUW3D75RreGvw7T4uppwfKgeujwk8JmbfkLQMfYT
Id71Hvue6yatfYnDi7HF/N3lpTxDT8fy9kJmCSYguMG6evpeK/8hfLqoQTexGyVhGrKs+QHEUt2i
PjOGO/nU0idmoTnR2oJhQBRS71WTlUSzMkkZJ/ElT2HtFIfhHY0SXcbW3AoxZtd8H7YVzI6KMST1
F55h+W6YosyO/grg56q+ovyy9itUrMhlRih0ZtSr15T3CMGhlJlr+2+9C8WUC6kD/2lgvkIX76O4
7x+f5RMoaIDpkG1bxQLLliw3gIkJOxL3aQelOuG3A3j+/CIbhpjO5lfqQuq/zas9FwZPFWOe7NKC
RnGRVZvwp+ZZPRLLFpu1vTAK9/knqnCUtqWF9A7+4tJQ6kXIBGSx360kQs5AsT2a1iIQDbekJM4d
USy2rST6hGt2RjTKEgmlC1DMzf+f9uyVYsPV6VlAZND6yGf596WLYE9EqvGSWhVNbWpPjy7sIOax
PabdQxJcX30GA+OjpTa2bSDKDSqO9rM5/hk0OvGo4Y59mQ5yyiPrbAjHFZ6ecMbn1KJayHwkWdmZ
Qk/tu2z8f5hLU/NA6Lj9fLwBOo/LmhIZTMqxkpR/X26EJMCglZ8tS2aHex8H1O6eUZ7F8mofSlhD
3O9mqoqeK5tuXBuKzmoeajcrwDPLUuwLQZtMSWUdzfYTMyrKygdPizdOIWNsZl4fsIZWpg4Ezj4d
mcncRTav5K1qzaPR7OdGRkoz8P7HXiomODWqrai9Bh48dgOqQvCCL+VKWAg0lcBfIRC1BH3EOrUT
QHIRe/hRe7mvgu6hXKcXGgwfS2dGeNniW3JGcRpT00t6M44mXlYrHt5SMCs8PGrRc5MNc//NGgfB
LhHPaehMgvcrLXaqVeu9JHbIS73gqqjwgmWOnGFigq7jd+VHPtu31G28pf++imaTA837ImpfmkH3
iYYb4VMDBFRjiom1ZoKfAH8qOwcV8OvSyuLMY/s/RqaiwhlfF4NZFGRK1kY4VEIAwpQjlARU3T9m
Sm/WfBdRiq2yKWHOs/YMipnsSwnoCEcrO1xItjH8ZRbrA68wDDP+yoOPURzMFjTVzpSvXH+ifPFH
Kmzrb4AVNm1c3DVE90jJTTesX9wYS7y8UT+4ydEsv3I1iccXcrL7UQmwk2OBpF2Wz/Ojl5N+XVgn
YfESCzl1a6gBhYv1rDZiLHtSM5aIEeT21T18og+rvkMtTObD4Z+eLlQ2KazS41WYQ8H5CwRRenvl
WPYNSST8rzoHgjm5ETWcllPI08YxvLsnF2QIXu70qkLtV4lLCvO6F03eCosm8T7A2rrGRfpIQ5/d
OH8MOUwkfLjv0QH853ng5JdDgtcf+arJgCN8o1VcAO99OTzAmIrttFRiGvdlA39VHz2MzLvS8IpK
at/J8ykVdGjaQ4lycr2IZw8Oiya/0+FKr+ack/fq7hxO/UZaxIB2PuPJUman3lpxFSaQ97lzBeVW
16ROY6B/+U4gIEZXduRdWHOk2HfL8EJlL59SNCG8F1gygBpi8i8gVuPftdk9hScZ4OsCN9ysQQdy
Bs8LSc6BynwnBzX2wJzpLNWLYtU6ioQ96QLWaU3s8DbUTTZ6ZTfJtxYfDNXjMXmBQDZS+kUZ6E9W
SAFgkdUSTGxTyjMNCSyXCjgYtKybf1N9klyAOgjtSz59vxHg91OFTmvoo9RPfJYzs3ASvTB+khDq
hX18yWiYcHgRrojUiwK7DmKnLJizZSk9O6Spwcm+IokRn7YfivUpqVi3xKLmglOwmoJg99K+kcGf
ccAhv9Y3d9nTL86jmIa3aSmFKBhiGiAnA1GpfaaK6BkYqNZBrsomspJrN1GVA+mJ7ZUzhRvbNIUN
Xk0hePnSwX+AwF8DKTD2qnNI2QWS9Pe5em1N1KeKNCa0oUGsUHnktaTUcAkzmB2zgFNDRwYNv4tu
rIxVEV6f701/8QIbFEeHaabB55tKqe0Sl6+JHOpmq9r0lHEX6mH+1vss0u8KP5SKNR8U2lJqPllk
ieAXrcj40YdxQgwoVdUNuxJ8LeCa2h8xHjuC6cpoZKTkY1uAJVk0y7hqRuZTilr7n36ItqYUkS4J
fwh0kTX8yWVdU8Q+Pf7YtjJw7JiXlp4rP4HqL89aWC+/kE3jvCxk1XISeoU/5NLcq2p3zkucF/PG
i5EAA/XZz68iMj74sDcOvnpHLdOSp9YwQkPevXR7gI6p1k6nFNKr+ezWO8U6LDPfvAZrYSCnjMW+
SJ7+QXBDNujFTp/RwWACrI+1YU35UkfHZ7sh/mFYBEB3PIby3PTSNNaF4CaouQr6+AVJ+sxQmoLT
cZcTG82CX0jusgc5SbdPjWcUf3LWYrtoQlbS2oiNZrGjTVofc3Eb4uHZ5YwnRNjeYSip3wDkVqhB
s/cywryeY+dPEt1AFckHREslLT21T0t6e12lHmUEjJomMDCTg3veCrIKiT6uk1nz+n6Q3IAc1BTd
lyvrZZSeRSCJMAIZ1TSVkdCyTnEmbPndli/k2zabgJcLcZkogo4fMTRlJhnx5Qwi6SBaYFHmpymd
NbQ7PspBN4DjVuOpRAndrb2F72ID1nm9cKYJHL2mLd8jSdrYaqlwVgEXmeecFQrfPaWWdoJRgPWz
DkrXiawjSV6KNZSa8VFEvwLms5mLMlutS4TkB+a1bgm0kw8LYELZjV9wi0oVCvk6Fo8jmlyFuyal
r012teCQZKWCY89drKAdvLmwMgUcPJf27A2MvTyT/U6BamWFtDnUH7U3C1aU0rMlJHQN93Y9Knnk
sCS97wjSfpwW4M7lEjJnQ/9lVAZiAktGCiYOsdAmtDXHCR86s6utb1Ll/WtaAFQmZ3hokdsQ0rXS
ib7lv1Pwqyn9wDH/hBok2EN4HaJc7qlceEkGmX+3EbxmFDAaxmOMiWT5YZsQCBCExNmTFvJKpuy/
aSejfjS2UGk/xXpRAMpJx1EWHQUztkdJXuyWCyXfAkAaVJBYlfwVc75AW5NxctMxr+m7+PNk44Cf
FOoBYaVp9eehvyn6LQEPSCE6GFUSa7e7MSBv6TND1D3KPEn5LC0B1l0MMC6F71P/I0H1PS4TzYs7
E6QBdwpYariGLGHgbN1CXPQh4SLe0WM2l3b7EBFWQ8miohJlwz5jr0YueU5ORtyz25TImyRb4TaS
8OIc9aOkstElnnNH3PyRVk6QyCTj4TrDuJMp2Wrqa7IC1ev2Gku19wnN+BtWRu1w5cT7k9VkgJfP
04hvJyHzEGf41YOc3j542v2iP8pE5iXK16uVtM6e7MeNOwwEMuLWFKyTgZJBd8LFudMFFqdEl2sv
mFXfuYWTdXUWkQpydkEU1bk8ailWVcqLYxshxswWZaA311w+CCfWqfY2JO7Q3NeUkDP51hqr8y79
50Gd2+SBZ+PBXfPc+ZyxZLIjY7o2/hcWiBRBy5cV1MRN73xsFEWg4Cw4L58aPu5ZdsuSmdEr+utQ
l64v4LoqL83KuNMfOrUdMGYNWbeYIHwPj+XCKKcZitBYChE7a46E4VizVza/82PMlbFcbPoraDKC
rcQhpu4nLIJ+wGtICQ/XC+1WPxYeRZqdHV+GYHu6gGsjFfV5284oW7RRkrvvncl800HZ51wPYKkz
DU/T0fNcoUeLBFSqFAhTwF4PyFUjfIIUT2NPalm+BuJV63zC0/sAvUHfGYl/yU3DsFNbcIZpSfaM
2llyTH8pAFbZ0r+ir6b7NniB2lx4GBvpsDajw5gVRdAhGSo7kvXZ+kcaJlWsW4OfWB42p0J6qIF2
2KP6eLycMLeKxOJvpPn0kQ7W50BByWKwn4annAzmCoV2y/DZh+vPc5/x3F6sf0OsSIZRYU6BxQlL
quRlRCnSxn42qIxIuURLUOw6Xn6NvMJ+sHoZTJT+S2PBXMOwoYc6D37tf3rPvnvOb8QbHBZqzK1r
yP6ve92gZr4dMMcsHtIaG569NxkZ9GO1UP2kitvegSxtQKvm6oBmIxCR45bsQpoGiqlmYJ6D0hTK
bux1/ffrG9FzwI5f21Ns3w4HlDNP6R/RFVF1uN2izRKOP4Aww+mpDQWmy2a0NjiG6NWNccsvGua9
fR+DxyASNODEWoWH1/Nkz8LLYqJQky+BTUqhuDtZIKzn7h7iwm3DJ0rtWEXWRzQU1e43UpEWhMU8
70elvP8vi/GvexnAxRNmlXqMt93sp4no1RzgOqz52uNAnS3u60Y1SXbeskbmRLEVsfPULWhq8Z2h
Z+l4l0hbUFR1u2zGNWifpF2ziXUcoXsS8STr+umr+bT91ZoF0p3ZeT6gG0IpCPOs31cepYO8q1qJ
o3Iqb0HAmuvioKvUEa9LCQ3tjgLfZQyrEI5OmFHOlgRL/P9nRCiM5nOcKX6Mw9An5LIi1BFN3GQU
GKq0QVgxQJUwwkVPYNfyoQsIiMABRJAQ0LpxoHMlhCHY3r2J8rT6xvOu9JcQ1MFvuMOYOIQ2gmxH
VO/WXVQcFJ8dLPnUXJqrVQqYgJK4gu3BcS6YGMu28WwnXZbN4eOy3pJl/A7un5z62yq605fnMNYv
DnCEjqjZMEIbW80XD1JZVKFNOjTEHNdO4rwa8uzjU/YE0D4S/ebiMaK95KjEJ+TKrI0xQCBxZNnc
WWYFqqNr6q4eP1s1jRDeztHaC2EcCItQI66oZWAvmPJBSTW/YRbJE6x+GVdv71j6nkfm3cXwMF8p
GhvJvEUSlcoJQgAi+lvV8hRMNQ87WBpUuZHJplAjDGNe3vNQbC+ceAI760lXb/ef7OCggSLtlS7T
nQfMNIbkMVukckd9968KQ51BQ1ncraZuwf7InmCiIwZfgTzx4XB4V4e6uAoB6eztRmTXmvUVAXay
AjlUeHVW9rTTd5Wwyjr9p9xNnvPyEPeyQJWREbaImhlFMdpV4Uol1iaVzU1PJ1FuPOKZkacRqeb7
gjXFry5U3Ud8CFjqPuSyWY4Nx8W9QfGf+MfJKnrnEbMwEV7pXFcSkG4Gd2ht+Rrdu3ZdrORrf4Wl
Z2EOI0070OG7PiWMRwnkBQe0FxQZXr1IMD+awjfB3qI5d9rbsoOFdCKyqEMDw/MzLN74tHTq5cm8
jXoAZ8d+x4MO7b376LByMNMw1fxR4umL9b16ECe5054Xs/oneVxmyL7sGIjcJyIlQzKwjycowdo1
sTEQaMIzXjB7imwcysitUXylXBxFec+6hXMB0+OE7eeoXDMoW2/RiUy22THBGfBMtuN3IsMslT4h
+DabkPvYcoAvlT8rJ604qe+PsuPVBMhwTJdJcc0iVfVFeBm3XAhc81xo/Zu9KapvzLqYqwxuBLGA
815voTpUSCAR5IXvXEIgHSYOjQkJgMPC1MidxatGfR1Spv+i5R4ZrebIlZdWkyXVy5I1eCKXOdEm
AX8Kb5osgYT/jAP/t9LnqrX9eUzeYrVvTTl5c7O8nE8tQ0bsaclUtO1Jg1BMqtD8QmNKgxELtfX/
jAka6efcpK6+5JnjEfOZSi7DGrH6popIjaiFpg4/tJ/Q+D3JvBuf3nnm/i81RvK+aJcRTu6Y/fkv
AJtzYwdOOI8RCiGm4Zn+RxR9+rZNj2SsZOjLZXTHA0BUMJZL2tUz5Z+7Ck9Rc3qKDGqtvJzB5rM3
Vmcnjk7Vt60eHpNCFfPduDabpCZ4zVHIhUI3u77FMcLYlQp6EWUju5AbPtpzKExrmxwoobZY7XiM
1A/HHYBGUR9sfRqzVbu8U72pBObpFLOsgmsIQOKLQLvtLs8YuR90MIM0xlxe35lwtS8rgVdU6tub
J07o/0mMSPi8T6SWSme1nxu0CByOXbFseduPgDcn3gDqylgtfCURPBrSWjaIP6K3P+31inZtubUK
//Qs4IBseykOiS3LLgibHPSOmzX5mUEvkVOSGk1yjz6Faw4LbNT0Zplcpjg7F3G7hU68JPBgZytx
s0o5HsB1JoCUWDCDzc+YscI0YHRNC7NiPSgTHE1nBdhiW42KQ5xHKgi3AI+zgKQ1CE4lUYaUn9PS
U3RWvsiHRTa7fTO1pi6Cf5VeE8ItBhOn9eel/wn0o08uk7ofYgfteNtef29yUB+I4N0HCkAfAsYW
CcEUd6gHlxXTn9SkamFsPaoWtnG+U8nMN4WZyiLwWayTZgVxP7b3LgMiHt+Gr9Qx8PyR5rB9ko/M
BdKeOa3x4x1Ogeu7TlGgR/DynZJ4fOcFloDw3U1ZRJmro7Mrdme9/KBiFdo6X3+Vb9EVdY4rnRB/
sGRk975QeQjYpYmMmCjZ0tjSwTkXmEuw9TRYyNdKnZX0NwDU8/5IIMOYyaghcvz8ilBS8HupKLfe
1jTDQR4i0/9ZRHZ3/o9QY/831nIzhyKFyMb7PPKwvPb+EvK4IqjxIwdugIdfd/qXCsVwSQnF6xXB
BQ8qew+6XPAmMefJMnHhabq2hpapFPJAy5tj6CdLkG6DwgRFdryb0r6mWruVeRE5Y7O0bLefQbpF
iII4b+84GVuDkLnhszCAyLfjjyOuwHzwbrPs8qZoOFZrvacwts+tO8ub6choQWesgCkRy5iuBSqv
Lp5XeXWi2UzNAVr1iO9CSOQcoXcxFjNbSm6MtRPRPjsK+iDtCyLQV3mVNHfICMx3hD3NaON0qVtr
/WvZae90hskNAviv6j3dVlaz30QXMb+93mfmTqH8SP4JTgeqjbe/ZAbCP1yNZVngprE+tlX3nZ2F
OIdZHsbPsIfEgX8VUDRl0o1EBRg6sfYey1pPOlVHyriXmbO/woHYdeRAsBUx9JxXDiq1SqmuuyIE
ImfZFYJch9Ng4fFrB+reotmWM5VPxhkyWFAJqFncfDxYmBS3fg7hAAsPBHEgL9q1QIxwV8Z0Ar5M
ePA6VXliK/ilP1R7CqGSzdb6AzI4Y53wrOqokpjHVdxLi/+qw/FxD9YEOvgvekk81RWqjszA/dV3
pjIO3Juu1dE6SkbcGIJmIyXhFNneBuschbssM+QgNne1ouWGKH/5YwOmkVLGlFruMffiP5nOJ1H7
Msv9U1xFlvLuudaM6vqPmtJ4wo8VlZEZMQteetrMVoVNQ7NG1wJoE5HGASDZmv6QI4gINiNJyXUh
3so18gkQRXiXByyp3NuYh/bGBXFgo8LmoH0E/lXFx8z01kkMtcYm7s9L3IgE9PWKhFCs5hibvqhf
yHrMzNtrru7E27t5bIFcwR+ZGTmX4ozzLDlXOZ5bFnT8kQmfqjGDtAkGG/pNFQqHHBxWOOlsOox5
S578yBPM+5KqlaZH3QjljanTADLpTAMD5YPKN2a7Hb5aMGMqu0u7rzGTalbcQWb8e99DIMAN9LMs
2FG2LDgwNREXt5F1jxO/ccxOwrOKAH20M05F81g5gyxQiPnyxKOHiudsmObISVhggFMlxiDLIiE3
m1U9MZS2eEYyvt02B7gtUPJUlXov0JkaPF2FzEw32c81GI+Eu1SXDaQaaGJ1Tzb3HhZ7rlFJTRM2
tQrCli+m9/WUMFQHUCRagr3JpM62yr1wFNqrAInnjFWwfONwpn2LgBZxt85LRJp8XKe9dJiAdAtv
QaX/dFe+elzpnImHmgulC+tX4tUQanlrs4RcEUGU80NdF9H2PqAsbgt5D8pHJXDX90/MRE5fxivu
QSKjwOz4IE0AJ+8lAeENgslFJCwRWlltCb5RmYzmjsfW6oicfRkoWdN6YVSzIZnZKn4xmad0Acjh
6d3EiiimiOPgW8UHqw2T4Etj/nfnkbXTXH++tK96kcXnRqG5mBmjDd+JLWKVJl7REg16U8jBIlU9
DToed46NGBtwCwNM8pbo/lBWghZh+y8IGnugb6TVrsNv4rHdmoBHWLX7j7mMlzI+RRudbLl7fTgF
uOvw3/hrdKszWl1wuVut+Dj6z21OlQGtrFkRvPUXyLYENUgz0Cf5XEO/KL2suvgSrusGU1seg7fg
MGd58gyfYmaPV0Pv1WATGYlpUPnyoRNBGKZ3HioOPZg8eRA1NMvkL8+NubOgGzEVfC4E3Qsbkddm
JcQJI4hH7VVBNUnhtl9Z7lClfqs5SQGEwXMuv1QfSMZk1THCANDm6Vki3/KYOmu77kVX0mXPDL10
znobg8U3KTQ8EuA7LHp1XAzah8dYVaMFjCJ939ECBromxVHvPl0C+vT0ApdETTBIxh/6gV0+BEdx
W+7jx72hXJLMkTuxG7i4i0TgQb9nAohm13qo3m1TWK0QCFJlvkGhGC6PxLnSSiJ07r/3/EVvsKh9
O0YGNysAKMEbQBpEuS4weNJ3bhtDRG5r5w4GbKtK5AL+pHNzj8LbafOrAbgafh12NjOjJgKEJ42Y
tsKUm375+GMok2t6DQ0fV6jmiSc4oP9atoYgtmgypJsJk8ZVVim1iqiYfegkkG0Y7EI9AEzF4uVL
jOLeZB//VfewaROTXWSChI+ojP3OaziFBM1d+nm83wKGHb5hGoIL98uEC4QLiz94s0do0VFVQM3E
fuy4tgsJE73hOOG39+B75aMx0pdjXKhrCRKG183quSTeq3UA+wHR2cJm0YfZauBkC/IiBClIBMgG
1soj3MHB07EOB7tOQyz/bK6l4W2DAoFqtWbV5D5m/sDWE9D2YSEcDd7F30xmSXs46InnL8UVyKb8
gmEeIpjaLkuGyi6wKUq/3cjceZnrU4PLZdDhSwuLIsLbGn7oar7aMdamFY0cdSo9JAHjwo9++IJQ
0sB7ZUkKOES6VxsIEjmcgGLGRkYF4747bLaQ7BQVcScAeVEtoznxxmYl5wgl/WQ7WFI67A7t8kRE
Y6+crTCF0mtpxbJSjYfodGRdm463uFZ0OfxaXkpHEk3H4qdD/2KEV1IgsE7FyCxWMBq4IYDXE5bJ
z8M2nR7E398vVB9D5Trr2ywS9TnJLqkHVLs2aRjYALLsEVjsEmpIDn57BZn7Voj7MrimaZ3aSauG
az3orpkn72G/ec0ctrP+z65Zr029AX79ya14VtYOl+//l9iM+MyQNldbejoOakdwxXa18FIDHKnt
eOTD+KezWdSHLtkY9T+Yt9NYMQdJmPfiOn8Tk1l8EAmWsjy64SOXHo7gaO0rBf7uUCLIUOu0iXZa
lRoa9nZsxmpzZQo/UUm4y0Hxckujs8GpW6AEH3R6dl2vkxk9LmNSFYg7XB/WIS6wnLeX+en6cOH1
7aQR5fs1S6KT4veuaYiRZJJSdN3QbPonPyyiYcrDToP9A88+kWToIVuaQUpUKZE2nU5uG4yVPd/w
Wt2xnJUzlY6p3VG6O04yhyZ93wfxdf4pXn83+X8ml92G4g0aWmegusJVcznXcWCwlNaUl14LC1DT
pfONCBJQ6YqRhTjKRFY/WdorQicRJISeOBMxRgCPI8CyAmYMrLHNawxNTTz/b/RrrKT652WB64Uj
DZPU5iSa+gjZ/XoLL8FziwbH/ScKQUQYfgRedxETA4h5zmNnXhIwYsFMvFE7sTMhaSHMvOMEfDWo
Va+U4m6X2FMJlFHhaqjo5VUxUpLULCkuW465MBqLm7M0VAbqtT52Mpmz9hSit3MdE8AqlREPrema
z34SNgLSD0B8HVdbywgfDxMU/lHSHAH2KD9CDJsHa1aRTfjoWJmyVIItVcVqW1QTsj3fI6pWuDQe
xnyaEYDsz7V2zwBo/qrOmWGctXQZb6QWKnzq0NE0TUM1kbG5iRxid96zu20CDbViLUDOaE9GZZdH
bgH63Hp7VhGLtmFCDyS3heKHq0lYi4VIMAbB4XB5PUbTPpyv7AChm6BcgqsQE+mrrFlhcTadp9lR
QE7uLwdXejVkLNGgUiWRAqhasPlfmiUvfSL4mugoyB2nWD4gaREGvKE5HfUNiOcGf9h5vEpZC1c0
dGTFYSIduwGKA0cA/1JL0tipn//nJL9Uq3bAEvj6mCCEZw8P952WlT+HL5Wi1ShKzjJlQYL98EsK
4PvavexH3tpGw/BJt5dUqTcuRB7aDLsA3w7BMRxXfXDuf9w3rj6nf+mpFGpb+d6UM1Uem/t3KShI
ya4nyI7A2YC4YJGAPqvmLTwHKU+x0mFQT8U7RVvHqSm4pxbGJEkQn4gKHn6PH7Cpfg8e6gmmzfBQ
ulMRhOPTmXq/0qxE3GjJ/9MvD0RNBrFD+zJPQ/DNyZH/wf06r80OnCa+HR5GxQU9W851g4kYSy4S
1SzJqSQoK3aMiG3G3s6nF5KQD72IvZ6CHC1A10skBUOLbKMzCBi+YvxuTcTIP55ZBMEuWNqDqUvn
Yzpc1WyEqT5unqdBoMZchs8ckB68F9/a5jGQmXrHhouc6Jf7MT1wi39vP3HPUVa+cWHkteooEnyT
DgGJ0AAxViQsaJJn0IQonSnptxOUH6Oc+L9YrqYkU6BOffMAd+6AeD1XigcUO4LTgPAXkLDglpCm
wdN2Dn+mHXi09IXMThPPxWva4Dup87TE+/kbp1vxS/4nGqrTjqDCh4xUBeL5fbIS3Rx24Amyq6X0
zBmTI2o3HlI7H8Stm7aDfXlFNW3IgzCDZUcukHEF5aon4kw/vS5W6jgcpdYyiJcGtA7DeXrGf+aL
wC3sAFn6tQye22WilHoMHRZyi87UYb5k1aAWClpDbw/gzinwbM1UySdRlPOGRrwaqwp0YNrvIgJ+
z7kCimAWNrEAI+8IKKI/2mAfz0wbqASIz5lKAZsrjQzOaRlNZWZ6IZsSMqVgEpKfaRag9Kp5h2yb
L+kIfPHWQ3Q58Zas+dp2yyoIhjCMnXXiF6OBW9PR554P7+KV0u447nXTf4+9C6CKOe2yCn60pJMH
1H20hiD+dxUbTrh8qup86/5Zv57RTAJl+axMsxXaDOOu1kOAAQ3+PHX6sUlQWE2H1rfpMueww/1G
wNBXU2p7U4K3HCiXf824HVfz2M+gi/5/dN33ZzPYB3KD4708NsvkzcggjZOPn2njNfHVw5xWioBY
JhkFOTeyAdRLFf654mT0Sh5eU3gNuu/6Upj0jZRM0MMsIh/dStBVK3b+QNSEgIHRODSnbl/0eMia
jPG0rvrkzMJFVr/cxVwYw6KsriwwiGQb/+ViysEs/yCLhcTkzGQ/S67LVHJhLR4cDqBG+ngZoseW
FjNdmLnk+GZNEMFzlwKmiCx9LeSnfShhgZ2wuA2IT0WSgbaZUNnw7Zxyxi/+TdQKiTa388k/gTzJ
vch7a1A6+CXPYOk8/gBvgzkD6JCOFVqU5CmpIgWzf8Jdn0LZvwN1xOn3VaBbuKIS3jw8EXylVp8P
8uEfv2xLdTB1qNmEsIqO0PLuRs4PE+83dAv/uIfFZlb3jZI2H7g1cLxxkrmLd7enVgLu2UQC1shA
mp6+z0R/Jm3b/LbSo83Mk60h7ZcrW3DEb280xvTlQx+Tc5NpY4Hn7syQ4OsfHRS8eH83ChQkj5GC
lsHk2uKAvFElNaRRfe1Z4Xn0zHE5UepjE+Lqwf6w0uisE1dyYqeovBVGNTmFCq+oUnjw/i/zu85a
jgS0qOxfE6LXuWGu5LybR5J7UydIvtWtWWoQqx8rU9SfU6j3YburbJYm72js8ty/hCBhUErfE7XS
VH+S2ug8uLR6fYLFHWpAemmBHbwvRkkESD9sEq98WEd5xR4auUgYjo/WbHO5YtwoZzXGyVrDJZsq
yYMf6NxNLirq5cCDbwTB3shYH2C0mVmIJ7VbYUWi7bS4RrUc8rzUolvPeneIZh8+HMqrtOdKGw9s
FSEqk5bKSx87Uuhuky5uFj0piYqeKcOHPu2lii+1R71ZgECwb4gxBUqvtaYR8LykCtBEGMx6+CUX
WBXez5pxd1aDwSPH/fNA6bP2o+puPl+uiz3zS0+pHscpB1IGs59jw3MOnw8T5W4B/V7F5DJ69vX5
Txle7Ieo4vRWI7GirRJ/nSw9QbLNnZwBVEq653+bolqJP7X5nFUwPZUzi634gNsyqeuuJZnw2rvk
GFnAiZo/AIw5Aebb6UrpiXFMhO9q9uptcX7znBlLtiINgqJwAa9UGsVYcpF+9p4i7zLLLRI/Zku2
USapnAS7xJ7R6DCv4YYZaUgl9NvaIQTfUOrI06F+4Wd3S5l+71hmmo3LJsPYsp5Jnb2eJDeMw+OF
vrLrzCNIqnH4BqINliWnDYBvfrxttw/km1D0vCjVEzulWSJEZWmkwp8TMt7YMk6EXpa9v/cj6c6B
0n8P86lwYM8FKX95kahkKwRi9kxz4/cSIElNJBva3QUxp7STjoQ5ggdHoqySDgoHCAQBXf4j/C69
27WcCCfuJJALW3OBjcy91v0EU+N7UXkI5wG4AF5am142YRVZGNyq5x6+e+h8ZAwOSidyJPyNHdZ9
PyrdYKPPUR9Us/FnB+A6zHZUHRgDte9qfvXeDv9Xe/SBzljkllDyfzoFO0ljoLRGmC/XYYYnzgrS
TIGEGDgjlysooPREbQYTLlnphtV5xIV1Bs+bmCFlot4ef2l9Eq77c+LYE2HvDxkDWeO3ZeWsVhnA
PNuyFZzj9FJqbUX6fV9KSmF6kq15imL+W6bPN8rXUdYAqX8pVrmLSgu6sY5e7XXYb/VhWAxznei+
gsR4s3Dmegne6s7F55lVH7SSoL1wgdS0AX1Vy16QAUhMuf+vbla0I0j1/ZXhrBRDdAaf8csxzl0Q
oAIIrHK1bX05yr/gQLL/Te4GhAvwKv+yxtBXYi0PYCEazLGMHpLhOtSEpfw8oPUjJYEvU5sv5z8K
huJELx/Di6LrdUPYuV22ZQRiuBNDtIzRvOjR91byHukS3ZegYmQ3wgbzNNG96QJShcB9qPWVc51z
+QhRSTx6CQ8r1Agta+WOEZDtNl1/JO8bWhjLKhGjTO2rGVnUxizrvbKzdwZXYAWojeEETI3JqQ7M
+0uaoJAthgPwi57ZmbAyfskIKcK8zVoRNNRbcbFQbLn8peCu6qZW4hmvJ4IKT2LoaRNHTWq+AaHC
uM6aNpDfHnvG5XjmxahMQyD7AADr6bFhcFOkteE+/P2BTnOkReSW3SlhiLXxrwdmQevx5BOyGhtt
v+f2ujIxeul4KwcEhNRaSX4Im9rl/pIhWGxdeDADblH08eTxKGTOkXfisFMorZ1ilwgLcTQR783e
OiuCcI8CY+5LxzzPIK8hu8A6lN7PYXjCx5Ol3x5brr4aPIR6qGFbBax2zeU+X4oBrdPLgwTNq2hp
QZLFmpyvPccRqxS8XPPVRznqUwIhc+76emYWQcBJuXh4cdwxnm7jS5n8oxUhzZEskmTiTvfQ7B/m
AqTzEc1x9DwmBVZ+XQGhj0C2vBLKy4Edkx2Lm80xVh7MuiD40K3oX5SumGwhHeGL1JnAz9H+5JL4
JfC6ot3AQWdVeGOG6k7KF2obqj9KkHOjKE39+d7ZBWQQpycZe8WleWxzJAaV+xpQZE00HXRmOwL+
Xm/iDKclOZLQNYxVjc3dNpcnb/NXcNg0vUOAeKRoln7P9G/6hSGOTd0GMO6c5ejQwdg2ocyHIs0G
/emCIQjYGwKNxxqkZDadGxRA3FTpE6tCWcWUQdXtnPJk9G+gV8QT3J6XwdzL/1jHDkFwDc5iItOu
mdASONrl1MDAeUvucKX8N7PmPx9axUfd7Dh/tjuQ06hyfDKppjUMHxX3+pN57rAQ6krD10HgNV21
rByBKD26DyWOqBm7ZwFZE7TTroOxPw/seLq/hRenrVtqpKHeN8J2WjKJhtANCLcF7v1z/RwdUuG3
kw+7UQzKxRZ/yK+kGYbF0KHSzbUsuj6eZszEISRRyhjoixyXi1AQCieh0DTXUTRZnNiF+zKpbTVy
IDMMNvQ/c69PlFPoJ9rk8UskHej4yts1QqYINqoU2GMzlSHp+yk30NAbFV6J/hPMdRakc/EkGZeH
7UW5s+KJLkKIwOvxxPGLAByWlnjsn1iKdJ7WcdND8kGyPdPdHdYMbPLx/ehnQIAsnKdc5klncfLo
FMwDrZ08xAQFi/91hz/AvKXDej6Agwi6LCWXsZ1EU2tSSrreKcnVwiHjN7sqozbMu1GNZLjZKOnN
MQUUEsVGjw/TKuqUtoKK8N9XDwFkpcmASBDcz97aoRlgRFWzwBLIY5tsu/2xV8VEFsARiqaEZvse
zFjTfEBPIuUQWy7qkwZSfMQsURqnuTCL/b2fnjKK8p9QYtEUSCbNsrMhG8nYFiOJGT+KzESu9Dt1
tToiMvfO4yQ0eOLTxl4XAhi9h17leJPolAqgCvQMJ3Xj7pcKFjTgsWsJ7N0HdEm+8H7aCtEA8Cj2
+vCQ+iO/QwRo263SKhUtKKeXbU0KQe3C/1EUOJMrQI7pb5oQKmhGEUl3iXzdHzZUj+ZXwHISPdkq
0nvn/xvZEJSmMEAxZS1767V27gtAdWV8AdB8W+D+RAnuwENQKXL0keXBr2be4Tr2qehEZHcE44sB
Mbv7PhAB7bn2cNFHrkK9R6u3W69BybO21FL8BP3NlTX9bAHTw2wFAuAEFtHQqnKBagjAGktf6f6H
PgrbtKb/ozpGwbT8SDCV7n2p/QupnirFda1E1qhQijcFkDRnC68K6RTIw+HwpSBMadu23LrQNVbQ
ywT0Ve5fVMYX4tsd9aPIjs3LZjoKreX+fowHLdJisFKt7zI7F/mL9r2IyvVZrWkK6LMquaBrSU8d
bS2MpY5ez957TWoPFXrwNfeZ0AokaO6EDF3Ak6awGP3km2B/3KI/hbirOMMKc6xRwiILlt1j/84f
7EOCTEw3eyVG/nwLnse2NqOF9e3INdnXCwMqTrADk+gIttxHXRmoBqPUA8FesdTN2ve9OnSJQLzl
o7v5Xrex/JajynsWLCOXv3LUV476OKbWX53kVj4k2yuv9Mm68+6S0AWS7m5ubvIRmkPhW/OFkCDJ
KQpWUMu0Lgxg2b0S3agwfeXguhndCvcW8imnn1aZl8F5/HKe8HWhT280w+/U3ZCz3abfMWZe2D5P
K6LjaE9KV6zpbkzUj4dmkZJc+AqRO1yADHsdMQogAgXokQq0cAJQgeAEAtSKVH8of4Q0seAkhp5i
KxH9IMIw0V4pKH3B2YhzTp6GBu1dwW8bkmgd8nd8j5WxPFNaYKinshN3i8GtcCHyv5knE5zAtPhd
2e3cXFkXC0SQK4Fq1/7ia3DaJ1xFnu/GWkjZXDnrD7S6YZHbevpW+NKp99Dus6xR64SJZVeoqkXS
4UCu0g41I11HVr+rX0cuOx9mN5e0Og8yDx3+prYjWNAw0Auqtubo49Hd5l4i71KhnBU/nWoKygNW
67Xi9bxcfQAxrT9cvH2Q4Z0FJK63qdwnI9G/2Lu/lxmUwkUr3LX52d2qdvLremnPr6NnbbvbUqHa
X+Zj2yv6wA2VwF60JGEpy7P1VMAyZQhWvzJP7pV9g1kUJMj4Pz3iZqC26QE3iXltLIuzDwdR/8f6
MiTQAJcML4DMx80nBRQYgftVJIzjKGRocxB4oXHL8GV1907eVGF1UEHs69TbF1YQOuqiPXc/un3G
e1/xuWKfj5g3nVsuxxJqCCrsa91JmbP7u3U3Omr+fA/5rjG2btNRuGTJSUB86bRi7cHo6JrqX/Yz
s9z+zc67hwF1U2TPYd944CtyAZSZaZu54n/Pq6yy77SA4iRisPcQ2neFZSFhhkOyh26784ypkL2C
98jGOBeKi/x0T2QrFfzl0z3LfxIIjVGxSTLQhvxpPLBRU+cbpJjlGnxHZTUQ6+gP/0cKK467Cpxg
XDTU7ihDJRGtKaSLAoGGmCNKTnlvOTBUUM3CLG0PGWSEfVeQ5kk3YOO68m8EWjVsH+Q0HRKPFO2X
U6K3g9CPl5hIdWOAEa5WLhvPpDidI14j520Eh6W4fu2tbtV3NhX9RCf8ywIWnser6tGCndo2n2Rf
Vmyp5aISg1Nv1Yh/r/QIwaKbHy9dNgf8wRQPpC3lO7N1hTD0a4+sm00IJXApHh6eQLrNWhBEJP2X
EYHkTPhti74GrEQkvEBiUaQOdOUuhftJDWzO2wwS/L1WmDREU8P+ZXjbDs5RRnRSQ97O4Gt2V+Iu
rIGSUmh+vpInHY3eD0H8mh9Z/Jbrj2VcSoJcVzAaqeSdzP4SuB7oOl3ztZuvgmqu2pXi8c6r89Zt
N9OxfgKWaHKUdFehEFcD6+EmDyn9TZFlrH0Qwj4wYKUlAmkZa9mbKoeR5693WflTzC0CUude5iTB
8R2j/RhBQ+ePx3uv6jl1wa/djhFuH4YBr55E06bv7wOmHg2ComdKf+Kx/deA0mCdem9VXomzpr+W
eystBnV8kKa8aCWwko1xioaNC5Y2UIQA1HWnqJ0VrhsBn3aameZoUmHvdkqYIoQTzA0jsFjT326J
nbdnp/PydtrCgPYxkuwComXdxKsJ/hU5B6X1DfnbxDbx1bSa9pIPzyIN5qOPhX+6S0DYecHFRhSS
ICncnj7mEiMVAlnO7Se6iF+ABmfh8zBb2hErvec+UEDkqcaMIhYEwxfzg4pAypttDXW+i6pvg4J+
uVX4+WKZTVgDnKb0mUDX7opQwiMSJFUmjxdWUuDFi+jLnAvKt258L4UTQ+z/WM5cMTmBIkuTOav/
UTAB8tQwEaWvL+04Pa4T6ToTDunIlT2/pwfgX7NNloGBjvs/sAag6SmvI/HzcmYQBh9LZnxIF5Xq
P1q6QOQNXoNvskJsLakO3KmBkSEAI1EGX77CXubbY6a/DAFVjMv0iwaX37/6WB4uaNe070ZqVXql
TIJF7UyuMTsvSoos4L0Mx3iNyko8DwOxvYHD7Q56XN0ZmbKICSDijuy88l7hoyY3HIaRZ6KsTpNe
IxhdsdVDJ5z0dtW7LXfzoV1TpwHi74eaxnMdykMwC0N1DlPeb9k6YhytnnKJLoahXNZQjkya5qcz
TA9ogE8n6jsLEu2QNXKKEjqm/nRld4CtY3guaKKE3lAxGLWrzxZ0nVV4BD//50naE3STrW5e/3q+
+gGZtxddbl/bjWvtqLK4ccZe4lw+GRBFsIqCMc8WzhRtROaiInUWovM87T0etR4SGRkq/J2pT+YN
/8wDeYraNyh3YptYjoQn6/eKdkBfn3Y/xk2DU4xqUHJJkBYAqPjF22LrXTrS2L0QjbSgEl2orRUh
/E2MSSQAJ232S+atPfGMHnUM3bowkKVAd/DJhV7l8YZXE0eP6h79szV5qmki0FyHgVBPpz6VErZL
auhpw8H7Z/Mvt+ZD5yHQRCTUFf2c4pEOGffWprOvg16vq5heIrepbiQiWp8a2P1EUoWsmNvTGpp6
pxhV4zShlAhhfsMIdsj0C8HvJxdDITmyFMq/8u702lPMl+H54CFiOpzWds1sITj32QmyRQsDZ5TM
XRRpo0vGkoldV9adXwv2i4o0zJN2G7Z6td8G7Td51Px4/FzbkQAfY4WN5+EY4riXFivGIYfUUntW
xR9cYWoZCMGgXVQVFOcj6/G+sYRnMovOQAcgMGvlRRUU9LbSduHjoiOAvZNJ8sQS53JrkENK0Uf1
1BH0swHh1U8Swu4DucNRxFWe18g5q4O4SXQwkjdyYNVN7EIv7XlT0FxRl03vE+VPxyMq2v/Rg27w
JIpv7POXMiMEDlRO0p7qqVQ5LmSLkHmYCGC/jW+nYxDwWFlgPPBMrSc0BL+73xj5a5sJcosGvCW/
eiQE9FZOAMYSNvOMIOdLseqn2zF+5l8EFE950eRGRXBHzImPb8NN22Yi/4kNzygweS6zltEWmmKl
5NENZLW9BNv0yqYaNScHvWiyB6Qu0Zb71w0/8n46ElQeud2IEaJCzDbR1udYpgRSUFsnNyn58n5w
LFCZsllO1lBfZef3lP0GCjvrwvzIcV8YgbOGAFcuTCZ814Vdg7UY5hRW1F+hvANN8wezVqQ937p1
7jiEESwXs05IjZ05+SUQzkGOTRya1MYdgaN0+Nt7bJ2rv+mOhXN6SVVVckHrOqJMooeu3Is44rbv
GAEVfFWnHDa1SSb01PACNenCgY1dh7tb6BYZ+6lIMHMDz2sA3eQmvQtAxwlDvTZjCyIQDk0AQSwd
+LYaFcF3GCk4kToyG9Y+MEUwWUB8A+DIicSvyaK2rtaU76kqR8KZth9VmyX0qB7xc3+BaVse4FeL
td/u8180P4SLJ0uDnSXBNlF2/xLMlyz4uvgZas6qHJEgh/GRXLLlKjI4l7be/7aDywKEXIpdxm/u
dl/GNMEhQmxhEH+VLXWmn9gMSkBShB8RWuKu5yov1Ype/3DshR1tmyg3+ukuNVxZzm3e5/3GHGoo
Qcc+p5P+0bPXKiMhb35nkNhie4qMmdll4lkrV95Mc08Evh8fd1bdC1sq/c6+Xtd1p6VwAKxlE6Il
dIlV3d+CNCLd52oYsGDkSP1otYhU/FnFb4lt56gJkdDizm9bIiPd8H7HYowi2zNxX0HJrw/goq/t
EJlKP7INf6E0H6rBRmhcSIRRihIjUI+PJuIUNngKeqtoIPSS6aCt79vX+IdLR+EyYXuwVJABrbx5
DS/qPqVZrk+gcJ9EV4yjhs70WvgxCv98U5dOONFlCxhmSp6UvKTY3ZoTB4CeC9eaMZ0TytjKfwWU
nsd+qhNLT5nAwGlYPWHWp8kYcy4fx5TXLB6updl4Fpe34k/gih2P0KZnM0rXZIlaEgx64CF+NxaU
mKB8Zo03j8B0VdrYypfq9XV3kz3r4m0mcLBRtyhJDajQfY9PYn2N5W+4KnANS+Zb6EEWPPXX5krM
O5og501WkKSxgJxu9PGKXf8Xx3j4uqy/Cnj+Wptiw9F6B+bexPPshPtrnQVk2is/n8qx+UZRt8r6
1QcB3oJZxX/qjbffDWAiATkiHEh+bONPE5WYGt+6rHS6aMGWTfcB6EkSTjyuJuYQnyVmGMGmpQjO
5VveU9DpJI6PUl+MBwyv/WCasazfTh7mdPOFXy5relL0vOO7T9aflfR/m+8P4tD663aZO5b4cTTO
wJmw3CvIEMbHtsZuhxxMfjmGQ3mqdYfNa4ZFNjQ/sf1BnO24hDxCvLAf1+B3weOh/3CS7HO0pmPp
aKNR55Qvs/Yg4RQtuAEHhZTf5dpO6v1rZIMAILdgeRAcQWt1b94ksrsRV8lRtJRu0I9250HOyb01
BtVD84nLTFYSjai1AJF8hsdwGxC9T2Q+m7xgkfYqNZbOzOckfEO+6BZ+730QjxH2f4zB/avIaTtC
3FEYohlryzhQmz8NmnrLcBGbhh7+RqHWiAgXTfXRaLkQFQHORFVvWvmsg05Q5gZozSEu3AsrCdMG
7narGf0c+he+S9ZsncE0yK7oaX3iumFY1sd2/dwFOikkRU/PCCtLLYnBSablTjn7r1PaAqU/coTC
++DrQZOosdMwsvelYvq0pZKEHnFPVrrfwG2+ITovfZq9xMK53wKCRHdA8RWwPypUY3l7HtHxDZjO
zV5VkHInhtP2NqSg93XlipU8mbGy0GqwIF+fID1E6G0s86N3kJTcbaPDvZIp9KJz9/PnqZMxZUuI
cQ76hfapQ94NjqxxGTXMwZeFSw5h052IQ7IfrrE5xJt6tlMjAnZjH9x9uENr+sME5mi4MLV71TrD
HT6gYlfAaoYQL0trNetLYwMV5J6+PDLJzCUiB5k6pxvjEDNzZQMR8TcPV3mtKGmX7vc9ZpPH3rWc
9/JMs18MteM4bfHx0068R/Uh0OSxIqTNSLsFvTkUImsxOPmwL2iaL6cbNSdWUVmlArsmrLxFrd7l
trKm8rYBoDTkqqd0E5RTUSe9MKgMMtByIrR9xrz/GRmdxaxNVrVDfCLsa/t/OHslyksPTAvJvi2y
bbg/yGD/bWe9ZqgwqAbyiylc7cE0c2JseZz1cPoVP6qj7IuukNQgdMxfLPCO8v0q8+kdCC6e0IgP
Q0UCYyNSbaPTIDpkz5DwTS8+eJM5lsP++oti4PKwXGmRvOY42TrnvgjsUznWLHvEdv06FB6I7xRR
3YbRhntehTuZ5wA3eJb4lBwITMw55Xd3KvkASSwm9HKRpzjRDvtOoKoEQkOS5L1Vwqk7npiGzGI9
cR+F5R/PEvmLP8pipJAhRJJGG+lPmK1GkO/jbceBYZmyMP4XsW9jrT4v6G13sXZTsahiYcg09/7B
gNOZiOAUeioRTUNiwxg97I2SOyRumJsxcDGkkVJdpGzp1K0woRPt1HsppwRKCsu6mD4hQuHtQUFy
qacD6DprjXoYtY7nS1UExAtS/m3pjILJCR4tHjC6DpXAO9IMbpilifCyX/G0v16jygg1miLFU5t4
d5e1Ydqz1XBsp+jEu4S/NjEr7GZsP+0y4uBU/fO9WZOuvASTp1ALOdsHbsKMX59Kx8db7ADnwNdW
9euUBPFW5YqdwWDz6suUUqgJrT5UqAxqYYgURoB6e41UFkrM3y/3SrxzhSm6mf/cV4DtG5ElEno2
JzHdM7kSUeYuwLlcV52VH6V/9gb7ErNWcZnsSFxAHvBVhdNw4kQdRKYbKgVW0iJXhEibHUu0IHzi
jfARV1KyQC2L70iGnQSD1SqCzhhUgCSm0WHtb1+sH4yrDlboqD1IANsbaiP+f9H20/XRnb4h8kuF
TuViKwYZnKYeDJTp3g7EiXAoS2DEjMOQV4zYipGzly/JYIChXg643KUR0tBspxsR+3Ctia9cy/oh
zTEWG/PberLWwHcNVjF7HD4m9us2TNvH40g0GVqYI77aAe6jGL1lWozMAykScNqZ1Mvonu2DRtAS
9NdePixB5WA2E2RTT+8u6YPj9Ok6zRAqoMyba9BiOAadN7zMg4KBO4bg7wmNv53ML+QiFy1gU1Bo
D+gdI+pvHqbEnQE+WhY4q72OtRo7ihaiZ5Q1Fc7uZxeKoS7030z8x/XARtN+HUET1HMUOAOGTRQs
eil5yk23zp6wRH89r6dTi3d7B9FH59KBrIKLITETENzNen8rXHhM8CUxmL/JmF799RUWBWfZCe3w
jjERpSc5tfNvTpyhX2iw4TWVhKtjX8QeWqMmwvmb0ooRRqkeZkbcEfAAfSFx8IAe1RN/hkAZd/jq
dbIBKVm+zI1OvqpvzEB3iGfl9Tu2SROTZuk7A4viEUFuZ0NvCxfdzC4MNV6MWoxkhcrlYkPQ24SH
aZZFm+vx/0dMiq7WTxBBcjVPFxTgNla4JJqeXM27sTT/NJ1uOHYtKpG58WdKrTwvoGCDRZTJBdAk
y+SBHcUE0ABAHnnbevUmHX11H6vP1j8EIU901J4GATrGpui0Gwv663EMGOhblUeuT93f/mEceu6y
yuc+BFOajoNPWujLU8XATRXzjFugitc2zwJ3C52mfSd9f0kmVJDG4/R2CNmZ8o9EC4hhHKVFGyEx
k5Gr0CzYy6EDFSHDP3dqxf4JPqyHaYA4Tt0uBrav3sDZDQaLXU3OF4iOvQ/iYLyZT89JiwXXXBRm
lyKCe9S4yeUVjDSNrKi5OdnMkHnSz4D7kAcDFzSUoNUntz5e3Ks5CFUCmbn5bqR7+STWzFnDGNj4
KUU0Zhnf/V6mb5W0mGABlSFnwzCKhhy7nyKiGoQCTF65DzEohqAMdYStq0ZkPIn1/9Cx8XtXHwXO
vkxD8QfxCkuOHTN4DhbHPeenZumLbdOfx6Rt+2CTakOCnGUv8z/iqVJ6fhirEWbLrQrv7NZI60NB
58SjmO3NQXnYgXq7ML5LTAlvwKPllccF8TZAK7L2gUxVE3m6a3sgeiL0plh3RGeB9Glb+sdKtFB9
zT3sviZZKnF++Na1j1r6lOxUa/EjT6sHSDlLqWGy3OuBUG0LkeDVpV2wvwp7ZCXWsbipvDQMT5nP
n9wZv1Bze/6/7GUJbVpikCJ6N09bdH0AtjvE6Q+o+LHqoYGpnG3jhVdn0bbnTG8gykbzxxYbtK2Z
oQ9RaUYH0FbWb4ZM5tkFUq2sqnHSNYaZTtMDygm2Gq2fquNXGez4UgoZG7eQg7DKhKOMDY1FQDBs
6VmHsrCy9v69pVjAxbHI3LBNxJcHNNFJqm0lALX+9dZVGn/BmOE9+ZAyvE/854VChgB2EHdb7759
TJeDuIVLaJema++UOfJ4enVvNRDV+z1y+dDuapUKVpoUr3XIO+9g20U2RIhbKZSqWuE+zzd5HIom
5MeMvpyCvRlCudAAPxYMZN01yr95asxgkwBTx+aZX25lYH+GiMkgnDExT3gammGHNWYhKCAtdr/3
skIb1KLpdpVgpPXw1dMtujLdzkkqjQQX8qNZaGQlEjc446BIwaAVnFODKgObrzAiXDzkQLBt1cjX
3Vct9AAs/a9juUEoVRAdaHgpDAe1djEfboENTTOFsU1s7a6umklApSYXznENSAXsShB5kvDMgjZZ
+dUXh9AV9ACT3c+hiLxpuWIqmJKEusky3GwQqqaPd8hc+jVFVh+9x33/0+U07j1qFRevWyDPF97U
7apGx45L0chrmfen7znsACnxf+zHDyx9wCEvP4p92s7hnPqm5TAXYj2m9Z9vfpwNvjyGtdzdEvbC
ds5geCDjw1CuLoTTBcd/r3PKu8qf7g9BKJw0AEjl/7P8Q6D0YPYT548RwDfMiczDaQFZk0190CEM
EQU2HtOlYOadE8lyBJWpb/fi7ANytw2Q663FF7G9nUwLooB8/KSJ46RRrnET8L8Ljb3jmzomQBw4
NWqoFKFrhCyD8MjC7ePIVDWXbTsg9nYnk7CWWl/tXMktAYnu/2F34LtfnV0PZwgZ2+QfD87k/NOB
+B8a8fh2gHhiy8GUNU8kbxiXs57b3imvo02vbPKauGjRe5VsZTAaBxWaHqgcTiX/urTxs6cHtue3
9iWa04ec0XM6qe4Vy36FUN6TMXjlAQOj9FFJuw9lczli2SIQxjnDu6lbWI6bCknhcYgjgSEHe2mm
0C7hQtSeX4Lamt3VJ00c2jl6B2cuQ1aIEddvHkOXKz5y3MAaS9duKfwNKUYPjJCG697CIHmasbS2
Lzpa4Z2TBI5kxK/l8XF668iIDMAo/jp8DviiLMcBtD36W0Bb+Grb3nJOsc9BzKkgVmt62nWLvzgL
V0Iv/mAC1QJayoWjCZqwGjQQBYqMHHuRrMj8KOxF9W8iJpmX3N+B5Y9NlKla/vATpo1PA9TdfA6z
1zZqFIrRj7x8zjF7s3IBrmrGOZ2mCjRFmvB7XmtS4D/6a05uxwUpNqM+EhAGjowwahH/ib3gAIRs
SPmilw3mcrHb9cIzKT/YkMEOoLvt4gkMm+03cdEmNbTAoF26s2T718Hb7KQR9+uHWUUUHjT/HiXe
SGS6USZZ7NaMn6jBqcg1UdoVBALr9MX3DPZginD/gVswj7KLb3NhP2rRcUUKXuD2E5fY/ArCtX1R
YJnSLxUT59MLEDOUxWvXeFncCfSewScHCKlLAsPEdMpiPJG71uZ6MjqfFrLatW/Ct23OODXMnebl
IphZ9bs4K4bQC5Ummm9Z2B5wEScE1Xg0o4JQxkbZ3/DzCsAidNAU4OkTePmZMXlzCkvKdE+YRc2S
EvD9JEiz01eTcq+byf0GOU4/M1sLm2xSEh8kplH0yLqIpYVRDeGc6vTew550I83kC3UkPiju9XRJ
dSBk0ixTJfyZS7TzfDM6H2338L/HhKAAxlPDK6HpSBzS9Ddboq0pEF1B5Y4jJBZkx83PbMJlhuZv
EaL7QVidlTGvWO0gWY0Z791ID4Zj/z1vXDSEeAS7RNINlLiAEx8m7g4POS18Ok868ahciI4Q1FZS
Ll+BA+flwrvrPDYqY9RY2sagG734Fbphe/d++zweS8Gq533JhirtQr+xGCABCByyjglvUw0rAKiJ
uDX5e7wAt5RK+WpEPfgu7ajBTQrlkFiQeJHmnyxVcMOJu9EskTbXTXZu+B6AUzrfWl6M0INRKfbm
UI1UNbIlpgvhbVOdiE2zd1Pb9IsRiIHjytsNDXKY8uFVNekJS2JA7rcWyDO94p+oD52wNlw8b7e9
CIcEsqZNlHnhBLs+TkJpomyjXRSyJK76ppMh7QZk/KHW7SlWzgI1yBVrAe4VccmEcPl1+DYlGtkK
MAHpTc4bok2Pl8MazE/6mvpSNvzBZvHkZxLJSjOG7e9y5GORc6ekEEVYcnyzs/lFT5qSk4w5q/at
id7/MMxpseUEA0OEIb4m7pICAIeiOVuhHqnkmi+L6FVq+gFugvqoMrqm0uVj20LcGrmWoE7UIHtb
Q5+BK8FnUnGf4FozwsOnbl8yJo6BvMX/gYd802RYHhQ3PYQ4P9cqIpSfaPoocSQ1NDsRDkm8m4Uz
RrLBp8DZjqFGW1jHXVGeyreJrqAkPRgL5gWxYAfdvOdR/JRwAI466nDZ25FRbO65YP+ZWohV6uAu
3OgZAxU+4qpLoicYMKEnvyeDVLL3jUZNYbjAXfaoJTN6qr88RunMoCtCwbjisb9s/Js+8ZAOgm30
75Yo/Hjvnc7gBvdnIoQz6SGORyJjrcWfGvUNjlacRIWsRVpZMqBWPu2A15s7JKEuwi8i9gpUMk1H
ZbnZsX1CVsTa89e1dm17d6xJJfvY8NNz3nOzV/gJSSs7bLtCNbU/a83PVYL1GrV8rvfBJhgSaZls
6ogwk2Nhrw4bm0hVsXJbF7uTQaENsFfnq9Nw7z7lfol4dSEb4Wy0Q1WiHPQPxJvxYRxvkqjwG0+e
/3hzabSEm1wQ93wQJ2x8EgjD3F8r6MOPASzWMhvLWTzV0XbUAGcr3oTuc2JizV1/3NuO5mycHhmt
M5FxiW988NEbJa8k97FR7yMTwgWWCUMQl/wubI7mCiRfaCdtx7E48La8C6fKQKzSuziKm1AJljio
bGwUDXA3P7dv0bhQnxjg1PCC6uedNx9NsM3MX/KRRTyhfzdeuqduWMh/5FUHchY821wHCxts0dNw
N2d9Be5Xby3K3ukTHqkclx7y2fIRlfPuRuGZl4nNC4Fwl7a9e6Sq2SE5VfRQYecsBxRwC2wc6DLW
AxvapFAaB5lqon3rHPA+E2IdIXT+O9UK8JpOiyfsJciviJqdzpFp9OQuYxYnGMv0FXJdv3mDlLHZ
a/8sJ/8gbCfPhqguVLoBLFdIzWBr2elMxuZ3AD4/ACt35pcNPULB8D5BPeoaxGvBF4G2RewWqMPr
PgsVM/URR09JVl83hp1BLJJSJQOyG8tJpBx7P107b+QgdbE2jlimvsNOJUBF+asdfF4JMtOIKUgp
bRsBg4XxTmFSre5I8+Bph+kh2/k+7DkhUNiQCCc37yCVpuZ/9451VFHrLyg9QzfLuvZF7FD4FjUC
dUgqiR5pfCWh9aLbZVnJURkgCWO1/r4J0Uq1lGnmnYuit8iiQ4Yc1Z3Zlt4CGeUUCtJ00CH0pJ1Q
pDJG/F2Yp7reYJEbRm2lYGodkp0J6Sfu7ilDu6gT9XTtUzbWtlFr6M59YqWeeG+imqAYyoUQrKa/
h8lrlwwJujS2Vf3obfcdH9+Z7vVvOdy7l3psCTJr4oG5QvAFoTd5oK3l44xnslnmMhd95rWLKU9i
zDxyYvLpPOEGeJX7jUNe4ynpLyYYx+dr9OY7KqnmDUM0sf3e8p8tYfJJH34mQorIeyifoqTrb6BZ
Z6ItNREUFe2umOkhIzulyvTcfh6Z8cfo4PyrZK/YCPROf3un1DeeBbSfDNGgulsYNHLtQI65i+8x
/yXLjuNhwm4GKCSelSchgo2t6ai72xEXVpHd9u/7TasyO1fix2FXMTTu/uqPyf4oVG8e+V5hdBlW
QajBnxtm/+wOmYyDAWS0kf0eE5lNNXhYB9h7SYkMyMG3xkI5Tfw/l+M9h9/a5Lr971EIGhhT4xrS
F3KyN4r0GQ==
`protect end_protected

