

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SFpyA3WDAkH/h6gENMNzEC70V+GWX/AuJRjC9uuhJRzuSJx7LjCfMePfd14YnV5eJpUmzZ71W3kb
9tnOI6KXTg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FappTG7uNGFdZRwaHkH1xaFvi8BC2aKkPLd6PQ4xkTkeceiv05HkyC3+B1zcjatywH/Tgp5My5jL
RzYpXDHCiS+WLEnVqDpcElLtP6A/XLl3ajXqKvZhmMUVZsEI6d4wI3wE8drV6caY5dK99YnGiCxy
c/wD5JKxsx7IEFSu4qs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LRNAkwpKrud10Lp0Eq/NqP5B49JnJU8WkULh5UDIksixm1tOfz3iui+8sx8gHS1R0x2iJMsSndD1
7xzPuxZn4a1eVkZa4n4EghKA1iQCL4jIUagjOF/A226osIvTkxPBVZ56YpbMiMwMMgRLER5z0xet
LPBfedO96PfexivUiLv1asz99hmC5fi5UUap1VwJdrnsIHsC0bEW3N+9FFvOSldno8glOl5txGSe
hOwrv3syYadhoBtySSxq9fjTH5UTCT6nikZqZkVb5yhHF7eaz/U8CnmNnm4+vrB5n+GG7KIVkI6G
7PqaCstXyxVZ0I0FOvUz/cqAZvJcffVN4NdFGA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u1B6Vk0Eso+5EvY7kmrlz1476LggIIsaO8lHvFGJ+HKHly0lYN/LsIll2vy/lYtCwxTSlrDsJgNk
NtsXioC5DfcQQ4kEDu1f339J7HYisXvM7Lhemt1gBNgHhAmdUioIYx0fpzcnzuhwqs4zH51jdAXH
PU3S8K0B/J5Gty8ttFjVJwRIoxIqhWdYqBDiUuGzr/SoWf0A03jx+7IJtD5tY/voAJ5g3LhC8YQt
AWy8nfe7i7XNQN6Y3WxajBwMrXsrAH821hCM6aadbQ0v9Rva24HNcIHmfKUDspzFekOzU9yGfpW0
fWulISNFKBsu0+/BoJRhSZ+oJMcibfGGrXXNCQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ufS+qjgKdn2oE3oh7EcYzivo13DkHjOXZdvg+7gUZzbjFQGb+M3QU6lNcH0LrOEXll22KbI2ohfG
TzYR0mnCNIzsPfjq3uw6taFIWJM74+oLYtSXEeuY6ANmuCGlqaVPg2smc7PFDAPdH082wsWirRmd
5thR9q4u83J5L0asBhDI9ZTgri+q5MwrlbJ05yQiFPUliJgl6amNWt26C09sTCAwIMPW69iBKeeW
4vt5DSJ6XyglFS9MDI6DvF+Cy8vysZSNzc8P7lm9H64JZqo1p7yTgGY0TjifISAPXC1fHwrwfQXY
BsZz6suWdJqjyzpfb60JVTQ+/k5D70Xj1MXLQA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TI2B3m1FrAeKaU6k30ykyHfDnWZXVLw3GYVFmPwE7PU79Tu2R5dzZ8wRPsdfoPSTye6ipaIAsPtr
CwCMHFOrInoC4tES+00nqn8BAlNtkgIns4JutCAsylfO0tbo1jdQM1s3ZfLRmzO8TErqp7qh34cJ
cDScSpPoqwYzQG0FgIs=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pRy8ixMxliZyP9cGiEmLhkLpE8BPUs0NUJLS9EUfKEgqPIYh3TC0iGkIkNMUl3FvP77e0IxaktFA
/jqS+a9b+rZb/lQQUSJMP1pPdZyeKNO5EYTlJkeq4M/QPt/jHeYrB9fa/fTRWFaLSO4suMctHSMB
vZbG6s1wo4stlPecixWiLDS8vMBqt9xY7MLA6d9rFSok/TUkwwve+vf4FZtQpUFEhypIh+/V1Yj2
bwgtk5lfZpX3tS8eSCYcpYqNluL129jpVqEYjJIDkcuxvvuRJPiKMpRwiViOhJULCVRU7pAOu9+4
kiLxod5VBhsHJGbgGwc1XTZvGawHjedADbu7Tg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 124208)
`protect data_block
stHg+psIGYDnI7a8rGIQBKkSU5p7JlD50ZwtmtZN2Tcy0ssA94sFhrxT15OED40MI35z59FelUmB
UsT2Bs6Doez77bUjpnmPUB3IdyQOQGCPcamR62XXl4aWg7ju6s8wYI44JJ25az7hWxAd45qV3ezp
T1V3+Zg3giHl1OL+mh9OBDrKCColKxx/0WY5tBgFCJIT7N4rQc5vDZcl/L7bINA47DHc3hZxAo3U
8GToZqKcJejKE6U9KUhM1HsHQmZ1y155Dpj9VfQxEMSM1Mas4PYEKhRUr0wPHAlnu/ialUsp8qpY
4Oa7m7Z72CCu5FuPLunhRjpRYGrmsfEiSeqSG5hbVMFO3CNn+WwBf0RXjcmxAhMUnt3OGTVo/Jcd
YyHqwo+91/TDAVmsKk7sM1RpdzpN69ZJuOjks9nsXCh25C4a6Z/EwvGdkTjCY7cCOVciYNwyNaWk
Ex/Y4OkFhfFt+jeuJ0u27xbln8LtCS87fWHG2t0BXLY2dDIfh5bzL7lWoN18kcDPmfaW1/3mzt+d
r16RU2untt6r2wMpdrbis1+0KxdYDjMEEn5ypXcMM+a7qW7WY5X4qduoFK8ru6dz4dJ0G31ebY9N
DjoJ/UATyzYArtXxRdm59p9gzD2C+sC6OsIvyQxyrU1A9q9WfF/hQ4+jtLfT39+3ht+K3+u7cXnp
7ne0/ch0MCd9H5A+mSo1ZEF4Cvvo2+tatzt//IpKGBhXTq309YGBoai5LOfIPLzdJ1WMH79DbZ1c
pJSyMnqHk+403B5lyKvyCoyMBBI6NO/DXamWcxmfiE5WpANjpTbNUKoerQBHyFcw75R4l7/eb2nZ
cqqPsWrKl76cexgmeGN9twqbtZujBHajPvmtVh57Lx/YJZhTWSRTyy9HcvVSlHxC3bAvNqQv7Kps
d3OdB+9rLqFirniXS3h08mOUbmqkqrmQIEoTCCHFyNzRKmoGdRAWh/OQeNRXNw8RJJXxUA+ayo6d
bjaLw/rTuoww2cqhSkCI6TSWs1UPhlXuzVydWarTXgKX2Wrsw831zPXSvnns6lAkll3P0avihzZe
bYg5hNqkLbmeLDcqnfagHJE8JwJXSKIoplQN/ByWsPY8zLhlzJOHwfUgb209C2Bs2gqEfNOGKmXD
OHlUTJyGG2M7xBDt85ANDnLETtiIdiRyH6GLGQL7nBsDq42vyfqSaF40TE5/gZ3RSqcB0hRf6DMe
f6ETqxIFLVqnQcXb8EkavUCqb5jcv+OdFJVGBlmUrK9LB4SG+yM8X2i4zDXXGWPOG33xwDRXCA1r
TWXAQqiz1BELBvH+GEYSciwyxo22V9Gva4UuWpihxn99lTbs0Ma2+p6fGeoU5x7KFnfjO/5G7eI2
PD6FcJRqN1plEC5oGTvfO/5R6S49BILB+ex8cLdnUWbgCoDvbNjy+xGTuc2K3P9NKfmQ1T6FRXN/
/8EwoUxVGutndF44faAe7PaaYBgQsiijI4JhDSxMEhyGNl1wINFYmRg41lL/56hryce2x3z1DoIM
wNRRxqdN8xv3YqXfDfNrIfFKrxHCwduKcQQlF6v8AfIJQxLU1xxbb0StM+q6XJp0ejPJm4LjOXE4
3uViAACi4fVSlzWqxq+ZTkojg6GdZBDZj3aAMCFHLtzzdIZaUfQ4RADKb9ljaJiNlmCXENOuO6Dz
IIDyE093I9CQVhorbJPpiGAfAPq/X95n6NO/E0ZG8EvzdVylzS68YKcTlgdEEo3+tJizZfa/wTKH
/d/kM3HheVZesepqFc7fwkcedtIT1f0w84Nz+mUZNZ4M7wR7+wAXnr/Ft+XdD0xmGkawW7z0aZ6y
ru1wlO/hb99CW5DtLaAOyEYSuoLKKuSL/i+9GZ0uVdvLsX3AR+wI/oZkCOc7JtQ6+fXRU3oWDusR
g8qWwSyDcupj1x4/nsWEcztdgCwBMKpTvpcq6NWMkTjWVau8SreeSLi1RkPPTYx27VOZ+Qt92rFx
469EKAoWf7Kw4eGQXjJdQWaHS9SWjs3ftffXKcYtKgQwFaI9Z4yroKec+q+59zBWaMZ+592pI7Vp
QP53VjRizUw2thKOjVyyTYj6ohA+8z/obVFDpVcpRUXFYIAfa6b9qp5NXCXdcyshpkno8OWU1Hdm
bCu1+HKcyljSuPHBTQl6CYr1s2C44hMZU9yg+ecFuP6WyaWW7xaBupY07AfWaPXlZWJpxMbKsAVJ
9X5DpNdqbSlzFTHc0k2XJDRphaLroPDw3ELLY7HI36OyPRSZDx15qnK0b4Y40J6Bk7Gmo3++3JCL
4oTmWLedI0z1ZBW4fvfMMadf7H9pb1uVU/uVpgvVqrwcWGNVhhos7HiOM0Y1Ytoe/wOPULKssNIa
KHYbNQljjLA7CCmPMFXFpPr7Xy6nmWn2DzrGWFx2t7QdR4NdubRxkjupc53QxTg/rzkghzEIZXMl
gwTzFe6xvvJYQzTcS+FPLey7qKLhl8JipjEfUDv5h1Rvov3+6Bph2K0XvoioydQLdhauctgeQaEU
qhdrw+fdEKsTBJXQM7PelNGB6t3XzN+BOk6FjyHFo0x0N+j2hTFvmgPIdGGC14YSIxgszNcUUyQ9
PU3sWZUG4G1GLnABv36BSwdsfC80X56uOLFxjCP+nxKspmI7fzrEmv5QFl5Zinp1WmxaGgaGvdFS
x7uL8ayYfHLy3zVlv/p5sEgQz7al3aY3rYLgr/DVpoiRJEUWpi7Wzmfew29xLYIXBNdewhgbUNDU
7pLfeu+HkSnwNqC0dGE1aAk5FR0S45nmQnB9vWkZfiJmWG1N1pGe0LIznxL+YzApjqgtB58XfyJO
tHkWMSzLEjcx9Ycn6VeAfxznIXSiPdQuuAcQdQZBZIaL45B5pfyT+GdTMy29Uu4Z3ptC71ak5j3l
7RuCqvQrGJbH2nWE+SVe0oVO1QZAFoX7yJGlV8IGku1GSApExW3RE6HyDlIbfaDbjaWD2cZy7g6T
1FfF8JBjew0zYO87K9PwI5d3mkHn7CL2miCgscXhgFjyKIqZsgl1iJLLFgDRbwV9Vpv2SJIWZ3uu
7RW2WsaizXUewSMmKdljqJf7FkePwbFwP3YWArIVLTRYct6bibuIYYHYm4w+cteJNhd/SIKNFl0+
BVL9mBTbtq8VXfAJKPsR87z3eAUktPS+E6Nsq6OFSGYmUUZbG3AqDd8+AmzGqodt/SrVym1ncucz
LGKGI5Y6aCSVwoZw1I9SvlkC32bqx7I8HGez/uRoJdxGsUGQrlPDDb0pqCQ8e/b1bJ4eXUE3sPVb
cFT7FaIEGDt2SS2+IFaS9Z8dnhCirKfVO/nYoiVPgcqo+rOafkFVCGPl01TrEzeS+qFxZGpYmjNH
2SOXoSiltOIITHLnjdgJaLUKQVt5u75MtnFZDYQti7Jiw5EaLGrAKWDYmE47D7kOi7TiePoAzsKH
necMVHUs/JzoQ/TsUPwzlQJ1+AP6lfurXE+201rnN24onqI7sgJJqYcZU+Tr7vuS73b2f71+69PH
h07onZFm416M8N/ScftPc7C1peU0uFjeY7NyYgG1wXZePG/cvWns7JZjuiKM2auL1huIQpfOavff
eL8jXT9wFx1aATtMXBsmncWTWG5KQaDsLfFqHberOCqAPskBP+5Z9iDc0hCOswQ4fFFni+Z1rGBq
wF0q9xrifQNh07u2zqqG4Gj43zJc2Ynpc412ET6xcZ03VAz8Qr1xHOBKx9HmpMhbOnBviMuvS8zu
IvWqIUAjWkT0HGWgGW7BxE9aa+576lFtCzG/DVPkNqmRHhfHihe2KQrzFR15i8CIF5o+KaP4N0Bw
eKbMOjHD8TEe00k7/ZJMJVr5irntSmSMrG5+Sz25O34keNoHoaJUlfr88MZBeM7h31gUjdG2iC8/
/TGTbyxiwGxiug/FCj8PJ+DKpQUmhdJfKqZRr2z8y7USof/Kp6vB0IfyLjSQJcPy3K4rlKqo8vTU
SeSVvra3Rr5zGXGrCjCym1gESnYuXyzP+v4kfR+WBOarRjAe0oFdsJU/rYUYZ6/H1Kn5ICdwwJIk
L5tb9hVPiH586mrLdbbOBy1Lmqna+LoNQh6v51IRNUqkYncvZicMTJpFofldbNpswjv7Qcwrs3pq
TbDdSi2AJWd6MSnFjU2e1annnpPLqy/t1ufgnRydX/6dQuzm33U6/fYHcfaF+aA7+T494zz85915
kG1ZFGXtfnHHRvOIp+plJofkdP+OAlIJ2pc5YTfMYvrYulMKTKprqRhM2MUYtCxp8aItKLI27aOJ
n2EZSXcleH15wx60G3nH3J3gM4/QWsw7mp0EPsbmO41KGHzfgNNjkQTrc/pFHehlTQu3f4KKeUo1
awPIqH7+AaYrgUEdiRcTXxbcYi53jL41+8mRAA8eiv7nP3mrmg1Cn24Upy/ebamIHoUReuXVgSze
ts/tp//vheSmWoRQ0ffvKi1DyT5NYcEvQr2zpPH4AkN1n76jw5fQpgv15EFjwKFgaNiIxX3dhMWE
2/ZAPNv+9kQS870LmQqKV46klJddX1fOx5laJLo2X2F5xXQYCHlH0GXUXuykkHcbT0+SqTF1PJ3k
Ka0as65pjxy+IV0PkGe8Ws2vGZjOxKrHIgkMhj7pO9jvg3ZuyppVp4ws6Jm/FL8Mo17hbfPpm00u
V6cGxPHVtCLjxpgQrJz8YGlTl3BEVryb3avGaOZlVzt2zHV8GPhfUcCtXOc5N7x8zn4dw0Vnehpr
Hfvb8BhVMDJ3vOxBUiG6iy9UeMMl+W8YrzKrHnUE4EG8MXf64FwJ+7etLmSMKeEuka57kuMF/cSZ
GVfY2n0PUjv0qvb7JqhsYTpJlp9/GclzWWiYl1lcXcnM21l2Z3kK787euYXhSJIJGm2cQnkO/X8g
1j0M1o58sNuVLICmKW3MMONskW2MW7u5/SRYmqoZii7OD1/UjWGZ5sC+KHIMcaGAL2O8MtUMksW+
ssXfCNW0BQ8J9rGp7GHAnGVgN0PTnA9VUmuzgRuegTWsxOqCOtdFlEV8BCYNZQWRQevanw+ZWS8r
3hHK0VCgY7i3nIcmM78b+m2PF9fOAQtRcdeWtxwkwe2pONjHi4sYTbYAGXRfzfxJc1lnlyQHiH7C
xoPdbJrWovCTFweT9T+e2+v1xrzvm8a+oUVyzqVllfWq2OsMrIArG+10qaBQetYJvSCtwmbY7d17
B52BThr1O2gwCG68Ahyutv4DpsBg9blq2XlxTNIYOVbosE4CDtNo1OA+ql+gEBGALtI4NCDAwQvw
TFUvOvZuLnjIpkhYeu2JDg2qBcG9KR2j3FCUw9dV+zT707TfwkIRBaGvG0L7elCHKM9CHhVnXy1o
fgGG3Rr2SoUANZt+F2O/Lk+M0HNfqK1I0P7DDwXEa7W7BltpLB9BPzY9FfwX010DFipB7951N+R8
GRhJWL8uXb3kVpynKTHntsNcycjc5dmSbEbVv7PT7lXZwsXUD+hKUV82uqGncvxT0hBPlkO1NHIf
8ArgGQwfHWVVrb5J8YS0B5wZuH5skvVeAd6RkmHycSGh6cxyNnXugzSa+SL5kAFllZxBepyF39Xu
IUsvi8Q3LGwJHcL3d0DJs7U3rfXYSbOf0KH6gocvMlpSrOAq/7qHLhgv09muPdL26WAE/8+JSTEb
sUdfpUgFWuyWQS6hpV/6cwLOFZpsqd89KJpL9DovObQ2zA+P61smyqSrTr7FM9YdOC8VWxi0dS8M
t5aw4p9TtMT9diAU/n7H9csHcwnX968/4NLWpvLMNuOZS6mmNy5tGJX/aIuS4nCyoUTQ9ulvCiEO
ONwre2eblQp08daNypC/cnqT+eq72ut4XKYRJ5Fn+VIXbTS3FPlUnhlhF4MiUAXng9y3oq4AFFlU
BUY+CByZvvfpHMWj/jkXRoEZN6IW2PkHrOjDT30cF9y98VNWbcoDsuZHLDS2esyWm6R+IorIvVC1
BCEbmZNDjRlpwa8agr4oaiO5cKJJ0fj0Ep1Bgryj0CLBlD5WdNtmuFT4cQRbYEpU51oxFPxB8lKP
gudF+A43MYGdq88+6C0eq8joByzxOvv4Fcx9kxKIaWuNcke7rT1CUmqldrLfH+sz0sYlaCCE/dsU
LDJvRE73pYMj6Sp5kk8swSQv2/GcScnqk/Jkfv9ssbf4dTEWi46WdqIZx0onpGqDzurw/cU4jd8W
bL5ZJdmg+nddVY2jkvSZRaldNdKWM7hMRfLv6wOL6sflrzg0VMzt2TtyQiMVwB1cyddbRIJH5Shk
ImIZZXv+8nNcfZjwKwGclZAHKcTWHBbPeLHmNn2tWtkuvk5yoqHEz/Sj3D7CAtfLKca4DJhTm1Dm
xmdExsAl02zN68+ZgEhJaWjTOQQS6SvZIiE1EgaXvvChNPQ5cj6uVNlV1ItrkCp9dlSjDlKVVe8d
8EysDZSJOwXaDNEylYyQmgUNYtYeeD7kQTgme04uSI+XKWN1+Oj2JbzDpI55fXv5/nSb0+jtGmAM
AxcdN4GgkZMn2SFFiDiZrD6zZEbroTl3HcfBCHGEKK2q8XS6ZPank/jWDJXH4nRi6NoumJZAU6M7
lNtdKOr1hC38K1YYLVrkV/pmgeH4HsnpMEojOX9sat+Edx/PIA3mnRcRc5wS9ERl0aGiJqvoFMjf
JChXUC/g42a8AKPUL33/eA8roKA1R+zvITVyCW/2+57khpyX/V66p8XyBe9DUE/bhIqzbyXfzizm
x8RnxliS2Kk1a0KuQzqkjix6CHnnz67XkCsGgiNuQKxO5NqxTIqs1OlTZtc78MeZ+elImiZhxJJj
zvB/uRrMHL9GuWkyUcETiL2+HwzKQF88991OoG7wec1NbfpnozKknKegBe9cxRw6Kmktjdc8y4ZI
nm+z5ranuq4UJW5Avnti+JHZEq7sZps75vQIjpG19T7LMix3pk/CyGk+yOhq/pdLkrlkNGoJAoj3
jgnG99CCLibYaEAblbqb2Db2knn43ByQcpDKA9IFKtekIjtQ9B6ujDqosCl7lGwEMZI8QizZqb6w
65Y53qfs0uh/IrEKN9MWXti/tagCv5UgPUAcXpXC/3wjmsvv1pkW+t7qi5kPC9v/sOYGUIOWkD2Z
2QzgPzoETV6ILznwE0LCPsVDLkwDgL+042lzoUzFx61NmDbrrABh5MMygJcKBgrNIgNFB/o05d9C
7uITDN/p7FrcoPwi3i8BGBoNfLhlWaghr7uLag8zaP1xbaTkB+buOrLsOedMBz/zNldYyqJHXjlY
JbXGuo/wCN4szDkEtr6/uSGvysu9Te4z0EggQ0A00lyZb4snY+/pXUX0C92MzlR6iBGtISFH6rV+
JbcbgoNa+A29qsfR4daEpZ8XfjKXub3n3d+Db+V7MsVnCYqI+oQkdXEMRxT1yC8ZSPoncosYdPDR
8oXSpnT7uXRil6S6ciXNpfrDPNwWWxL46FwRj8YTaMIkmmRT15eW6+mungnNzKTKKcCr6ehSnA8E
XcxdS+iUBo6AG4qE6yxtpU20vT4AXRHczjHIzLoWtIUGOjFaUdROgso3brEKNHrMNqhjLcrWzrvK
Pj+CBLek3Y/YICudnes5HSL9zU6DclypVcl1G/Z3vCBmGntK2OWC6/QhCBiKsNABSM7pU7M1ZcGd
va0ug/zMF9GpUndyiUBi2nzdijdsyPyu3emy89gaVn+oGJnl6w/yHZZ3bGfZsVy287Uchq7AeMVG
X4MbK7o7CEnKphTnJ5XwQdxuims5qRSNrjhJOJdMlrZgfVcRK+sCgmUKxu01DUO7jr/3+nyDFIx/
hl+8AhCjahCoYOHOYu5kH9Pta9GBXY5xqjwV22+Xub9fgl4idu5CEDymVudECRR8yAmaDHRcCMIu
ipD5Bmv2uKMvnXgzkP3M7K6jK1mBW92kACcwR6PTAX5qy6Uu4gmQL9mvQyMToWj/gmXodXmU73/7
Q6JbmvKV8jcOzOB4E4XyIU9vVPAqrZcH5+dC5zPHiCmEKD0dGC6XLxMwDjPRgCZIXy+Leb3jTYgD
1Gk/8oN2pdtD1XnFRsr3GdFFLpVC0qQ/JHmT8/tmYFJsld2uRdGW8AeB7UovO3bPealHYeo5ZGyO
SSnPYzB9yb4Xz8XU3RNNd1L58IXycMg80Hmfy+AgpmCtN6P+S9X/OhN3/d5gimpiphEdlA0Ed6DB
qepI8fMFDDW3SgjjgwRUcXKQsMnBSWOJhQS1ctU/1TAiwpVhIsz5qFEpIDaH4wQ/gJR6hI0tUWyL
65Ok87ULvp/9sg0IwTyc/hQycbg1tVorPk2u+lmqDscpqurmhuhEHoqiz0jt0iheHf68rHvToOSC
l4C5toVk0MQQvIUaU7IpWA4L3sUPlUjohQ6n3eFTXAMM7XTNUiGqlyIa68UWyPW6x06MoinJaNhi
816+D8UlmWuDTNSy++BMznmrbIXKMW2DNlMiRhkqYJcDJnN3VBztVv3DAItGacZv/zvRKqPV//Bx
PTDN2Wyjc22DSO7nFjwkTCcadWA8M1PGhDuzns83iLDbL1tcFuVeoApfffRVhUjqLhmpZJ8tuSGw
lTO45iKQqWQUYVCJfSzMyf8r38HLwR30zWhxk6FqVLURuqFtPDYyc07CWJyw1JYSq7cogzNba0hU
G5tYq9OlHQUSTlOnW+H0KTO4CADuAzGHzbcmp5+tDp+YFObylpKI+FEEe3g7E3/rEhVeHSnmHNsE
je+elLD0dPpl4Ir0q/nDPlJr4EJ1qR7yTrQcUhThzNv6vmJ23zt53hoA4iol84vAySBJDC4tpLtE
ZGztFaAPap68XCke6WX5yaL6zXwMnYhe+KknyCmWxELIF5PePfISm49mEk93DaWnncH6NjHPo093
td0azV9lI3ioYK5yvSnH4GsOro9qjIfV+IqUQxBbwp8XS2y0WATifKqOiRJ+HbVNxkFJIXzhkpgy
EybmFApi/mwGoh61UxuPoCSyqm9RHt4qaXtOtysWKmLHmhwD5SKtV5zxdhq8z8M0nOLmris8f3wh
ZrqMXsvYt/zC8lHC/uJq4tNYH0oxU8cnPUeqaGyKfC5vBFBaHKEzcgLvm/2uj8gTgvgGqWpHOwcP
KZk6oT2CukC2f9O6jYW7MtL+q6Fu/q7DY/ol2CXI6hhRxKXNyYtF6fA12x2E3fYIvBX47QhgO2so
1Lecv9pb2oKPYHXvP8DglCTewPSPpPcHrYoxZLAj8SYdeeegqwfLUGlWNHqX+hwR/F9nEsBo7XhF
2eyeH+5uC59r/KFRMpEch7NUDveo20UaK3nROfXF9JcpOFlQ8RmFEu/8aqibdOgIU3ef5Ujn4Kpi
Y0DS0Jo+ncrW6bOE4WDPbFBfpbXuEZdptSP5m2l0hGzpPpU/UIwUrbSuCxTP1pRsBfjGR0XENSRd
8rUjY8WIP3TZjsrZjASmNHf0KRekmqBSJlF1rM3wCTndIST/Wbe+/qqUK1B3+cduEeJ1Wg5MRxIc
VCe6Xli/Ne+74czYqUm1MMD3lqhn6vDluPd7/CbrEVt3BbbxZFOOTnyS/l7A8nY3N6JqYlZQrj7r
EBWLosEsuDr9ms6qp3pUbWX9uJAtCkC8OQ4F4k4j8aOFZUdvPc/pQXDa/AXKLmyxfUDVqO6v4/Q/
ZMQJvAC4AVlu48VpH94yJ6xTa9jAoMQdeNixwoHxPoCEdsMQo+YjArgyCWwNKjnR4tSo/xXLvue3
7BvTVz0qW8+4w71/GnqCdn0YmM9hTevNiNfTsJ5v8ek1YG/ys+rO+3avYZ2qewFfefhtURenpRgF
Y5bFM86lRgtUkAkBykx1Q5zUUw2HtCFJMnbH6qOiRkHUa4PVn1Bn7Szb+tHaOoWArK+sBWGwvq9Y
ABxEe2moLtOBPHVj2NqlA2WWTcgunfBAMoegN5KUCSoB6UrBrVS1uh0TJakGBq89dag5inTOkNum
dXsDU1ZEWIIMLveKn43LK0U3DFBCcnNCQRvBlpreyP0q7tkCLAP4n+xqw6m2EmLNHYrgJMIQoNgw
oPP2Lzvk6nsmXgFzOQGbIcyMTuFHpvqv4YvXqIqdSAWT+O1pjXbyFbNB6z53Bxcaif5DFidjma4L
DdJc1k0vzY7iE+dVifokuaXXN1tcS+GsvqfLTbi367bVXM8V3G7eDRrylxI4VPZhoc+B60oPt82f
vEmhLZtJ9pmIW6wEEE6NoEF/9smZwor6SpZBgG57FJ3k0XA2pyhZ0rfPp5fAkVdKRiNmBK0/UHNH
mIF7LNIvduLlxlRTpIKRSR+XCYlXKrhVpBy1tP0VNtxrbF9X0P7AoYtqufmzxlisW0K1rICFUQhJ
fmfTaInQZFrWiajmVOoMdp7w3y23YcKAgbITLLcX+mLKuT+rZH81geqwxx9fgdiY/NXimjJVMLw0
RpkwPhJA8AaNZLXZEt6fcSWnCRw22PwaS/JjVcethLb/y/PdvS8ey3FNnN7dRvQ6iDmiIe2e6rFu
Or+H72w6JdjoT9UsXu4PMCtCKzBl5WOR3N1ZEccecqNVrh/bCt/hMRM2hhrz9T/vXxnX7Wm54faZ
+tdo+1RGmBA0k7UxCRGfgk/ssuDJdal0P6cbtjCuM4NpMFa3cqVOlYcoDB/mn/s1zqmiDdM0/Wgw
yKLfM6splH7mPluonROSXzXPEojMHJBixmzfAj0q+Rno5B1hqt6ZNFtDkA7sSfRWRjJ5wQypCUt1
9eE+h1zX/m/UhzaHASXj1LcM1sVYsmoMDJ4C8xjh36W64mlJ/qqdcoEcbYE7C7z12evEP6wQdCOX
kwO5K5uhXYvqGI3bIOmg8VoRgiV3VSgdP6wIDjDRZUUpj2jI6UzIjzdbVd4HqV3yoIlH966AqgYt
VQOeUotePu3+YnAh9wZDb+1gRyGQyE8W89Uy98OMflGmcQytrkC3c1Nj1nfgn1B3Xdx5lAcUsjCs
uIcpnYvklmdJktWmSKSnjyJKpeTiVpMjjJLCP9kk4G/yvtN4y/B2C4SqwnMN7ESvQHMk2xGFVzw8
k3tpYCxiQDakiqoos17ukIeec6qPyVinbn2VdDf4QeUUskfzC1n9NEp3vOZgFEh9rRCq2TES82h1
Xk9M7dWrbCaoUwUE8h4GjqX9Pge8mBmVEisbIeemajPk3j/J+PZ/h7ad7aAIfCxfl2SJUi+OkiSD
DcVCJRsVxdJ+TShkoI49neOsGS9jbqaxmrYvnc2pQwnJGw91mLRZPpWA6jC+oFGIrFwK8DO3YUN0
0aHDvLYeRinqBkXPfBcm02mMWhSMuZJAD4RSBBJloPukqjus41Ky/9wkqXSOWddQ3tI7PXM8t23V
NXm0C78s1zK6X/m5k9rit8SbcYjhApD0ycuwsdsYYRz5v9S4KvzpB24VlxOlwCKy3xF6u6aowLm0
92IOmN+ew4i29jZA4t3uKQEekZvUHGXRXrJl83PA+KMGoGurDz1vA0zq+wddRdtHBy8RR3do7Z3n
uCnRWUymrqH5KAuaAcVYXLqDKN8HazpxoCd8dpJ8LfTtL/naLw8xd53gZjjNEPDqTXD/6bOYU1Gs
b4VHai21JgxgAIuLnoHo4K5EnJ5jNRegV6Zw7kacwhKa65+3JpK9UVo5CfJzza2QpXxcosq5DGy5
gjW9fXZlmqijaD0DizY+nk54AlUKXMax99GMVI33xOJVyLleuxNNakPZBWUQBSWP1U0isYztn04b
VOdXvclHp6KjUTqFORcX7tlXEPuT21EWdHOaVGpUfx2h+CjhfGwtKJmRoUWQ0CmHAxhiI+byUcGl
SIONHzKNZUhxHDexxYA4xJBKIcIs/Pt2GLOITolklsCMuMjJSpvBKxz/Bf21wB+cTFcTytViUja6
rWHoMNpt9+uj6I1MTNfCS7m6ns28Sikbw42Qj18VcKj3XPAG/m+x9yuPjw+bqxTXKxoBHL3ZA0yk
gzhDt1ewj1EagdqCD7VhMXzaItACjijD1fyXqdVCuHdhbcESOxP57ueFwhHjv5qRgC7W91e2AvpM
H/yySBXPtacDSu9VOSMLOFKwfPuGMAVd/M5I7ouHNB8pCupyxRKRDzmXWiUnKVN1h+pC+XbQYjZx
y28Gf3pT2l+nEeJhwU7/CJsH3qCZPOvwt9RWgwkr48x9gssa46B/Y5Dv03ViM1L0zghCG7SEqK9n
aEN1kzaxZ+/TIZ0QX3LuIzaxqEhsgBpiluovNC2m/Ec/gxqENRP/pSQnbigOeJpY3drZrVA3MXbK
e6wYCEo1ZKbQOzIH62CsTN/WoEAey0avewhgQ7TjHfdfo/dwujsr/pB5+suIoojFgx1HQiEKgttj
4gcNNpAQXa3BXt3p0nz2iL3R6h2PFQOAygbMzcu/EDJPH7IJSlhsHY2zMwzUIqCOXHtPJbn3NTam
1iz+RwFElA2vOTARmweyH5kHukNw+amNazdlSdTlx15iLsByYG/hBBYpzIoRHSuBXUscQg2jHTP+
IXkKvtA2YaKkAD6Xgn/60MUYTdFIKDfu/dK7nwFQPytVbUf8EnV2xNgHiM+C7s2zCnw3+tAWH65Z
qH1uLlG+iroLnvLCwxkiohPCYdqIY3B3x8psgqttYbTxtfO/JY1Oc5+zjAivuRGCRbqnx9ZyJY7a
7u+uxWFzKqXS5+TMPDQmYH9DlSwn625AEztidxOg8OFv2hc4LmJIMkPRS0EMFSruMVe9tkalFddG
z/ZHw4SnD3/8GFK8SlU1Wl/tjQT1ulNmu2j60vXWhwJ945L/H96EjiFjeIynrluOOqUTRkNiXIZA
cgGwQ/R03Yv247+zOUVLoqOYoJjOLNMkN+eRkxaqCzLjI3MmJLXAUnScR/D43/RKiPWne3WX/cVH
iNoBblLm+RbiTJmDFHcBSXeeHrwoLJMd9l68zyTOcTNUuco8ax/gsF3uu6cCKNqUgESyOC+Za+pt
lY8T0xGybG5YQBAMFY3vPKPzY+gK9S43rMCSGQ0xb3+Eh7AbJOocouAlzVq/4qea0HO2TN7RL6/q
RAzKwWBpPmuZe2+VwlFZvO+wq+gaW0VOMUpCiAClClabf62LhLOLhgbvDI/bCl3vuo6QUmF25WiM
04nOCtX62qDgZ4inHqXMuPHlLCIDfexIix6om6e/DEqtNC8j0+WBPXxXN08oFhITPw4q2m3NxNqd
M8QhcJF6TfZqR8aioVpIXq6s5HxGlXpKPZgbV4d7iyn3YSFjSN6jPM7QVv9bbg498XHQnYLskcd9
hTV8d5W1wv8KgUiIaTRGRKJaEM/0uika9UYO1GiNT2lKdF4/Ia1BGea9iMIZRMbHcwPBNMpEs6XA
ShiAA8e3JoqMHgpGZ8kDDMrdvw7NLyfY7rz412K7YVvu7ZJek8S7sr3DamTzzDi5F2T7Ol3m1KYJ
lgL9q/zcCA4VMnnRaiSwrYj4S3nNgZT6gKE4KS4SYTzad3RP6+3kBTXLw1xcenlbcdTNWuoDza4n
nZPMjkhEMln4t/PvVGonc/ve/O0rUMTKgzw907SU1nAXW/g88O35u5kePDKI4xrlP7M7+uBENCxr
Z+B/EPCnFptyhQWwi0Ny1NiVN+UqQ9s9Sf4GfYYKBm4IqOSjZthFjFapo9LevXp/j2RRoKqJ8o+B
YXSuNHKyZyc5369N/QZSYd7OLgXz4tUEbvNXi1wSeFfwGIDWeOKYhaXCoim1w9HSzjCnNMPGBFtE
xAUEcQZK+FWP+Y8o1jYM6+sqiVxWomRziDb1TJVicPmRY4pdi/TYDfimZM+9JfZKlCsMRwZL0BXe
ry6/JhkWMN3ntycKBTZdyxOSsphml9GnPH3JEiK5SfVPe14Y1L58GIVnGjlYYW+86NR5xhwpgbVK
cNKqHjDADhLxg2P00YoBfju1fEOcW6mH0ueo5+qfvCB3bXatwUuwlUJ8W4w+XiMY3f9A6HojALK9
1YThONUafcSDMeu9Bh7gDUhSaWeYhZp792r/giYsFFsrUgnD4OnUCysAcRCc+0zjz63ETva8MmxZ
J+yzHg+WO92Wyu7EZFfafynmGZ2gEhpEtvW46a7KuXwRD+kuhlzOyap55OFBYLCAN+RmaPCdj3x1
9Uz8xt6g3Hznpu6yPfbvLNs3NJ49SwjsO2RWFW7AW4GN7vdt+mkFhNsltEhCdjmMH1glPSHvcjcp
aJSHZegoUnwjPgvdPUTwxzl9b/1JuQ7FjRLPhzGK7/J9+9Nj8+FM1PnogdJE+TAg0/vjo8MVMjn2
9zDEDTTx/r5qRCV1UyJCthHUFFbtRu6gngwZOGFpAiR8vW/ePwX/RYKRozXO/96Tt35BvH6M/P4I
H3D71NIOvyEInEv9WQ5HvW9K4IQAmB+Wbqok1QsKPswMm0GQM351PH49S7F1IxJ1OGs9mOCub3fI
HJTRiCT9pcozo0x96uYXMjYkHMTWpIz7rUptIGW49Wk0zZjulxoZFE+t1DpZxEKB3BH6/C2v2/4l
rJ7mjMACqODYeIZG+LybUsMHIie5dSRET4b7nE7OBD9qcyHeGP/d4NPabEGP2LjI/HRzMXfBPZ7M
llQ56cx3IaaeJF2urpxTQ5ySM55QbiyNfdlNEGsFiLY3Np36Z+tFq6aDaVZHUMNPA+Ydy+7XbPyK
dYcKvp0+TZWl7L7hmS/jGdmUMF0I6+pGgazfsxisoHnnFicDr7xg64P48+WPJywy9LZkxQVYBHGB
gZRp+Yw9tLaK/702qDc8I2JJTLmTTne8aNCtY8V/6VsxokljEQ49ZldV9CgXy2mTHSsFT8A67HFD
7ju2gaReA2vKzp2M2gEuKZSifQij5YAIwNg0FQ/fRK/blQ3lHdrIMVt8qPeYJ6iU0O3eLGGY8dBe
uHZW4+4XwqNQPwHA5MzSYIJOgnUEhCkhhjWv6do9yphaE9/muf6Ynw95pPMnQTpTjR0l6XzrgVZM
VYBAP1Ecz4O3zgzYYJHWxe4lwtQ5nwYpYczVyAkJJYkotjK7XytdVcCofVxilOlNcaiq3tzLk6D5
3NtxF9f4A05p8E3XT0pENSKpqPVtl54YCo36rylUUnhTN/Do1dIck6J+K3AXOpuTbOR/8Dq7Kd7I
GhipvxJJI5gYaA2z6d6r3roUKfPLRA9TiOZUxIzYUDEFvZLIl/XC6d4H3rtl2o0U/fzkR+slAgQd
3OzS/zMi+1bEX/CsEWyBLDzWwSH0M+a0tPPPLnPHfU0jXuy77rXJFOzfAyvE9O/LOq92P2g3zKfY
YobXKOq74ps0h0z5PT1mVFReLe+xq0I+Mk98wkG3WripD3OmsrAI7NgjKm1xCRVRfN3jQy58A//D
5zEekgnQRif83ACcsf5on34Dx8+6mQMyvxU57VPhQu9kLbFvIZgoQo74LXzp82EP6K8buC24SgrL
+RiESO1b0gha/p2LVsYl8y15Ng4HQzlGSL2m0P0SB581b9aXvuDqZRlSqe+8DuEhlLp8Ae4zx76W
cuFfBtpAYdG4o6EbzD9TTbVDYnoTQYuu08D6vmPwV11pYohSpKIQh49GipawSLcgpfRmWX8bMFx6
bSaiFU3Ebf49yMmKmsvZa4xH60WZTfgKe9h3hqk/y+CeCek6x793MT1v42ri3l4jiVYHK5qZbxj4
4N93a3u1cdzj8QxUBnKeh4NsS6x8mLS+yW3hhkvC1/eqc1+aDrI09JwnLVKESvQWcSoGrtd0eVUt
T3fXdVmGKGNXDijVTDlqliI7MBJdP/8KfJ+ZyOf9p1IBLgOay7lgrYvOjr/r3NNhL7DMn28Xy6Th
3hlaNodW2a+V1WIfKKDATM0A+a0LElzVUA6pseod3mqjxC9sMyNYWD0bDMIM5vLZ5yIcT6hnQFBW
3judVrMdh6yDIfc0+I2EZvnJCYPsGPFuqm/itXAd+1Pw7vLtRnSxtn3vygqhB5QxJUC8T0OkLQTt
afzo2hZMGufmje9DDmaFJJyes348vFguSeSNBeoKDB4vaig020+N5/t2G+VpfSOO/ECdCpsC8PLZ
NpOUrwglaAjrbxfqTdktt1M1a/BtUhjMhBKmhEWbEOCqwf0LvIXoVbbUwObede3gmifgLqdy7bE4
aTzI5haVlzZjLS22m4xSTrk7WuvqSUK2P9gErK3o7YEslWd/YgkcqTLPWzz7M5sSWJPYG9XtcZOK
nfG+wTCoU1UfH6ZqTtCx2whTHJMiGRtvVEkZD3r4LkhB7rrfM5STOfX/QuBHVzb7qfPy0ZDMwD1e
3vIB1v/kwpuXTXLqggK/pfvzQT1WEQJ72g3RxFoc7EEwET8E4r6O0bgoE89jV+O44kYupmvc2AqI
J1FiNEDfdmHeQekzFtEZTo+q6HbMNSzv3/Aym9oqNX+o1OdFPxzZEZa67rcdWje5TxgcI3ILCgp1
o/Od3vPodmruucxw3XxT40kPJSG01MW5uKKJIWasXaAMtRRrfFeNKE2lqkZVE3WdAh58mdW4rrxK
iF+/AfIs7geDBgK9tgD8jYI8TY7odiiGgqak7W+Y0M62VI5gwtm72ZqwER5UNHcib9CoL9mJdiTo
mVKDC00u9T1yRKU+I0aCqTpC41pmy1/GLjvQHX6vw6BiD/Wcq2/Z44HOah0R5gDH3uAbY033P4M5
s/nvrmWiot/B2Lirkbot5z7jGVT3wfZd+aXdhm4l2IJU8wzXM4+QFKxm2SNXEjf8w8Ly7igi+s2n
zsr/bmaB/7qnJUuMEQLZlBBXaH/qxc8du9k0pWbFPbDD93HBb1T/0XuK1jWo6nyF0L+jXtOtASdx
hDPMGrDSU1cHWwpx4nMMTmCe4fwOurkdR/6QSQvbTEjms4eG+z3YLSB1pM4WZwvBYyynapEx/LTM
VusU49mslgAZxr4FZS9TFkzvm2tn4iyskfTLhSCJyrxnhp9AN9m0SfFv2bpeOkBHnU8rnE+TIlk0
F5aoIwt7owTxvnfrSnHazJ7Ko7Gk5eml3z83TKH0GnK4ExPc7UNYBdbzJDAEVyg+2hVLOOi76Gxt
1Bya7PtGIKU/kaIx796bTsq+O1nWeH6VKhyvuKHzw9w0q1umc9xF78zEGBhIjBT1sjcdB++Uo/fj
Io76+HRLwSYqxdK3reLC+wHGOInR/D0hXx+A5J1iIKOyvlKHMcwTMJCGNGfJWNdu9y/CkoMo5i9P
Pg4r8F1/HJmV8LNtJVVQfMk+J2o+QWFG8iEW/mEgC4C9b0jCaTx0s+ExOjfyibkJGsG9V0TSE7T+
Cc1kPwamyyqqS6Qq6/t8pmDEKfPYfWfSCdxMBZnuRqTZ0IJu4ZcbTQpF4YWDZJu8NL1hAcrEpK88
lRmjn9v4pMgOJDzKGkaEne/tkZOMk8qywOLZrpHuIj0AvRzdG5w1lggdG/VjrkpOMiSIkI9ZnmlG
xwPDr+//Kbpzlb1ixTXd8ClNiOGKZwGyIGwHUTcwb+WcMvkkVYYx+EuelNC5NGc9WLeaNOG9xydj
8Z5xiKjoTnZN8UW8OdpTku0XwRJ0xuLhFkZS6SHWOKtho79OwuUs6dVrb9X97bv+SQZE8nP823Rk
MNPm1TSJS01OYTxFl4EdrDVWWzR6vkUSQRc6s31pUGlTK1cI7qFoTxYpM8eP7lNdoYL43/RdNO3W
6qPCvPnXR9w+FHmVSnQZMTd1FYPWXygpoVGRrYXVsYxf9bGFGhFq5UIWBDa5VwPuYvxaf5go7+YA
XnWJQkDcyKCnGfY3UhobbunNjXECbPksIktWJveOw9wSWM0mU4xBkCb1RfKDlmAJwVtey39KfutF
1rFhbeZQg2VWWt3+76QryilOdc8/lNbe+x3DU916LxTS3KH6lGyLAM9XieBg0NCYlTijy4PZu1Xs
UJFDOzB/VGNbZYf9NWORrs8gi+Ksm/QE9S429pGgIVQSMpudv+19VuHSUlzwPvwRfiLpU2i+cDA2
51imIpG6T+o6c7hBfF6/npZ32d6rQnyjguiHpXs3RFVo7aQI/ZXAYugQRRv7Z71ntzwNj0sQu9wp
nXcgP/rrZfAs1b6p3MgViRqRPMdZ8teUIE4ZDfb4fVzC3SZr1RgGV1kvajvlBGOMpi3VGnErt6Or
IIPogZWLAFXeLIzAiiGnepXrokxamaSHXpWk/5Q2AX+rquJQMW+s2By3Ve0d0KnE0CuCgGyS51ef
KCRK7a4hyALg4i0266Fyd3sz5R/w0fitlSKxBbJTKbV8dNw5z56Jf7wZpW3RADzxLDgCOzTO3sea
t+nI3omgk1t+65w9Yog8Q7lQMTVxQclhWh1jB3Yt+4gG3XXorkf2s4fpMcrZxZ0x2ndGBSkmCNGe
9TQK+B6KEBJfco6wgYcCPjHTmuXOEGYwYVnbMDJ7zDHqDGXHErVOW1pzbcN1hhutO7jhLvsybfgW
icM0DmkY5l93Sg7pzbm1XwPcDA9H2ubOGW0HDTFPNH+K1nreHRqJaGh+DQBN+XnBg9Tr3eDx6D3T
pwydvGBCwkSEfVRZt/TEqu8LPWCedkzIPk5oDmASIIO6Z+opW1GsVwg9COpasjvDNQmdaHa0Yr31
8i8bEDiALJEWebgT9j0QF+tTU33f1XZv4C+JsjINg1eP/yg4l9qeRPK49+5fRTW5Seg/b9nZklPc
fLMrp4mQs9gmKjhxjr7gr1FWtbHnOcnsOd5gY3wPBCLa8rcdMSZxeeHOKRJHKXRZLuSKNFGVvTid
+b3e2KBO080J/pKVXKZ4LsNjdR0XRDX4zd1CjwyAJ7PdXWrUnSICz3U9cyGmA9RhVwWwE1Sq49Ts
LDVeforixhRx5vtcz9dJ6TkOFe76cQT/PMEYjebD3fTKIGkyUudJ32XNVmG0M6HkCWjDGphrYTRT
JGAwUmLiE1f/pQhCSrK4XUY+SJ4ovnbkgpsgaE7xK5AeMu/BNlvzcTUf/EPly2eOGKAcw8JEiTCB
UxgufAiw8hYMFvGUXDQfmrIsMe+Y9+LuolnUR82IxAQYr91elrAGAE+xm12vPvnBZxCrkAK+XVi8
JwJur7s02CfZiDT0F3xaTGCNDJj2PdgaLRHQd+PVCMTh+qlTvPiJ9pEG88HtWQd4TWnflzcSE2tc
tWgtF83XFgxf01VMPM0m3Lm92F3U/NdKJKh4jXOpEJ+TLmAbo3nEI2y/XC1uDLItdWmipsdoiJeA
xObaaO/lHnhiyc3K2g8+wgh1TUPf7KTKIRHIplDtPAQZeGB7bcqo3JtMD3g9s2wnEIfg27xDndOb
V9vJbV4agTmJJK8ovib+WjfFlqDREda2KE2SUvWtk2EqVcthFlXTC0BhQqTsN7aR92hz/uPc9uHB
0wtR1yfiUqERBkwJBkR5JpZ8vWySX0cT6hD1f9cwgrfoYn47Uh9KzJpRm9rwnYREXrhRT0X39gKu
hbbxzTL0t3ikAh+hsdWa511Br/xYjQyGSVr32w2MVRI0DtkaQSS16no0qjcqc4v8uUOXanl2QEYQ
ovtkG49FsAUDOcAMooWR0kME18x2mwlNCCm0IEOcMqLqobNUOVF4O0HQWkdasN39XH7feERfuoV/
EgQZOwjWHnrf5L7UQncmA1odwOVkWsERpEbKh2VRJ7r90KaVqVltQDfqU3r2zn+cOL7AhCHK8OyG
rUDbXrX3qXVWPRpqHPJfvrwvfM96IIdd5u+LU4Nv6o0fc6vhkbLkIsh9gFYwHRWzcYZAEIpU/eLD
QomaF2Iz9mf7SxC/DLXI4SelQslUF9yKHkGW6GRJEVot2DAr9YDdJYxWEmjuSJ47vJTyGw6eIdfx
Uc2Hjvy+l9LKcFOnRLfuq8HXMcED0sE1f0/9Lp4tJTyr74kxzb+YkAHHbwU44Q03zY6itWf9jLEh
cmOV2WPKwtPv2KUd0ti0d1EAZycNqPwZqu3QrynyVVErAQS9r8QmoCqD07Zzznez0utFy2FE2HjL
9zpKS8SWvm6YVJrHzKhgolyXDSGY7yFvBy+HQsDzEhMAXPgEJlEh7Gr0p+OA5vo3lSFClx8Flqa1
OSyY6b3oCxafH2rX2pGwFu4gYOG8YzzF2kOWXEa6DjoseAaMdYVh21huV5beZ2sOo1smUEZlzXrt
FPEFbSOSAZTA5Y/x4Y0wfH6XHP+MGUROGFd07YNIK/kkoM86sWnMeatcuf8VCXze4JebJC5RFxw6
2Py9DicvWie44jOVocPWhG0xkGc2ABZ9GvpweDFNXFM0FMNy+T8ZG7kAsbaKF0c0/rgw6uh9gYEV
P88lJH7sBzYQPuGqpmixQ+SgnqsHMmRL6XgyNeW0temj6XpkODeD/Jbp3PBapiMsB1IrVxxJshVL
bARi/bdj6OAFDwda3qlB0JU5Nz7jNXVsjsmIlNxQjkC8Q99Qojrg2fCR5caCmbA7OvThvlquNVIE
VyfUiBmnkosoJBtjvHmlalp3ZWJv5GY0p+6HzEcsve7MWfo2AXuWx8Qvt5VIfplIBi2mT7dansSn
UjQ5cpnRARELhICn5+jBYAkKgBuj6UFvqk2US6Op/+jBwIJeql5XhHgsJQja/t5Wn3L7jP1DULri
QSA1nFwuTtiM5eHDOczpQ5eL7pebmTxA3x2ZVoQqEfdG1LaJdoCgZjlZljkJpgaWzj+WiNy83uoR
yHkMw9kxaYfQHbhVtAh/f36/XxpdcgcWVrdsjmlevuhKNUiyx1mVcv2x9OUgyWjw2dQkf+ljeGXn
Si26oAM3vUBPih3HYhh0gy7zv9/kVwfaIiDZwmvZTSExuIpjo25ehj+11O7KsAWEN2NEDP8qWSwk
no3RSu8fVA87yZc5ZaAc5ssCNuPTDMRUxTdIBOBaP8wIQNDiEtoTPU6JGGuhnn3MZudHTAdJ1gZw
7YAo++F2wDSGXsXBdxz6h2ZQg1BUpJaA+ikOiJv2bylxmdnumByhBQ151gMpkB6l5RPPswl6GLAD
mtzr9f47/Oey838sjc3McjAhIymGvlLMWTX8HIGljR2fvJtwLMyonyI20gH0xYHNU5s2R7Xpd55n
Jd6Ae/KZsZPvk8tae0wwWwUGqUcF0NIoqRjGT4Xhgf4qDze9E2+3qvzTNJc1Jt5jl1OpAxa0YMui
siSs9/zBs00SlXdg2fR6nqHOLKjepXqfMZU36KJYzGvf0KXO3U4hA4ELHLVKCsF+tTffytEDmEai
p6gNXKF3L1BtL8yyr1NTqrfn5MeSt2/Us3BuyDlghnV707IOmxCjYs5RYQn33T1WIFGR7nkrO9XL
/8AjyDO+r/7ER8fbDT0PmlGXom59XD31lb0/D5C1XRjaAHGYmIqJxKW5ty5RKEwux17c3hdB+ck8
s0JLyi9ouDcBqVQaJnVwb/sWwJ9KgGRNx2wZy/Coed5MvDle/58FfwvS3uHjIzTm2kSyukBhbGA2
BBfQKOvpmbVsSm4+gr5x5lY9l2/fg6BZ9JqJ0Eb1sjDZQlKCWI1mIrUSlAsgMiUw/omZ0FYvuevC
xb+yBe028JD3O5En4zW9Blaz8iaUMLz0FLma3tIeV3k3VMu6CNLlf9P28HOnVVi+XlMJx2DEFlTV
2o0gIdEEhQoZyjl5u45U1QcAitrT40xsIBK2ZTGqo2FD5iDPfZWSQsEpiUEury0viEmJu48iWW6z
J3kuS52Bx8p3os6nROWpvc2Yrg8ffGYz9JKDhlZ3Kx0PCFKdONP2WMKdkaBfPqrlZx6+kg63kxZQ
jQ25d0CFfjtQIjyomhLA4my1ec2ncN4v/Hdx7b4CClJChBO3lJKYnZCKwuesboATSdQxsW6oUk0k
aKEZ+PjM2Jwail8a2i5MlxBZPs/t5xOeeF2j9eLW79jLGIM0Ft5bB6/KwBIjaKF4aU7sKuaQEFcg
wq6P7huekC+fd48v3Tk6J6iz2oYhxAsn6C+FqHBgrvpWcBvfqjGEBECtVpv2nNFtQX30VtFVP520
O000c+wfi3SiQkcAK7pygUmsuSROvl4b0j4OeLc13xvXxuBEEl0+pzPhL40YBj+A8IPs+cBXdolA
PIp3jEVO7e/F9olXDuCEh08BMnhfygt07PkByP/lmXSW1lgOhWcbHPVYi1z+DcSLsD69a2Q4PLS8
1PDR35z3oGrEnRyNiDJRIC9xCrN/4yIp32oCaKEJbiEUGNp+YN2ZywOw9syaiLV3gFaudQmYCdlK
YQsZoqib/C0nMqf1gI9oOu2zdfPA3P/k97+MZteawRuzWt5sOE9/kdnVbN8JflDjgj89U0abURhA
jf9N5Krnd0kMKi7UMKL2YcGY4GwzSlaRhsOcO5GSf/X0lfj7In0vf7xhRcKg9zGrCR/WS2CyZPiG
lxZkCQA4Sh0b1P6+Vn484Db0SN2hUB1YZpMhucq8MgYyWDVzQ7KfUvp2unhCD165owQ89czoj5UC
Wbo5hVYwVOAdOk/Mhb34B6APxCNEio7npzEOXVmwpdPDV2D0unMxthbT/rQBTycMcn7dC3/z0QcT
1FQKNvWQNcEHsFhvwO8JuOOFanyNp4iCq2IAMXyJZZLSGKlQc7zAAyM33Pg/VJNe/4INC6oW6pec
i0KUdX1H8iDsjbYibTZYn9IRdbyGUj+2TFAbrG3garas9hxYZXurARvXaO7ffWxboJWY6iiEpKK/
g0WX1oTzbjWsi0uOwRy3LF65daox+YrrRKEUy9ErwI0/1/RfhCHXCMXDHwl2jnL+QrdtuTcuVaSx
Gf89Ks8ze7DZ8LmJO2qgnEiqiVpIGjOEVB8meBeUv7SSAyddD2AUwAqa8q1OGFuOnZPYjKY0NrKZ
qElSixmGwVY7icXpTX0iv0o8ffxpTfw68pPZ/aFp4TkjpuLLq5b98XtxIEkpoCqwixAtBA0eBasm
tolNLxV/0lXQCL8FhcieOh6xJbpctf3G6aKLMg35Uji8AfL5mvTBvtpY72CzNd77IYU9znBNbog8
yzXvaWeiSGuAm0meMwmQYRAKDkP34gaFLpVl9le9CtSSw8XjlpzdimKX+d2dQpQadMeEc56Yn3F1
uZ0itFK7M7IYvoxnriTqYrOYgw6RivgnPjQV8KEKTL5HsfdwTXq29qYuPogxIzA4dHwBSIUY4zgV
WDlg1YtTo7p561GbqoRcAIPWajmBB5ZXO6UZXVF14lTpoCCl3Bdk4/sXoS4ridQ7vo9+U734Zrpc
Ego8++gB4wDtQb4OtPtmEgZadL4q5ohBfwo+967k2p4ELg0moy4QnNQvqRJmyM53xe7CPqwVzoLe
xCMok+d+JxXl9CUSuExyvP+msKUGEVh3eEyvB2TfZuXHOQhtc5Lc9lsoDlfVUWBoV6m8BIJs6gz1
nRk88N0dIpmR1QxoWJmh+253Axze1YkRbJ9s0uY5LxPjV1Ln8OdNNoVaW0+NxdmKS9zqc3/p/7k1
aFTWU+XunRcbTL+J6Hq8GLTt8wn6+txkat0xKK95/nAliXsMLPumRTm4W7iWuOv7tajYzJJEL8Az
Q225aVU6c1LyljPMITQjuMeU/MJAnjnQL15f/UoCBy8OYF37tHa28nQZ5sFnc1Hha9wU+7gMipCK
RyUh1yhJmL5eF4tniPA+CTOk2z3/C3pUi7wgcuC6CmrnxXlW1/lvpA95l+31NbZkkKLLiTWv+hcw
cWFdtAgmBYFOBSxIHj3i1LX7m4ZugDMRKO0NxOEu6dNuBs5wC60oLrhM2/ghh7SKh2cn2V4eqyiu
zfpFjHwgJiNlnx1YZw3BaS/4ILc9TxNo/+n4lI2C9K3JdFCRz2K5Akux8Bibbo2ELewJZ5vfxfr/
yazAEtGfMXnriVhW9/fZnM5U5TliGtS7xZlCCFK+1/JKDwaLITEmH4SNNGCixbyN+c0RTKQG7GDX
ZoSjBe7eCgjTIw5U/uuBnntDxAg5N+Gi5c/lycrI0CD3hYZUF0RGDCnsFju0jODIQokGEdu5sAey
PWNGuVb9NFHKdZI3OB9OmN8a78A0B4HkIik9v1/ql6xkXr6Z5GXolZCdZcdvvcBgdE5cpUx1qqk3
4sz1cREgFETG7CC7H59AacqyzM6kUiTeKUBqUHcbDUjS10EvZy44JeWV5WQXp3SbSnDvJYKsp/oJ
k5kC0JpFw5AHvYP2Q3YDKspA8eXDYbQE5109BWkLhYue3fRzJsu3CqjsK+QXGpRa/c9BbjqvOk4H
AUALmUFqsTYZYn7+DXeNcCpbkF7E6/tTLDjjnKoxA3NA/b+8lzGpQvmI4b1NranEaQeyroCvv5IV
DkeCmA8AyrE292ozrKOW7hCxUFjAQdRNiH3HW2d39/ivrfzaT84XxAbnn7/Ol7DBaGFQmguBYFhA
AlZPlEceQuN4KkV3VD7W9peQiXae2Rh/Oid4gynjTgQe4THB8B+WxZgpBAUIY2oSV3HuzOYU+3fn
L4fwvgM82t8KAtwdl8o5L+5oESH9qfgx3PF0fYwHKn6cHZLVPR6ffFTDifqrWelAq/bVtGNrKPaE
lNSK3l3mww2eZ6Bz1jjwZsZ3m03qZaZyUFfSrg5ICK9/pjYKSdK0c6Zr6wSNNAy5f0GXYtGDJ5bx
sho9Pdq8OYE6ojqCFzbs2+swvoOaOTLS3a5Ox4O+HIDVgnqlIMnJ+Xo5Y4xncnhnmWx/mDhSMlA4
lqjC6auBIsesN1ZFZt4VDuACr7OY2MZYVZBzVevz79ydFj6paLxpu5Z657qqzJuaDk9TxM16Pj6E
tXDIyXg6ZOJWxmMfX2lA0E0YbdrJZBqVFbWCEXPsPMXKfe8Sz4lK0unXcntyEEp5Dn2Sg6GxD2dY
ZlrlaniTVHf/4bh5JJVfwSHqYUURRT8RqFmB/q1V5lq8vo8c7cyMTgHYWYhfEW6ZtmL915jfC9Sb
q3l8VZl6lcqMUnpZCCM7oQSEdzZrRI+IytERdJtRnrqv5HiyXu3bBHHBZ5t7jNejYVebofFAreha
u4c/jCsm+ywop7CYrQRCibjaesR2/xYYDvcyEhS7/t80FOT/EZsbDtV2LOkfFWB3LVsM6gdG8GUw
v1hg3qpMqoM/2UW/G04DgwqCf2R8BvM2cfLDiKU5cbInMA0sgPmynTyF7JUDR0rhsuBURj/LXohm
BOZzbBYUyCIGrsBmuT1rbPPAe8AupMMp6ImqUqMvsBoTxcDBn9ZKdL/novje4HLaS3yIC9FPeLkQ
759phSP4i+6nf7XJvnoTr8C5jKJmMdzn1fGknzXLg0b7hsLHqHNlGdcZIS2JgohcxCDgi+jqqxp9
sVDOfjGttnKgpm0OsTTg6THnDW5ZjA2icsx0murSWPmkYFT+LRzwOVpTaeH2GuXmhIf6PpLqOOsI
K6ZUd/R6OVoh/Tk0V/nSTwnPfxg4Sdnt5t97TDY+N46bC+KZMg+wLThuw1BmHeURVYIIv0PNXBaw
GCXiJK+kA7wFvqKQz6/k15SUdOh1ROimm0r/J5r1EgzQYtX8gwgmpGKxijkvFKJ+6HQnO1BFXG9L
rffkFGBmCqQjnjMEWM8qWCgh8k3zRmr2Or5vR7YpF31zn5GwL0H+wHs/Jj1nAbhgFpSJlR0vp+cF
H8ehvsgyADR/vT/sCjjaKKakWhJNHgNSb0zWEjUR9FP75ZJmJ+3yh3ulusWZCN8EYAKYZatnZnh7
u0yaSGbYWMzX/iw04tRdX9zKOdGxmUc94USgvKRHPslwoun9CRG5fOeE6VV2lCu2z5Ufod4mYdDU
/ILNhwkTnZa5wEjSsT+rzdZSxCtfrxR4QB5b2UGIiUIXqD3xptJCsCcUb/AUimkSrs5gADdGMNFE
/xjE9avZIqtf9RlGMPQzl6GfzahZF6UzyOoOm+xnghnVh+uQonwl/eKWEYUmNfximOKXfPB9Hik/
vNS9SRkF2+c4UIwaYUxhEV4g6+4sNY5zOwz8f2YeowHQKVeGrqd7Pr85fHNepp3GzUNefD+ujNTc
eGAJlP4CPBhwGKPg3XlDnCwvfQvwtjKkhj1ehkT2OXkht6fMj8mG14npszHtIOJvuATj5ORovjO8
V7acLLDzV4TIXjFMaltTjA6oGYrGaZFG/pdwaKoxfxE1iMd2J8jA6uyfGA6q1cIoO16VzSrNpIVk
Z5oK+ZwC2l8TVWvG1kVXBHECwx0Sv5WNlzWtBoBNy9w8YKag/VAepF/Sg9EdSqyD9npBgDHnRvWE
BYwSC+b742MjnJnmXJTIAMXqr1pCy6WZMjeN/GhrnqOkriTyrOXO44q52m88Vdm9pFUj20pKfS/3
T+erZqk0nYp0isdJNqFZ2hVnuw1mgiiDSX7eJ+wuDpBAE04iDrDBmne28i2SA/fKNWl8b+nrorCb
Xn88MYDCVxwDb7UsIxdC0K4XK0ttkdOjp8OXGAvz7iCcdFAeiLZFneAQUhgV9LRb1ABHT2tMzc4P
likbrlxOhK5TYtbZDSyciSrQ7nbsOK7cPsgj26ysukLz/7EhSozhqEAdIIEMOFJpMNKqthtjpaCV
QjYee243gtnTbUNXF9ldkGsx2WFznza0cev0h98ArdhwWl/ucklr0vKmoQM5WyTqf+kmeucNRquG
n/GzHmNVb/zJiRggPiPS6ZXU9PnxC5j8JIRzmmyb6vwRxQlVCrTi8nQ1cVrwLuV14+PWs1W3UIh0
B3GZGrVgkkTBp/tsQi4735f1ICZpPTLo2qfKTo/7Z5JwIMzRLeKR0DGZb2JIq//+oC4OFXvQuH8l
eyA699MtTU/w8e+bCXPoTlXQvtBgZWwFtMjeTMWF+0Vx7B6A4O0cjukfncmgElSjt7jOnb1gG5H/
yN2UfMF+opBfyDyAxEVx26xnGkp4faGvjP+LAbXLgPiLnfuRpeU/CzrsAMecDf2CI0GikQlK/MEJ
B4LsZJtG/utcWOtqKPL7OYqWeVM/k6OGWZhthrGcPOoWWtdH3vLdeVufSbAr2Hs1HtOoVVWnEUVv
VH1HHastPMlIqbBdDVEUQOXB3XB41f4HTSTpW9DGnbzxYe5r6S4g4EuaTPTbDZGEhk6E9NyC1RU9
QfCwSyHuVyaN5Wj1XR6fXbN9pG6jNcQCc1qdlA70U3t8kYca7fAAQU88PCDRwIo8DiNe6OtT8ihd
xqmACo7PY7xRnUXBH6q6Q1uYP3ikN7hk6YaLib/qth7umJ67FlhoBBJIQb5chNQq2FcWpyf0z42D
nLlcfzfJD5pc3Ix2MW1ob3ps5BUDz/lZteGXK0u1NRK0B8PWr81nq5MJ3KaW6xZ9NIh17PmS5e0l
/4rpiKmubrz9AhCCcwqB0/sS/sulHc0PFxJS4Hq9oVDjUeGR8yyjQ/yFjrnCgJ06LocehcmTFKyN
aJ7pq4lzkJVPh41OYD9H7nTIOeVA45Qna1mCG9YKXajhH5DC8CBUVfc9wcmjf97KKHQAoVFRNvOL
GQTkQX5TNeL+3rTeVS6IAE1miRiG4adzjB6u9N7qRiFd7ERRjyRYoXOfLFQf0GaGq6892cR48aoj
RrPcMNUlrt/lnnHnVIbnz30OUwMhYd7+sCq8AaPW7/BkOa5aNyTsjXe6fAdfGwva42kbOX4jT4rM
J4Rc0YdXHOgmfUM5GTfLgCUWrvpRQm35gJs6itVOKyh+Yu+UO/m9oKrHNzODQZbwrpJL/Kk/9rOv
j3LglhEvP7U7Wm4cYFxBBiuFZnMwb328Gldkt6etUZOXiwNy2QuomQdzTiu5D5bjEtROOIBvIdw+
X9ia2rd3k1VDHC1VYM9N87gkMDdos10w7nRM8BF0c1i51z/rKqRfgKWrG7FwLG+dotp0ybaokmNZ
E92A38jhziQa5tQByb4TCtBl+tWQq+7RWU+EkQL5mmCNx0/j7Qp8j46qJDjRgOk1RUZIhHbJLfjo
jJwdS9DoLOhdkPKp2nUL5u73OwbzloQ+JryZMcqh5OgE8ozZiuB5F+X7Ij7bCYfg1jXac5TdUm2y
UXM9W7QJokVK7kWhUBJdk59JzHR9D5OANc3n/VrwsjC7YbkzKArKOjS/pCraMXB3PdN33/raMN+7
GRnZcWI8bTFwTye30hVGQ0mJHfyH85T8bsbrZot9vis5BrQlO0e5M9qKOb7c6hOeaQeblxUrzHmP
ELkI+4TEeEO7d0/pPLH4f26xFYkQnfr5PcRP6/PrikgTQDhlIj9mhAuWBP7JIxgQnSj2C0qh9pZV
UJrz7Vd5ilo9bEfBhByxmqH1kDgDapQ247IV4Qg96i4FVIqrnGTwazcHkbRppLJKwvMpm6/rhFpG
+w5PmMuZ0ts3+B6siFUV8ENjYgynW7KiMOGmcwWzA3Jj1EoBpFUXC0xKrqXTBYBfS9H48A+29EDv
tlyPBAcc4r/5mn5xMmS0ACA9OoniL2/guQPJ7tvzStYW28nBXzpCYbmkpkGz8VjQaBieBlMFei9V
MbuOXJfQUjdLNJuTL6OwJBumT3F1TlrIUKf2mqZYKGnFFjonFCUxHeeuDNEs/Cbo1u29fBgFl4DR
XFnMJh1r+NB4LGV3XJqdnK2dwW5oEjJudVUjYBvBcGukVTTwsNY88shyadDWPkn9Z78lKIq2qXlg
WM99NXiOZ1dNqO1+yRfAGCAnoNWrUBr0VWAkn0AWUtBB5sWIDdTR2vqHeWAF3kI/gqvN5UIMHwA4
ernP2JDM2XnWknu9lM0SP8x3LUkhJJuGYDcu4HUN1okiiCoOLPOsYZHwAUIO9J5QqFRkjPsASOC6
NjOEfY4gT8iqUy/slLqP9y+1T5WrpmzxiAUBMB1G+78OeiV8sDGJMIlXilDA/8FtlxuPeMTr04xb
geHgn2KTxuDRW4G31zslPrqWma3Doz288Z5p/pSDCivluJL+642lu/mEXxY6m4FmsbdhZuYLnh05
Cyy7lzEv808Nm82iLo93e9zRZj55FUTBuahMGtgtyx5agEgzugBDBeRn90DS9R3kAdXG51xiykJK
rA/Xww1CkpKsF9bzjiaNioa3la5QRkmgM2458yqODVgauNLx5d1WPEcfBtpIi/UXNTU6RDor2rfk
e3d05yq58+CyeYyJKuXccT3xbKeCUErtP2WaU48S36Q9vhl14LuBXXGcOw/QHvlGFfMNeNDKhGTW
T3v0snuut3G30VgXapf/SZupVZ3dh5VymI9F0uzMIklO+rue40WEG9JazNjMksSh70vLEal0zYvf
xnvScv5IjCgX4hjZNnZEISCa4U4Ik7/VfgzB2Ptd0KwRKsDqqeFwPa2R4KCCydarEJclOxpVOU00
HCAhMqsMenXrWit8izVsY4wKqcclt2cAQjpozI31R53X32q1mQsUvBtTRbz0T0GfE1V9X1q+Sxix
PVYrBuXj2pXg2FZ4mepsqkTph/cPXeidAGuEoN4SJet4yHeOvWfgi+/l3Aym/FeYF5XNuSain5Vt
xDY21hWGB6NN/9SX3qKtqNRjwUplLbLOGjUsvTs1jeezmtnylrxfKUAfR9VhmXg+QgXqdzv/EHtL
J/mPAUypTrA+iY7ll/RNB6Dqp+h2BkRonV2zhWpnwyUeElmEMfNtgaXYSvOzqaYE+hFKlEz5jiJq
wr1vug51ZRXkm6qmtB7NIdcNLphzPw5iF3hJMSr6fkzCKjjbbKWDsPKPgBD9FLpedo/WpP2gbklq
Vihuz41gGWc0JODRC5pqWLb/UHbtC0UcAKUJX5+dPMiZxxBrNmEkW7YQWG+ogPs1dz6D7GOqzOyk
TT9XAuU9Wy7MbDu5U3r5wifwG79NgASiZw53BjIkCXOcb1fnK/3wscxmfVakpTfPRFB7x/2wDDd8
X7Ga5Ex0i5ezN2XRa13DsI1QwfUmD4joi1/qL6NcJhBy7+j1Dh83ZTd+XmC0yY7FKu3me1LFFGE/
yB8I1sU1J2hdWawYv0PIVSCVzKHXBRO5ooTxprNcXJS/4uKWeWp0IVUkTUhllwxK2m/Ii7LT1PWO
O312X8+m1atKf/0F+j5uf6DnzmDotHwCArud5yOmLtsqCAaBJXsdtWYe3nDsmzmztHtB8G4RKn4Y
xC9CkKxTy9A7kCfCGN+qCFToWNMmHlXHq5Mst0nh9V4ZnQ67E2mKfNfNrxZ8iT+Yf/3MRILjBXUZ
D+0nWqUMVXBJJ4TpSxa3EnMNOmTsF6PseB1oqYE98r5BY2be6muPPpqr6y0uOKXDiWAbhXK0+GZp
0mjlMV+MV4sgLur78cMqLitqzKghOvhcY1yZ2VyCVu/pfQ+yERxwCh+a7+uEci5uy8eeU0lNjD/3
ptt90coEe8Ir/9SH4PLWjG/nuK1An0z2Y51aKlU3wYcE6LrEuTafuPEyNfHTfyRRwaJJeK8EMeF0
LmcPUs+TqFdwwFneygsdScg9TEVBav4HWB6d/M7PuXCRBo95Hn4vRXd07FBXyGDb5SPGzpviT6D3
TcMPAAuTutiltfmoQxWORSyzqgktJIrTZT7z/AKi+C1IBH5s6/j7I72zdHc/AuOOHH8bAKMw5wFB
Ih0zKi/pKi6Dc0g5r/jRGUz7D/rDnFI07ggZM4IXJ0SJfQZUQI2LxU6AYIX9gMSBuDC50ryn5s60
MM7d4LSvAe3iBzaIS0BbWm8Wj73njxH5sWu+DtWpgpSnFhEQRoBx+IWbW02auwh4UNlfWKpH4xpf
9ma6fuzStzWySubDEuwZTR0gBgiNiPKyWcEuQ/UU+lH9GVtOgJgn9p/rAqyDNY6i+0xrFR/w6Mx9
dn/oDVrm+7LFSmOEf3NiM/1cl8VJXSDvDAQiVvyNsy5AtJ/UsudiwkcchND5XvZQ22bUEm7gFdiz
AvTGxcYNJFX8jOvjK7kjlKk1TRt+/9aBuWL9/6n2rqyhDNAzYYQR1t/Wyv/0MI4U9VZlS/EjQlz/
aogTZIxQraGTBxldWzs6GlMEicDOMvZhhggw3I2pdKECRQkESPZNjmzQDW1Gu708qDYaAAThWyfh
i5sg/ZYoUxsa5q1GG+s7VB52j3DyYbGa7hQ++ZfHcfpt/odLqYUWmD256rrlVykiapRlPQwT5N6A
Dr6Ha2Zk8Et8EsYPQNj0y0e3MOKEpVNOIEKTZjCNCITX84Q0w+ZDYbEQIBpYIbfwDIIHRaMqHOBF
Rd6WX/x+GDdFZmBzUZ3/4l6NnoyLRMXs/Rgc4HBJUZxqR9nP6AAaJ9ztpxJqqk+Ep8nx6lq8PzRc
tVVWmHJw9BVAGHVz99bBV4gILaXBx2Ssz/6rJHNOo8apIi5K2Hd7109SzmYsW3sbocTmkXqC1xU5
Xq5bPw3z82xf5l6VFD0C/QjtjMRbBx9sLqRMLPij/xpCGR2PJH5pn9TtsLgD6ry61BTLV032mMKf
oeooXPhMQRVFbJCFu3g17kdSwgHqOreVS02fUmpwNcvU9mqfZBFGC16jZ6DxPePW7qyb7+ycZQ6W
Fff3WTGG3XrFvjUne8AlXfVb51fSszABQHsl0RyO9g1Ip3YkD1ZLVke98Uh/kSAx+TP6Pg8uwaBg
PzSQReCTvuwnYAfTLejZMfLxf8LPabTxwvScbxhsOfTSpeQ0m/lQYSj2enMM3oqyCOICDRIzJI73
TN4eyJZYe1Z7VrWBZFilfd1kBCF2j42QecvpJIzi9s89Cq5JmScqzdLbcOC8dwrDkLkUtz+bwnlJ
fz16s1atXa5fIpkkKTkXloDcVUzUgaTBxo8f8pF+GMTpLgfPxwpQPsi7baDcxI0pvdojzYD9UUNU
BXR6SkFJTR0SOMBKgq6csLy/uwwbjNuvZQzFpeB6MTrab8IkhZapC+U1wI70rb410cY2Ni3DY28A
IirfoQfHnIvkQCyQHzojuQv5K+WxsvK1ZFRNQv+vtErgb8LX59BJ2LleA8fJ/yQSH2NPevKx/U9u
RhlxbzXG8sUP88oDztFaMqygEY7tYeK8JCKEDJtFLji+fCL7D7MfHGN46qF40bzytOBjmDpbM+Ys
GRQjToYC8Ll3uyXFBeLXGguiwYsguhV/VFH9j/a1fmv70mZ8fwOYCfsJlZ/ucvihZB5RYFH9++0y
VwtdDWRdzbeidtyeU8GsBTsRJzprgsiadkJX5nNXKUDyyyXQP95h0I3TqHaEjqDlZOXc2khhQvNN
Swc/uLhKyWjJQ9pcfqFRwYhvdReZgmA848XV8LPc92Mqf7Y2GBkaD73YHbLFi9h7hWDOZtlIluCK
A1lyWfRx9kTNmShYuj56MA9MwUBafKvdHaZvoLNq9ogXonIJ/vVkl0419sUhdSVlajwxj7cGpLY7
Gn8aC7AF5eF9mf4e0ofPRaqjFBvClq1uS98rJNs63bObCc63bmByr3FI4KYPLRx/rcoyoIN1ZV6H
YAD64NhqWU1eVLjftIiVU6kGowphhSxz7tqWx6kdvP73Uaikws6nAhLJlrEhryv4m5wIwh67whYZ
xCdydTDg2W5XrWPd9MSwLqfVs6m/YrhZqq6oUsqKlxoE/DzZ+Da5vWypJiaeIzMjJtUtRX/pBHmy
Wy8UvZiUbNnC0spwHPumDNJrR8Ui6nEdM0nzDl1+9PVqrCHlQhUPNjom/q+YpBi+LOsdWKkZrMVS
43yR4MaBsWkIIKqtqD+NQtSyowXNwNESWmEPHf9SmI30lR5aCloJ6oLTHk8iR8zXrdxGxUHMW7zs
An3AC9i9cmbfRb9xWyxnGkpymv+mdSQfw7LxVAcPf1EKSgKSucZjqwYB8/HbOtCs7p2j9rR1R1OT
j8T8+cS9BCm3NbYn2IGrPqKJp2b5++RJdvACJ+hGbMrWdUsHi5zx7dNIZwtqDyCfOnIqRMADjo9l
j2AhNmkoEdBSE3YRuOfTHAc93NHdzTBXTlc6HCrAjVOnckst0ETGlr7yy8F6ot8GpV4o/P0L0HHi
OxqR8eeXJoLf7RtLEMysI4URm8Ok/qOUX0a+RxA+l9zXY6/2/K8aBeYlbaMIx3V+YbAQAfo6HpDP
WsqgDR9VaHWK+Qjric46RVn6STUMlUolsYvmbPN8uk3+A+q71Zqbvn44y0n/4Nxu4qcr4NDeXkVS
YBg3tdXOoTlXvsBmua2vqbU3sBQlsjdoZDYZdq8+rE8t2qBVMqlYbbwuB99i3Hp/4GDQvJmOq7xt
k2m35AyDPLln+2x8RbzKG6WWpjg5xG+cP8Ehr+3PlldGuSlKdILbrIQx0qUBHvO8pWdI1owWWzeV
mJACjpKrx0V4+lwj+hq3eBdDu7/frOC/+HrMau8bVaCVkLPC6qi/3Mub+jJKaA+fv1TwNSJfTDQp
GPqDxzNtI0fTtpT+Bv5xx7fivlI/J5tiOV/yB+92YGhSX/rUia3sfzUc/WXTIym7AhqwttITlDn+
1h76PteNSiAfJLzIolueFAulf85nQ7tnjv/lOfWsDSQ6dOI+KqOKIkIU1FDhhL1BT9p4eE09BHV3
3iwmIUAGGFCfi+LP+AnV7p7y3WPM9ND5JQIm8sgqFliaLjaRJ9hAHBQODvYyhByuDejwW741zcOD
2820j4lc/OrQ54P7/4gLoG1EKosJNwYimQivIvWaN6b6bx92KdbxFdeiqGHaQ6AE18MQlS+Ksep/
I8kdME7S1lpQnrBmxgu2nhHPM7DHG1VClewL7OFBpadRrRBY2sIcaU1z6jD9DQ+cLiPQrEPNsA2h
lUx/85qjBOGlJkP7qfqCg8ycjmBSm5Zn2TFJsbGoVnNtRkx9APyukc5mMdWpJIyDlix0zgNjMCWl
CPiyrk3/icpAPlr3ZLtmyhMgLUHM2FUf56AW7vDxLBdj6Ej29EDtxqItdhCXSRdnswt8AyHT8Liv
Hez8vcbt7p04bytGwNMzg1gq2pxT/P7uPux00wqVAJ6rqP3AHpGek5xGl8KV8XS7s7ELvg+z1WNW
1GEJi2upOQFO8SpPauqojE8X1M9p64W5pUiHxI6u2/n8TAEHT+bHROlrvkedu4m1O4JfkTnnlot/
bg27+W4MLDx20ZVS191K2jCosBSFLDDRv9AI8b9kTQyiuN7Q5mwTihE8OcrZxCECxPGw2JsCTT2H
KyuMeuBBUlnF/T1LZSHVE21DOaS8iRuPZTuxUT5CLS9FR88n2uKk44whPa3VC3Uw7vLE+kVPJO/e
2E8LK6NhuJGBs/vqYfZrJoHBEuV72myrJWlNokKCKTiD2OATN9T4OYTI9uHqAhixIvlXALmR+34k
dihg4TnbbEpz8JKfMKFxxxMebkCZ/uevZ/Ksk1neyocFPwErXFQ0zX5Z5wP52CMJe2pZPKu0agYE
sFeVu7HF6dvWdsOeK/AxsKiD0WExb+4gkxUZK2RJkXjzZdrqvgRK9H1AO3vLHx/iqH5npVPazDgo
1W6HDJEMuDgORJmeXbPlTaKyp37ZWjVFhTFvzvgO8PcnLp4218tiBoUjQ7jQ+NVhk4zuGM19r2Bj
v5PPmz5qvGDSQZ1RtRB6Wjb/3Qk9i2rDAzjzoCtmgsG0baI+5gsoJiXLKWiaLQelYMVGV3tHGdz7
ZFX/CUTM2hzheNk7lyB35T8JCAGkx0WWWU11nRMr+VSk6fsnkFM2aCfBIG6RF5voShEncTr8Sn/a
D+HVxeHH4liFnE4HqTW8yWKOZlkQbAoQDYuO7MjBB2++X28xMIDpqkJYjH0tWdtleob5b1dC2kZ0
H4pwxz4eOnh2KGXOYG/Vf8abdrtWNpa+5EyKj+5zbBiJzmRqrQrESVTdONb+57E79Nazjjc4vVvY
TezVzLanWsA1Vahb9/xdxX4sxbAyExf0/sfZnpH4t7FhUFzyGX2iv+HhYxRG3+CAkTa9RWI7kUJw
LPef1OEr/YCPE2S+8GQpOoZuidIEk6dLUjykJsFUtHCOc5BnNRocLM6tudnEdFqQwx0wrUACfsiW
OhrwYWJIt+TwX+BhTwJml0iIP+ihBocwGehnoisQzPYCO7ITve8VW1utdQaBp3nCfZDrX6xIddlt
zRs4kF5lHm0fJt9hLW8yyIx2sgeGw2W3OJY556bfk/tT8QjTktL7IkBUNieYgSSgPgEoQKCI0P56
ffTLYnmAWE8BQPMvB0YtsfXR5UgxtoxlqUElecZ0YvM2bL98RGBnDgZKMp7M2POnRW4lFcPrHrk1
5Wt+S73RV8b2yWohKb8kss6860V/j7UFL30QlJNOXCN19P/9odc0jfBmHVysWIPnGhdrJgYgXQQ0
ak0BN54JJ+Wwg7waZpFdfGljqyWc7rT5xWKiGS6SuLjFOi4LObWUqknSTfOLyUCwVR6avDXlmPkN
slIw1HjGRI5zf3bXjvd4kep7NWwiF8+iZLckIkNDYePdRM3gHhggDMZ9N3j6gOBfpJG0SdncXpEk
KmDdY+QObIaEG7fmY7kyi6hwy2YUc0D9DVj0V+tZp+GMYMVfl0/lHsxcilG702PPk4jQC4N+b6h0
me/ZNOPz5n6dV6uyYIf+N5rVuYlmBS1RYVm0b/6BLO14tER3lxBzmKzhlPFx/7am9ORhAQPKwLJO
YbUFn0rkNjSVxrWxuLGjgK+HDr3ZcB9w81KKYiT5BhpSrsfYwGLaFrl7EjJZF81zSw/PUwncKlDm
nW1ubcbtO7p5qaoo9pnus0auMQGQRpp3jccEJkR5ouyL3MOVIl/KqvKtFmsWNlqKXtOMAVnbwX9Z
/NTSgVOBZXiDONoLfvtNuez2A+VK6Mx+QK0Ig+XN5eZLIwBTRGp3//QupdzZePkuKTyb2LFLoVdt
hItpd/i0fAs/NzoP0uy24QiavMeXNE6AgEpK6kt+eWRsigA58xmckEAIObTcaOlOlYGtEZENDB4b
uCmsR74+xLE8o13xQN5QlmmO1wU3UbuV4mqaJsrJLbC/imDoVSPgt4efqqJkdi1SWd3Ri1YBHImg
sM4G0BwJ8DCQDRaAMMAsXPXXH9ij0B8bqSJi1XKa9l483rHiaitIDztL2WL1B8GIbY/jjxoN2NqH
QsPu7vvKRIuM2y8KvcAAmeopUu4liRL/XzQeda1k0tL1zPRR8hLE7Gsx1n78+iF7SD8kdbwKrRn+
rCZh8Z+aG+lcreTMxyG6RUUSodF5OdiohhHwp9dP294HMIcE8YJQS4N7ptiXndkc6Coynmw6clys
QQqNDPdD0Ts8QlMLLjFaTSKybUaJCR6oU4dxOPX6BQMfCqeCCilZ2qV2r1NRFroJJCG+Xnfdxx0S
sD0+2n254bSCKOIqp3msIgAfMbkr4jgCR958LcoA0YdPUZLnFNByzX0A7NbsZ16gIgR1uyMdOgQh
PhA1ms5b/3x+gSqAJ+2kmaqISvnzj2g+YaiaZI7fP1ZRIeXaJKBSdtD85Oad/xfqJXfQZ7wBFf/6
mj0DzJg+Sq0gv0xTPKZv1AqZcKzKnJVzIZJQEtMtjjno0AtQo++hrV5ws98l0juPM9lu7lNxp+s8
O6pEyne89zPZP28lll7YDeoxNO5cDoAzqoufh/mS3yOOkeSmLC3wlIXI812pXCScPWAMU9EX7KoX
JHjwMmKP7lLA9ReIVGUS2NxgsTRqQ12RoByMJhdKjTsHPir9r3EoXcIxwsCcrmAIF1uccwPBiyaw
KMaRsqUsD1bGMOjPEnnjlVw+Tpsj2zEJuqxeAkhDq0VCAaUq1D6pR1eISr7BLgPzqSpNZETWfzYU
ibqeFSLB2T0V1z7xR1u42102SmigQdB5DjmbqT3zKNVFRlKJGLlrdQtG2oXukgJlQBzaqS+x8WVU
ooG+IaAbRMxXTXZk1/iMEoKkmNsn4I7W2AgDip+6PSkKKhrvDA1GkXyPVSkt4EHnPCFJPYIKwHjr
kzbkhVmWJbeii9qDs+DbUzZU95MqmbIBq4UxImHA4j6Pi8Zw7Nnq0cZuadOndYnJnnDuphEgiFn7
CdKzZIIKeFbKPtvbSZTnf3otEsOsDgzQyZeRkWMX11PXzmh0wdGZiUQtu4CprE52Z0NaVZTxNbQ3
5XfGIfr9CiKqybxQVTLS7oPdmpj4LgQzmgOeNOrAVNsI2IJApXAqJEeE4fgHAFSAniUtT5/WCz0P
+eJWipM9aOee4+veIf+oxc2DjtOaXL917wWGpwLe8JNsiNsCKe/nqlULzjmE9WRUBJRzWhILqCeE
rHniIfRxl1gO/hnutjbLVkB5efMP9bfGcxai+M67naOn54/Bcgks7pgNvL6uOe5KRjGJVkVsj/8r
pKmGBelL4vJuXer0e58WdAAVMn5CpffDWp63nHX4p/X5rsod0nsNibgInNs0O731fToPa48HBtXK
bjv/e7Q+WLISL6iVo79hPfz08bHTDlyRRR4YWV0quuK/GUjNR6im1p5fnKEu4lazqW5KsLLFzS2r
qfiA1mO4oqhz945oD2ou5ChlsSiZ+n4Fm5yAurhxA1BjZH/ceItWBmtZxJvwCToWKvGM0qtIbiVY
V8Q/naZLZV28/yimpePpZooqozsU0ojpgqaZTBOCC0TAOV9I/chMk+xowoRBx+PcDis7mB5WAA69
377LgULEmoWeEgNNbQ2autXGyBq4zk3CBf1yjDhrKg7u4c4kJ1Xxagz3iWj926RXAkkkMuWOLMg6
n6A9mmQVMcup6I6xvBCLVwybygyPLo6UIT/VyjCXYX2VGwpuDzAVVwrQ35vmPRR6wgoiTTqnkFJT
8xdKQ2phHyPJrgnZsiuMxLhMV5olF0MI/iUKtsjxulQo9oXvIqi/GithPDp7dgP/SfkErYpW3v7g
J7INSZtT0NS1+8s4eYTYcif8BMq99bRo9mChTv2pprTpcPoURwPd8xKH64iGxT6/Ay1BEcK7I5O/
zHB+lIt6bETEiqXHRbRsgGTOBEdO63WVPYIXWp1SMVHvieLTUOwJkUMT8PkPieIpnGXfXNm6Keg4
jRal3wMd9qIugy4jZNkuWP0Hw6YsZHp/dXvTB6VKTuDYM2day6wIR8rJPP2b6NbMq6ZoNRd96mZk
T8vqCz7STsvHx9SV0kp1qSNNx21N0x/LC/pAFzgPUdyafzGzwF339pL3lBeSdRIuWgYiNGJRoj/+
IU552d4uVQYpCn355Ki0Dn3LbIiqTur2ZnVRgxnWOH3o6tlc81pebYsPqPek1RiQMy/i8trJkjJw
aJqEWB1/ZgE3TCVs8RbVoJW4gp7q9KlKADWpD23oe6DQHZbMGwCluUKJdORUAeYm3ORUu/yA2rFe
fUOKmLB2zY6OWq17Oh85P3MmNV7j0vHjua0r7VrerCnWHCRrRhe6LeYCPRW8U7T7Ww1x5jSJVllS
3USAJXFi9b7B61Jw+mp7PUMTpWhKt2kVGChZqHJoolEYTJIOF1SIIcn6GbLEfH0SFzSo75+5HHJL
XjroTnz1FQW1hNV3r3F7nGEo7ryVoNcY++4WtfeGfoSXBuTl3ZLZpBDaEhrJm1oucemQfHFQ5fOJ
Nn7PYbEz/TX7l8VvAiS8GJIPgHoBn4Hle/yoFbjh4hIB935vf1ULrtAQ+PLwnxm23xM9VNn3S8Mg
0Xfz89P+7sj+3QtAC/mUkZe0AMPWc6Z0QFKWG+j10pfI/flMD6bwXwSNJ3M5pb/ylFttlOEUASS5
5lC67ghWK+kcPTGO/2Kc0c3+yDI7jvy3rbS0XLEF7xoUXvXr0okOfWGM8R3oRZlMeUSIQHEZyX1k
XRN2dj3z8DDT+9D7s47LHqFtbKU0gm/5jgMjmhYHYeRFngs9fmet8XFje2T46dn/RsmsGf9lK0Zf
gXv75xVxNxBMxI/AWajVv1CkFRGhfOO2qzNEFFxbIjNvmt4ntNoj+jDElg9n42hw+50ylWs33unl
B09aAQ/TW6UWwUs1lcz+ph8vfhjHdDTlmikYK7nDDshZmr8jT9ULPWnUxY7DDIugRtc1f0GdMuFL
B1KClqniOGUy81xY7c2VqIYK+uDo/UhEXypvc+1b0L/6pwwWxrjG87kxXZO5O9FaYpMgPM1mujK/
7AIc6y40WCgadkeYuz0Fj9foBmOd9gaLTtBYIkoGp8n0++W3xmGcQlD99W8HgLUQqY3Gk9N/JghI
B7D/E57LT+DZFvi3PIuizqxjyw5JHVEFrSpVGrId0qDGFJGS/LTyN8T6DHdhvDpwv8ellk+YthYd
1ChTLCu6QXU3yF6OdyUbEDJbXjxgswyZT3bReKt6L3vB7OUJeSzCzb+YM0uJ+NIEMODSGlcGOVHa
3OBKAIDVt+B2GGOJY/89vpNhH/JMgVsjSoqwYgZYnHaTpymRUsrHN0cc9MlsNyXtNpan/DigxeEo
2tHo3PcnLC2J10Gnd9xYrKV1QfxIHx73ihm5K86FyNKKuCbmuVQjJLUzVHs30wnTv3raQd+pp5Kl
utQ3lSP0j+iFj/m/yf0k2nw1xJesJvcw0LwxvCkpEd+IO7iEFF3E2Rv+reFCgFokn677zIOUnuBo
SV3zD8sAOGXeeGxaowp/StEtVqu37C9DhR/6jGtO1kQxt9k5Gs5f7kuC5cezLo/MCJV8R86IbIUR
pCwwt1zDcq9d7R44589JlO7gWCBc4UCSmYFmrb486y6I1pjatFHWQtlQWJMyDWSqS/p/cBt+do/F
1ASUqz05s3OSGZGkWlYDdFelVhKE0bhrYz32EFzpl4MJH9AswH/RRtUR42ru/XecnXZu+/gJsViX
JOvHrWtRMDgX0KB5kxc8K82krnzVceBEx4Icz5e/sa2zaTOwaEpj2qW6IWLnYtSnekNaD1GRH1da
a1+EuhtZuPOeMAIvWYkRAO1yd/U04dPuYyLu+IjvbSk+oeowsKpB3a+FKge3idVlir1vft/s7Wf8
IS8H/vj8/hDPxiyZMS/s2GZjwS1GdFEwuXJOXslBqrD9QkU1gBjqcX6gEpdp637JbZu31DJVRgm0
mQ9/5+R9J79zUfVSuVPbP9JsPVSW2JXp++p9L3fqh6rlq4RnAmSMJhwqzmyKNN7yIlM8yitAkV/p
cWhyfQdCGp2r0gOjWsEwao7Cy3ku/svcWzDZkl/VLMGhSloI0JfGMYDyTcJoFrVxZ6sGPAY9DgrD
7QT4ysaCv7ERTAG/WFvlciyuA4Lmqdy1TtslivukaDT3rJ/rCJgqAB0p0YvTQmGCksptWlY5PPgy
BjS6NMbnQit7hdFPBdUdlATQ9+itTblVKt85cFeUyIwefSJccAlLZdbziJlX6Q62spLXN+zqnK5A
mjgSS/3glO1KQmAbHN86pZeXiYZo1bMosZKVwEPzbUps2Ab7zCRJ5+HovjmlIpvdUGWn14o0gs6P
o1WL1RNsywMnr1DfDoPbj7kB36mP3pLXQM9j1L1+6/kYz50jKuVr4pcCZL6j618Qb3FuY14OZOKC
rHmNraCXGTOLo1xbQ0nHqpQGq9/leQHOTE2CIyqRHW7wCZLUoYepSiLKUohan8yJK45jM+jXSQUw
14BsIqRBY96vGns3Ub6/6XtH9pA9bBHfr5VfbHsKupw0Bu0BGHaQEzDBHBB2DfLsFtF7sf0XTDva
rvP5ARfJ3sfeNohmu2/gvlEUpXN8G4HbqrVtkLCweSUMoP995xnsADtCiB2JYmZf+eJ8sv9BaX7F
+UwdmGVDzs/Ldw4hLBm1/UGmJ5bIW1SydBDyJc4UjEtDfwdo9j/bBpv2lRIfr6IOOcPie8KDum73
g7LKi1Bu5ztEwtZb9vGYSm76DZbnmguNiRY+MU11e8JiZGzlNU/FTo/AZvMznJVyY1iiLqAvxyic
wdwu49Tv1gRBnQRu2neWkR/vMSqigP+eXG21l2xTCWV6eNLdv1PbyrPwez51HKh9c8igZvIBxyNA
d36lpE6pBNM1RraLbjpFiYr3U8Q90IspNDDvear6Y+cv8hyh2DUwiy8oT4SlIZfhfDc8THKAxoVv
onkRDcobm9z2szghf4JlJwJjMNNB+/pxJVi3s9Ppa6uACesZp49tayhddFVqDMzKNzVnGPFF7syw
bT78rrndG+2NeWT9vx437X6k6t6MGUKE3G4EUylTFZ+sagz/bvRzWvGZ0JXAzdy8mSzV1ZHJzreZ
a3dLmfTk5SdPCDoEQk0Oub1UOlv0DJxMxSV6tIhwT3uJWMUvf3x99Vj+Ss1NsB5LeKPH1hlSvtoB
r1gEtqvOJMLtWAuNCM6RFTMnAODB7i+bRfWP+0g0hSf3FFXQMRttECTvxGBzxwaO5n+MXMdgTEMz
g0gfG1CcgnAPq7CvdgEVgiF3BSy+H5xM0SQuHfwFbAPRSqiTpMdFj2ep31oswSGncQCZl/i9YL1X
W9KpVA/xh3KXBgJebGayCN+ba11z/AcvGa21bYWdxqTN61CYc6+PLhoWjSnzqE1YZZlr21Ynif7i
FYeq6D2JbxD4aVjQUwQYXowN4InoPvAfYjtAh+4mO2H3LnaVgMxuJA5lNILEzx0tEGqKFZ1uWiQ4
EDy/7DRSCDY4HzSNKASVgMuACN5svDqeQ/9oR3gSyMTMKpMSLrVrxfmbFr3G6dZKyBRdrhAf12Yd
rxPOvSo6cPIykkk5scN4Rcd/4ij8FBNOp5P2GbExuBHUcUyEyu5DQGy0/l/vn3nBafcRlBPGhxX4
hV05v+7HTsFLQo4ykZlzRMQ1Xndrx6oXRWnryfNirxqSjHXe34LxwuV+PyTtC0SiB+46ETsECxd5
0FlaFSSHhCAi0ZMOhpS2IZ9Dq5ETix9cOq+5bO0xAvEb5o67TFw8HoCBy/4i7ZHMntfKOtLt/tQ6
ZLrcJ3W2SLWrzxubYsGaJih9aQ6n2XdrGc021NGpmb7OmzozmhSjmmnKTMDuLkAvanFJgBped4SO
ZRpG51Ij6Lml77PuVWXsqovTaBVTvuFxkXX8PzhPFIQ54iJHRQPp+z7wKygghxanYCWIecUN312p
GIipo7Rac+Alty6tyaaf4EVYBv9vK5Msaz6H2Dlav9PDEPo4loDUGpV6Y0zkLOkpFEKUCNSiuDyQ
1grQkLlg9C2NhE7CK2dkGcEOMOrbwQoBawJukvgZKefJd7yr2Q1yVhoITkIwdJ+Shfv3iVBw8joA
1xd6yl87VL2uJV290/DizyZNU/BdM+xHxja87Ey2E/8yFUC9xiR7CdqSmjrIMhtcU0JJ0qu715Lh
8zEOazqX2PqZHiYilWfq6sXF2JKkNyfGDbcHRsQVfwSd4Wp/fBJYShf6ZXUcELs9h83Ik1VGy0HF
HhHKEPhm3M0VZo1yTIuPYSrHPJjkftm89OhHuOlY6K88LUijXg8BXLj3sHYPORg96bOlXhV+bv8y
hHgdg7cvyOUahQpd+z6gKkWMCVIzLGvbEo1dU4HCvggOg7weVhWXWQ9wI9QhyuO3Ez5cZRemq8Vj
DfyZIQxrFJLQyllkGTZpRgPxFnpXsj3OJ2Czs0J31aYn6/9z1i7UauqskynEsffSt/Xvi2imJ5US
HvR3DsqLElgOuZbh6kFWqzVqYW5MCgZS0Mzv8smuSecRAgkU7w3gDQIINb5JgPp3s4okQwL1NFeX
Tu5w0qoccOJRS03R1DwPuHUY2A9rUrPcS+8qnn83IGgMc5JklILhVLVV6SAgYm4Idj/osdXQVBcl
oJS8vyWT2vWUsw8eDtOZEoK0alpgNbdfxwUbKp9PV1jkaCVJA1vXjeXYnzWBF97Gi44WM9FLJfUa
Jkk7j8aBBCdH/5q1QJeEufx5SSaNAvQWWcU1x6/AJnnxet8uqW9nvUEcfLZ4WKeH2B4PIHnIb4dz
L+fENAiZeZUe/NrVR1qCkWhfvK+m6a+qKEuGWfPYSwboMQjHXQ+f0lUL8c3bYCHW6MpL5NRSN4dQ
kmteIGOnaaZnNZXQP7dQiZQASWRCR+SuitTCLgWyfE3GOTqKgDGyqZ4+nUGadLpUm765tFHs/WMH
ZFakwt/CxHOrXrRQRMQpOTH5D4U47yzqAoq61IOp1xn0ASjXw2R/gaQ6xT16EM8CFfgMb4OP/zLk
PPMQNNZg23f1J2E2Dxy+9cLZ1gqlZ5r2oZASBYNUpC1pzLtOjlXbEZkg0kYy1IcwzqQ9sxmNyNNX
ZmyGmhtv+na6zO73sGph0tNl8l6P22MXwFjNLf/Q3lJvzNWoV6ndg1SQOxupYhT1nSV4G16Hu1/d
Z7D9dootHXKAFTfuT4tYFP+/iWvJIwEXYlUT5vgEUtxMQiU0nhrD4D+rf7yA6HlmK+LjUhZbmyT0
R56fpjNUMQQ2lDShCwPTgut2f4/Ll6DifYemJl0Y6kMDAEj/djipudHUcyFjq25C/3mZDGkuWK3Z
LfdCBh0s/OkDHXngMhNWuLuvDvmtaAWJRe10Q5bMGSnGg3yFzn8XKlS7i/sqY+Mhrr+ZZIhN5MPL
0yD3URo9wLL8aE9gqnyCnIsKE9BFUMlEmSDUTK4IiFfbyhycWqbZzfPpJ7Al2HJhTITw7fPF5ifk
lJ+X6HLQwIlvGt2yPqTiS/cwsOkV1XjhPM9AhNvf8B3o+Sr5a0ALtLnHzEDDhx+oNM6lWB5OsqVQ
Xw24L4e0OaD51qC69HCEQzEh5VEhdCfSx5tkwbu40RgqNOmA6rvepbt2AGG6xGuBqeOR9uUijTJ/
gbgIyidBI13cUswHIiRNphlGr7iFuf9IVOxdjHIVJr2AHlSYC8c4Sukw1WpoukH5/tzgdNzWpdMH
B5N+B45GA8frVqUMV+Sx/VsTVC4iJWOyEbBObDBuufRFH3i3fIIPdjpXnMRyqzHcyLiPsQv5B+Yx
stD+RMHZzWgnyzg9jmpPwdH6/lJcukIv+eDtlsp43ji7BQkoKIhrvVVVKAbLkGS6MRFR3JIdXBjh
tMuFAnx0QSGepHeva/uuwYGUBPqqqjWY8ENANGG+F63Kvh2l90PVVhDln1pRDVjOVXT3ba5gsorY
1HGuX5XcTmgSLwihDGZ7QvYlalyCisAL0QeiTdvRE6L5xJBFh24nH5SHjBWrWjd4lg6BgCpgEcuZ
KqyxIEX9mGz5Qc5q9vd6kIbvIyaFX3XHJ/CnL4T1l0IPNl7PB5oY7ei1SwvOEze4fjjXjJiemUhI
zj0gP2oEJ3hU+occN422UFeEnRaNLaQEiRTzm4cEdxNmyo6LlfCgglPSeZWdawvxWJYJCdk/BZHe
c2qVVOV8nxcFMXW6lxyosrTImvXjQVrAzW+OVWekatRf8pT1lG3a+OLGwCJYUnO9ZEM4Dl3qehJV
gSEZFyfqYJCg4iHeFtclcV7CAFulGJKxBHiGLfdWr20qoBJZhjL+kUyrffiv9r1Bkfe42bvsdqRE
iK4pgLYc+k9MXk5vXmmxX/hBrh8ItMYGPtgBuZSRqPZvtUXxwCLQMpEBsoxQEa0P38ZkZEO3qBKR
A0CvVK/4zzlHyk0W0t8ct+A9FMePrw7Pj7LUc14FvWUZ4WeSY6uIvj03zYHTli2crXyxmqNTOpV1
SwgzMvbTu9Fw0cw7CNsgfY4S3Sw2aHn/LwhnbvJ/MhAZvAGZpdH8TUOb3YwR6+TyZEoBdDakPljX
CPSgoZmoFWaVHDzOwJdvFC3+iKlCs9iiiMPIZrCr7Tx+5kZY6QXfc3GLE5v/DqYpdaQQU6oP3DHw
sAffholcv0DTo/Qfu3qi2eWuR2csrmGrzK41VGLlvr2ttBNUYHkfNP9m7AiMfsnyiGCPfUU9o/eW
4gukVOcRQDOE544cqCh9WVr5CmNKZi5NxaDBj+qtzAfVz2M83+D2kaY0DYC7Ha9OHeQR44LA+CLg
PwXs+ve76O9qwsQTGmYsDB48Fzn6IKo4G7Kulf+/SPaBocrg29Vc5NY5GJYYBkE1RxLTpFLcjBD2
6hQTnngPXTbrypq5DotFeDSBmu5qe25khWAWRiJPoDec7EkXNleRDNaFODBOkSXCv7YMSBQU6AAZ
k/5YdmQU9Jqg0KKLtJF1tHi/XOEx7uNA5oAPyrlycoxMQrsLz1kt4SHgbI4trsIVtI19DBlm+PM1
ayBOIXPUQTBRLhdk+OpyIMcKRk7tIavlLHGwZlAF8HQGKjoJIeJrGYukmfFJXYjuiOoDCWanY3yo
HjI5s777IoB1yQ7LLdlogmos21wy/QGqqXKBGo4y1UfzQWDbIdVr+R89nvYbcMMuj2L4igY8k71b
7SfqvpV/I8sqMLlNMntyeJNxtICsClgw2inPJ0ASQSJVtMdXqDk914MpIjY+svq8KRPB267/ibTg
nYuREh18WgelvpMSvrNIhkDnZnSJUTWGsaPtIuKF1iDyMzd+oRjd5dGySLUR+lwtgsb0Ce3RUx2z
r/n1NXZGbvKvcd53hXeSMFwsqe5tuE1QAW+HD1sOBjaH7UNwvgoPps6/Zpv6jecCoXMGI3jpx2x6
jJoeNTei5WVn7ALKXh1D+O7eOVotBc9RivGCsevQGl4y1qs8VeFAnm5GJwng0ve0sDV/b3ILecFd
0tD/aHTjOEUy2yRN+7Yjg2QQnddRR0CgcKOIzM3UbbC515A4wFI27WhEFljRkRff6/52KlpwhQqO
G4D8wSrTju9p4i3USUhUDh8CXXnAWGAAvrQIlFqa/ifgmLteXEzv3ya1WoPrdhw097xycGVJHGtJ
99dMimKXKdgKEt9lw55Ewy2qvAzXlz7gfWmPFhQ/bkFbkrOCLjsAsHXAgc3HF6oCrCaM9+S1sW7T
RXjeMLQCQKioGDMy5PeWmWJNx5TZ6/T7SSRTImjeaFJFhgFAiZfnueSxXhoUVkp/htT1D7lH9bvE
gEodWYOdx+89+N0sNPObN8aaPa6WqKUwbsS+d+D+etQn3PfnOW69zToVjx9NY61S/utJaJEWy8fS
AZjVr/LE6HeGTzalYUmbaCADQ5AoRYbM0W7AlXCasigkUqmcr0WHz3Da9Nrh29/ad6pr8DB9eUjl
tBHp5rHny8zoqzLuwGICwtmEI5FXxB4ZkcrqFNlyIWcH0EFL6ea846mz8VWdAK6HfMnoAIJQXxNl
QsVLhTeAkffGM0ORbco1aCDeenSIVmo0hK7NE4sKdBRUPjzObRNH1Zp3Cz2CfwFye2ejZlBQcp7B
xS0k0ZCVys3TUINcT9jRYp/kVw4rJZp82FC0UoQBZN95HRMsaTDlCW6pfhltt6Oed4Vo0rcSMqqA
FdvgBEP5vK59NGc/0A2PxjLqc8tX+jcl/SOp5lhzHQhL6fTDPDxN3DNzIUOazJBCfpbKxABdlxqz
HdGiiz5eLoLKbEki7qfWrH+EDmDJUNMjyUOYnAE5xSkXBjwKlAp0oHpwe6j2Yc6F9E8HT71Rn3a8
LMRfuoQymWN2FrpgjB2JDr4vqw0ktveG26eyf5+sF8x85azrKqeke5U2NwVTIeuGcaMVcSJOQ3rx
lpoyEsmBulCroYNlQEPUzrJIq+Yjg9TRjCmgVnQD6tJAg3dOB73V+ml17wpY59zJoMtp1hgKPFGD
+zMJ67R6ffyDbEqjHv59EN9XHXe6Strkw573sARW/8cuRZdem4+z6Z2/OVUFd1jUmQj+XIOq6CxM
PS7d4BmbohmLCUmzVFIbiNIrBTqnWTgFtLje7pJ3DBu3+jISinyFnJHSQLbetHOqtV4a962J3leY
3hGEHahydRsbX6Vcg3zVii3navp9oXVhhI5vKvAc96BjGrXNMAWxsft8ZBR8PaMmRM6dUkgrOArn
4iZtKGAd+Ih8AVHpe781Y9p0CA7qw9a9aYQ4DTOcZxcg5KqjBKnf8qpmmWPphM5BBGU9A8SJOEWR
QIl93M/ZdmpE9Gi2LOIM2LgTZPBFykPScJ7V2ALmVGT023IcxnbHLnwLzv5QUu3yEhjOt3U1vKWu
8csPFa/urea0u3YW3nZoZWUGd3+4e9lcI8HJHYNeO+kDIK2cEXE2y7pbFm/ltLqLl8vWNgp6uNtY
IBogSuTIratDqmxRyYEBiNoMpTSojViNU47Q8Uiv9682Kcd2eZctcmhGuQ7+e2LOrLJeNTTv0r91
tq4FQnJ+S+ptPwYWrT2DiH08Dm5+K9CalOeX6VxeXDBTfttalwES+9Z3YGVtbJMCmqb1mZ1GLtdD
w77BvQ5oICwOX8SnQYUgHGE2Lmq89srH0dTVzGRKvbzM356MF5owBmvRG5Z82R9lHbrQUit+gKV0
QjP1g1Fdf6icihH0h7meI8aawgfV/UWm8HA90JpXAnIXMo3tSi1WeHKGW1im9Mb/dVVcn3MNwCr/
c6n2JTRV+WsznXfFP5yevszDjVdylbpl2sSpuROJn3LazJxRdeT/abgOxfo56BzDUP12Kx66YeNa
HIZ+IU8kVnjmTxNf7s4fe0zWPJqK/sRAy0xRxopEfQxYD8vXzhFfPYcMc+iFkCrF+I92sXkVMRG4
A0tR6SXTUFK2nzdmWhUaJCAuhPjPcfQPeAibI7wLqVUwnrwKLhpy2LWDoHz4K1EK/6SZyX0MBXiW
hx0faftkIyMbC47yKyg9qS2NbUkICDeTu6euZX3j0SyRmpuz+fNnaM3CAfukm0Qzbazeh8f/Jy82
uHRiDenEPuWUNrk3ny2vp8ZfHTPtz8yZOF5tgHUklq+tUDo7lKL0f7v8p1WLGCLdC0QLdyA8twQx
Mi7IJy2mOiG20owduDguT3ssz5YI4rCFO0Ed9TxC/Z8s8iwYwz/h4Q7S08l91QBmrgzIen/Rm5Je
CmViyukilpOFPAu4TD9G0XDfNOAkwSM17lyOuL4KLF35y6dtKg5quQ9d1uus9H9WvBe/jC5BzcDs
ggU+N1v/xAFJK9DyOK/gFwnK90b9NbLI5lp75lwx1FlJIPB20I+6Z+ayaLe2jJzvu5RVLLsOKPxa
PA5hOMFRiXIeJRHy8/asGJfnjqs+edJaxuQdtm8bhRXWjb0zrR5KO0c5ChDoP89JxlaWriw31EwK
x7Dk4b2JOSnc1FlDoe4o8aiYynVsuE9mxk6ip5/Ohn1+809JapImQ/B2GhXMat8LdXBgduOhQ2JY
hfJ05Te3TT6R9U2U4dKQDoJAbuCdqNRupLE640eYtL0GeKcI6B3dSPQd6jZSumHoXDKKmkdRCrTB
SpKZs5qHVvPv0orb4giNirOv+V/xQF+SIHRk1r3UI+3LA5EMvWzhEPBISzYpFb/Ie0tWW1QsBGgn
/MRt8p2wjPguXK5kWz0JL8rt0vuzuURNeqkezCX5j7+Q/QGvwGXB46v0UKkIT+0PP3njHTDRsmVA
Q1FGCuU9dRU9rHE4YNRybb9uPDOWRy3qpA4roOwe/Jk+A6Ghiib4L5c6/hr1dJGfq126A5r1fPeb
gUXFvOGegUDuFzVZe84VELplUbd9sH1xHMRef8ECutY4dBAUYv1bmM8n10HNUtZAQvsTma/LCL7b
1JERD2KahDssZ6o8eAC0sUXgEZP+Bi5LzANQ6jj7jq22xgT5SdJn0uN5p9wLLl86DmvtqkXOshcL
uuNe9wJNHmLGlBG+mjFlaMYkU8Ip3uRtuaCICuN3frGc1xA4k4VBJK58LCsQbusfwson/TcEF3BG
SgVbXMw5XLFlYgGQlQCVMk9CobI5aY04GjiTgBwY8VQwU6nyi/DNf4xi2NieX2DfTcNo7sCZk2qx
EEwoEBRzjKtFH15497PhMwNk9T87kj/dF9TeD6Z2Ky7eeSdI+EO4pOWN1UlbOhaA9MNEU76Gz91E
OMyc1aW57CA1kGMNEAddVHaKrnkiTUC904/WPpVhdjnStBkXu/Xg6+HquYUJquznbyCgot6L88Gk
cergQtlgs4t6QteCrIPR1CAcbtrhGE80OScP63Ma0lw23cfSUUTxsex76jcopvY6w+yxJhN3Q6oe
ePzAVO2LUMk1tnXdsE8cypxh9CibZrMl/PHevORCbCZYBNoSGGCZIcawuu/ve2cb3ZOhJ7a0rABP
IaVWoWmamxZuIpu8776gsVE+SRMQcZ1j6UJ9peqYjWwnWhG7pmfHZz/EVOWY/uZ4AMG5l4ppQyPu
yEw0rKV8xhv1ZhhoatHEwE01VDIH6GtIXYfYtN4dGbgP/ppTPSY7Dz3kEv8nouFO0icoEJJ3A/RI
YZDuuajpGJ3XfyLosJlS9Pv8+ZNgXJcdUvj3Vi4Cxogf/xC5C640MxqhD1m9IxrTPKTrBPT9q7kX
tgOmf0//2lGiBNpYzt1dUCcbD9cA8QuFR6IkkDlnyJaUaC4NBqu3dzzfKhBrEVJ/KOox2k9FMlbP
37mtFH6o5WAv8FTYAk9qIipQ23MavN24oMHT5WjG+E8ksjSUmMYFlfeVbXcdB/s0SrJ+QyxCzvsV
2nYI2OxPPzCGoO7I5I+IpoRDUNO+g778Vbtn57aSVb9GNLYpXNTZDeActm4IvyQW79bwkUFBMbCg
u/60vo92MIGlvBkbOvNurgFQyE4lP5BBVZ2CsMo42QELYxT9vr6znYy9C2gFe9NWsFGuaiJ/ylUY
e0DTylAB8ERkgtOQVvSGewgi9a7fbx+6l/PfrD3VeIDiQwSen5dzwKTEuKygI9O1fmhRxDofz/r9
aDm+FEWmpzDVkkI+6wtbaT1pMeLVSvKvvynQk7F/tb0HzCfPaovHV1pxaXIEavH4NMF7DnyIDfuB
S8Wm7DJY2GcUPEaIW8CpJorhlyDozBZBJYkp0OBnPytXVDXmbXdklsQbP7jipRe/ewBno3LAfin/
jIO0u5iwgxEqMIBNEXyjKK/tAXME84uxiJByqLyf3H9+dU7hqIqRbMDivueCNR2hZREZ3kw1fY0p
aVlD95PfYJWIgQcRnDm79qe63QAA0tFSjyfPKDvx23Hkdq94kYag6qZr9piDo8LC+S2YEG37/FVu
bAJPS0MS2lNCitUB3eEW/qdmFjOIFFQFkK7nrC68ckTDkoN8dlAlFYOOT2M4e7BF1bTW9nmN45IF
7hTZL2PLdZCwUxZd4ZFBZF0z6JMoN/Dl90LGtIVq9zs39HQQMDxwSalc97sDZ87v5yMeu0h4XwAW
ay9/h202WAwkzO0JMZKN20VEhszUQNB3ZLxGcfWZ3aXm8/HQx7TCTk1Ymg/ycQuws6vp106xDMVE
hbAQmcpBWFnxED4he4+dJRpjohDaUgtIs9tkpjJnWNMmLeHhyfTSDakDEk2bH90ELkuWE1Bzvt02
MbUOrKlW9OME+zAvG+pVuZouA+dOt0BDsZCjMLxTniYtrc72X78Lpm1Hs8sqy1Nz2u9ymuNZ9JhO
I/takOA5QmZkE3GuH+UCVi2R1vf54KubQ7YGJRV3X75U6JVhEVI7WF37QMw/GDwvSEtDFpYUgGoQ
4QJUtKeLjjjYPxsgkyMwtVWZKC9VThDsTW6ahfx6bkjzbUyiuK+av2zWgjKe9X1j3YaiJpP6FUlL
+AfORtyrxBMzEplMb/upu81L2I/7cUE0EeTsUee3TT5ZeFUDVMkze6UTqJiItypChOwt3orIp0bW
poqsUC447zefw1E8fIwW3lah+CE/sdp4+CNC2vDaHZrAMHlqzIcxBDFBj5qAFpQ0YPhnqhpTD5TE
S/HCzILHyGHjbMCRQTSZmCX0+tst+cIH1pLa76fQj00qBiyR3VFAyAlZvQMfP9QeTq8mNWwAlNlB
1OntHCj0o1O6mx0ypdu1f7s7r9V26NDqk2iJqzGQvF3TMuevS4yIn5xZdhscEb3XKGIkfEcHHHmM
dq0/u17VNBJGFBF2hkdRinaiBfpbWLwk4FJSugnxcRSG2Zfyv6KtoJRE1VLXg8CD8MjovO4iIIGC
2nO+AokobYvmalch2kXyl/KrbMU+JFLFboadS3kIjE88YLSi+HKSKaGdg+b/06/7Q9Xw3nTgMXZq
tOICkPtT/Ad+Nhf6NhddF6wQBtUTUT0jIU0vznnCRbjHuhvxhPHNaxQ9jVw5I/kZLK2niYbymc11
R7+WvWYLqKO4QjBlAwmhfWVrpn8qoc+NhgoUq0L5NeTy5dkB9MEXiAt7P58mge/YIqxAqnx5zDMX
UQ14aHUydLJlmswadyDKE3+CFIVwlkON5V/dI2eJRZhXMN0NX9oIv9OrObqAH+qCe4anmKQGBI0m
8Dq4Bz046b8OyRVYOVzB3jO4sbS2jEtJmf6F0i6bVJWmtfq9xRxI7w8XPiAowM+PBmsXqKMQEmV/
qoPwq9b6Cf4KlaNOTg151Jkyna8dWOYjSupUKjRzJConTPq+fu0P2A11br7MwMA+qV+zmCnnr4MK
g08LLLKyN15KqtTXDj+S4J82yKX2yq4+XnYq+nJdycoX/hrbXq7lJwwHiVm7yqIHHv5l503kr844
VlG4a5pR7VO+ZyfJAhQ/XRemXoqowJgHhN9YRbcu3uuTFmqjSrIk1bOBfPTgqBpkkAAiumyFvghp
D01XiTUs3Fs2QC6uD3ey1B/QUxcB9vuson/nCdY7YmOoGHghNmjNuAcJMuLEn06z8eLFcyDHImlP
WgVe0ChT0HMsOfJuv7Q8itrPWvsz8Hz2a+bqAi120+28zva5BPlz4VnYzuRI0PRQ2I+vqm5T03Bs
vJ9BXvAkZR67ckYHuJVv54Qy1yE2BX/XxUxSeGrYWUqr15IjIoG4TvwerQU2ey9eAQ68IR7qaple
G3svxQZjdkJW6WCnsR/L9X84u/TQBwaDoDP6Pi55L0M0Wmg7UlSWHyoOLcwvuxBVcrUHxUBp6R4v
AE0PYk5ZGlKgD2W89Q2jOEuAGaKlWau8mAvMZYlHl7TYLxfTKirKTTB00CynHQS/M4giPuxElKS5
2k9UoaJLY2jOkqTkH70VeeM5T9uceD/g+TVqXoYSpsqJgExLntVfNy9kYqRrcxWGKtEJlw3XkpFB
ZYMoFtWN62X1HX9w+Nnz6Jemm7mLmhR7AEhOxNAVPlNjM8VKRhl5gPmSZudDhMT/y9S9hzjqM3wD
pCWBCM+sAm0o8nzJFFEx1FkEkM5XN2YLBsvxN12vaVY1Iim52k7BB+qOxtAXi+00U5JckoBku9Lg
UCo8QAW90XH6wkHOMaWpxxHLdnEKGLnp2AuLP1PoAapyZSJlEFXC1pJFUCA+WIBoG7GZxqLMH3Ea
qTHa4VFZ85yUliWR0h1i89rIDZ+Nq2VGsQuIyBpaLNtbJZYLG1nkG7oR8P7i24D+kRi/IVr66EZU
CgbA6DpqfH9LHtuTC0qAawefNMqNo9Fo1MB4QZ5djiS0EjYEoocKILYqBMCLr3NXs2C6yexF+qu8
JgpyozF1HsoHVl8JNk6Urc5AoKryuARlwhIpAh8ckCzp/pfW2QS2Ebq6eKCzzDIGxEaxFf+4XThM
hEOC6cxS1cfjq84USND6OiaoNGCoMljLw86i7ZxmuhBsQA2JSoSx2zGxGZZQZGF8+Iz0grkZcy/T
I/337BGA4EAYxUZgHt6S8vnc7nOqe4xIeW1SEZ3j+azQsmhUrDs0GLhO8UbDBY/3mNbibW9IFLbX
iGMLdY/XQcpUZNoW9+Ng++HXVLtdJlXgbG6kOiDyv6diiWtGTDLH124rKn3Jaf3eIp7Q3YQjjzVw
bKUjiXqpCHSCjE0I3l0RHsixQpH57C+e4fMIehnQdx5vfQ2KaYlvT0fxD3EAGZxGh82hnq+QcYOO
0HJExFqaIYByJB2Vqxu5DufAMRw7h5tIiUgLTU+om7NgDlqfOzz92nq1IoI+Ff9IuAuFdAKz5xOr
QVYl/Mqr9MSM/LmbJ3e/cFAe78QaKmX/NwbDVIJE5aRMVksoK+lwaEHv/BBpj/ResjivtgTIzeUi
JoeUvXxapjxbU+mrvn47MRR81t5+BX4gaqRbmYagK5XzTTVnCFnGBfbZVaTZ4SAObT0a6xaMwFK+
0jHQg/8iMjkYwsNHk4QdykQTjwoyAXs+Hl+1q3tvbJolgC68tMkvjhKG3nTAVhUL/HHIUVVlY2o4
rljVcsFBCr/Tx4ONDg+DfusqYxsAqdSn7jc/obvAfzbeXxNSvZM93V48AS4tPqnIVpTJM/i5VxIG
47BeieUFtymqg8RI5BUcz1jVzFXOMCjEg4cHiD85TjezGaSV1sEgavrcdKism7vOUlj2XOWUyUP3
BPdJgV4giIbOcruoQqtfQQG+3hADGfyAg0Nc+fyKxd4ivR1Bl+6tp5jIh8RWfwIWh+uFjh/+YgHe
66tm0pPfPbhL4D/tjglzQVcti3QbKFqsbLdMyaHOn0qDmnqEPJ25Tkes4gQQNlcXwYW16XnCtKwe
NaiBTg5yuN+kEUsR6cdegMM1XlK5rNAhN5rOqXiDEZXuGX2ce2jv9F64f19LCTKF1YpUebL4Mpy9
XlnHVH8q1yQLVuJziwxKrHuq7JLt1+1Lz1yi+pEhOnwNVVSTuy2n6At179x4Di3rnJ9pxbBoh2R5
LmeaDqwHMABcuFpOAA455OV9lPwPt2IYb6tS6hVU8huIJo5CquL3n+rQFvpEBVqGjaOW7L6WdPTk
2IxdjF6sQqJd8H6fb0XeyEajHF36ZtRojBN1nf86RjZVK0lAp6BkMxRae9+F60wB89l/lrRMWyBG
/1r/xSBih5xzaQ0Ar9x8v1ddOSWwA1llwvKh1WE8jblfiZjFoVWN3hjl0O2ecn3aXFKm1Egxg78w
pTTpqt7cg24/7rNmf43IfSMLOy4CWB2wWU5gsBU+lq0RdoEY9yo32gnCyWwXlX0SNgxrL+gxw2Ej
sfzMdpoQUcFYJmkgewtkfGRaBfU2Nfwcy2N5yRdJ8/5gNBaayKx5ODduICGQisGdki0vzhl/E/Jc
Xtokj6skIg4KA6dSDNVMysYEU9vQzpkhcbjP4QmEn0gD0CYQmO54DvYlizER8A69vM1CZzz019Rv
77p4EDA++FKUfTqk/WMcwHL/zA8tfdUrKb860dN8iUNxHNnw5lFh3IA2/T9vqmLOZRo/zF2X5tgD
pl9mrPpFH9REep3IJ4XQRdgX58eN1keRvi5Hsvx4TCd5uOlWquU85qM6VIXpI4DI7looUp9n7TtS
MQitnV4REBY7UEvYs+R0QHsIhT3vVVfW33zFLEaiQ+2i4isdfn6/BUq8dPUA51odm7DMY5dUb/57
wuvWc7kwLy0/XOerJp579cfa1ctIKOa/7echUNAbaQHfEKx1wkYEi9h4e6KhoI1akU/DnJwHP40s
k7FyxjP670VmkBnbucm+yG1Y4WVDE9t2THwE/RSAU5jrL3/HFUePMIAN/etNTopopPmSxL17SHHh
B5zRi+Cgx7eugxWQYyGx/wL1rUBYheMeoxiR//3rWdaC+GIo8GUO95tjZqwik/mhDyrRrS6nzgLK
2cPhGaL6BH5kEqyGB1FD2ryIXGZ1JqIBvbqqMOhoDMbvTXLlpRaUTC3y1OtO81xk1O5CUsO2N7OC
vFGdiETAxAFgsNZJaosYuz51MihoNbTRc+GZCZIN84XHvYX29oOVuQaHiVwYS7W02Nq6pD2J3mf3
DQopNgrSKdWCmidQ1fGwZzawqcH01OHK+Fbmv650cFjhRqb4utwHaPrAhRvXTopgm6mEGvYKU/W6
UlJ1Un9oPsvRi7mcevzv4cnF7wogUSyI4zirMCwn5RD1p/Yrmg26wU7FU0d7AYFTZ9dZ3/DOL+JX
40wYGSn6E/1SIBfqRZNfliBRifyJulR/CyW37Vcp6qub70Z5GYCNM433FnEUgZztr9dKBvEyZKCF
ATtof7peOgg0+Cg5KcOO7edkoBdtoP5IFeXuhPmbpq0S31QLVAY4XToszlUf59bK5TfDlHpQDRCr
FruMX+ibNcILch5TLrt1DehJGdA70Yffcwne7IVlb7yQftfb6d+NQEPZDqcYPSkHfKSf5V86dMWH
edUlHrCfWszJ3gU2FKMeTMWQivNwIdDiJBv1wj6M0C2iZERSb1hIgaNauDoJzFkR3Z5+XgjDo0vA
ZqTY/qCF0ejpdWkeAdAqaOiRJsgw4WYosHTslJEhv7YJyNq7AYJlIOKBLM608nCmmOXgx2S6ckvD
pSMp/J2MC2Ax9frqWVhNZtpAIv1FxFutEAMXIb5Gvw0yDlYDpHVXusPDT/CROxP2P5PuqxnduLX8
7FD+jwKGtQLVg5c6/qDaJLPlxbqZTU/VJCiZgxZTK9HiUnoycRaFaBySupcofnrsZxFy3KOkkulJ
fFjkUCmoDWJj20bH7CgxzXGaSKg1yS0qhlEtT5+AZ8qdqVNxK+62a31D9FoqJLziooo8g3kYNy9/
EW+3plhnLh9bx2oFZ/8QT8ZealvzVdx4qZo0sn0ucmeAFY4vjHZxwDtjM3YNhN+tLKcGZZAGqDok
J/BWus/VjxDubQy3Fgud7PtGLSfhdscVXj5roTIqq921HSNByR7D6tDEDDaTheVgx1al4up0tKBK
edch+L2d+qu0LTQ3jY1JLdGkKESdmdkA4AJmrm5O28UFCEItc/D0FRae2053wwT5ZeLC+OvykOQB
F8N3Dw8n2dRkkCmE08SGs3s9XGUN/Nzwufa1vhxtlDzJukv8BgRb3pe4vUZE3M3I3jPiCBriJwCH
07w9BYI4yALpvy38rBhWBz2am18uiWRTmrCYzwT01EBN9A6Pl7R2R6fFgCqn60zE8Rx+TnlChpPQ
3XnSigue2b9jcyVbhx1HkPkcf5OY5KzRaRSciPGJXOHJQFxXte2cEbbsWJqglBDbgkMQC2W/DXE8
MbZ9xrmJrfHEp74YMprKbGkXiZsMWjpnLzfU0x8xGpBikuMPmGJZAmWEGDPC5cHJ4NBjv2JAgyhj
LG0//6fzViNrmkoh/hRwJhVxP73LL5qfTfykOqjOzE2Fi8HWAvd82NlTOqsoiwIgEeMhV7zSsSnK
AptdiZshJkQVdgjz5pxcgp1U4BqQ07V5HhfddEsZw5WzDLcQjcASiQKLtNClU53G5cYcxGT1G061
4cm5wmyojZ96fbZMSj9K1mlOjkYp/UZIUNXiGt3aJibaiYhp2Pha3LHOloy7LKh4bm3X3wt7c2K5
chtLtTMQ/7I8UmX8oGRxU0tTjagVtBsYnvt+y+LpawwEeMh4Zh9I9NSN/CSbzDUuHa26stODUY+N
JGOhcn/5mWi4bsZDMtJqWDLfsgJ/ICtq5oo1zhqHGsX8VEOAbutRoOcbL8/KAKeUHKDDHZNChAk3
/GU59nOI9B7OHf200LS1m5OMiY7T0poJy+oN2fnar0cs/hKOsF6e+iOvB3Jk0Yh5COs5ZDCIiX2/
LUhZIkNyLK1tmiptGCsxBKnALdT3O+CuOfGRa2tlZC2c3ECbe823eFxWEsws6OxJceq4FfkbNZsa
jTqPBTBdsNBEuBe+rLzE5VPWo9Tz53cKIE2kdmzfWL+L8smccVfPk95dmzP0DYG1K0gSsfKcQNYO
qOO3PyeGuGu6/bf/dEizEzPQjW0FREwjiHs1hMf3LtlzeY+HPS6jaZ6o1px+A5G1doyVOm9g5orf
t87M8eOU16Up+H0GQhPg2PS7VZZdzsxNmE78HCy9gZjvKYBZSanZwPvDgwNryQwFL3HiKHnpsazE
3RZ9FI9AZS9Xsg6afRojhIyuDRkA9Qb/FDe+xSRAI+Jl8+r6rzsT44k9M+zyTXkJWaZGDsQWuafJ
7caUNIjVe0YPve1g1do8aA5OsVF+z8lIt6kyVD1gDUlbkh3yq6zZTZi2tbMpBRJEa+4eTDPqXAWA
+LncFQwVkVE9j+GxYpOyNqEiHdGOr3vNyZPUXWjTBb4aHUm3kJArkg0KhYDDGHdoa8iW9tGpcQkU
qrW80UBNNPnPypj1hhJ6BIyjQp0tqjCRYkYb2HRR4qM9Hq4/1eNHDidCB2WhtnsFwW1yFnV1eAsu
H26UshVRZ/kBfIlwZGimfoZNY83sBj99c9ItiBfpet5lGOtHRdBzDXobaC545okJOaXRFOD3xGR9
ibFI0D53G9iupJSQ5vPteMNNUKLaMMdCQNgIr1KCeAJrkywvQm2M0jrUGvKTQwRovhHdtXsZHlNo
b1FE9LYpAVIm7Vx32a7km6g4KtL1mcXoyl36aLf8zfB2qdGvZJTRq4Kw9+S9IjQtFiO5Nf8+MObI
czT6pGOBFWviHJf495AWMNlufGyUdqXGkT5B25YrXPen4Ezrpd/4cXiPPxc8QGrVoDV4Q6IlB6Qs
jkWSJ0Dn6NLdhx7QHADay4oq51nI31wPkUY/GqPqsuHPA1fHCHRnWIl61tCx0FooFRyKAtymN99P
caEwgHtyDjNdsKZlfpINMAsYCcPGZ8+ID+qbrKCvuhVj0WULR5QLcAoZ49xioz+NY5iCMhfPuRld
kq7GQ5CJ0hssbQ9MxN2pChBeVfpY3v4IjX5/1g9sqCVQAtwGs03lexGUlf9cAEV/W+DTfNYgxabs
dXQR0A+aGMEGB7ODKpWdo4fqIJ5Yu9o4Zb1L2uIA/C70tICjqfRBf/VSFKKIPTD8n4xfcvaX8POW
ENzQoqVi3f2JkleGWxpnwGPahNAq5x+/wziCbYiuoQTfGyQqw9R4UFQniOlwuKqeawitPfKO8iMm
84NoMnmzzaNDzDa50RH/more9KeBkQ30LHMnZ/yy3dIIXGXAxMUN1bPVHsOqoBxZjsiHhAz5Jb07
AabWUurLNR0I0cKmd4Z1EVCbaRYTC+UHKkEp2vCT0nY2wxKaISyeCu5lU92Kc2GqpT91rLSwYI2I
iRCJKtyMpLO0I3sg6kM4uxMV7L3d1dD9R3CLhXegp4bAU339buPD5HdkZYGKFXI7rWbOK9k0xZGE
+TjPre4C/xHFGXyC9uCcjsL/8wqyA+bVsHBlXsr+BUOOKcm9XTBza01MxTxZlqC3qny97xqcUJsi
8BqjjTqYx/aoSDXb4tt5DdGuhwW9pWRmXuALRcyUvt0Q4F2WQJrWBn3y+kO2amSl5WxLWGl5qSxe
utmdk0fCdbgQIdEevPwEfv8Km76F4PUnmWF6/5e6BbsL9vpsRcjCzUluNpzypc6t+piEN0buw/+w
EDR5Y/yIHLW8OlzBrxIcYZQYXoPiCpD3UAhGBbQcZTo8a2+TVmcnkCTSNKDbO2vGQ3hsg/BLa52Z
mjUrF/Phkn1YWmMYXyLAhP/OpRVCuO9ItmjbSUahdz1iDtsL1lJ3RkQ8oQoWsF7G0ucW/BI3W2gr
T+uGDGS2moP7z3Xcf9Va4VTy02Ct0LFDh0OzoeTC8wHIKf301/Vmt40irxQhN43Iiv9FT1UGwCqd
+b3U/1vJM1btbmo+xWkfohsOIB7fjt4Y2Vx8XCp2l5t1Nuvdjf57p8elR6l1qBdELP+QImVBegzR
wRKvPKfLsDiYynUjYAGi5M/7Hrkmq73biFH2CcP6JdXQGwEK8eq7eXU8vmT94sOkZX/V8DCgMYx0
p/BLZUFgG98rFissay4/gDDsMmvHWBoidShpA5bXZlpKISkG1FOQpG6JKLZXybq72HK7ENwja09m
NXJo1W0fWxFz0Cmyf+pzXFA10pf/FKKCzKkZg3hhH7HfAkNsCWb6pcoX8JwFlBiO05EUjtMXZTzA
tbmt3mish46Yba1mTRnGzTTOMUwZH9gl3gmFZHGo+RNmFqF2Xt/pfyfPfEPOjtm/6H0fhZxjttEz
Go6E55CntLoKEdkUqPEptB13WNR5TFDIFX2Gt5iPTILq2bRy9mns0L03jjab9TMYpedvUXW1iX1o
8LtE5kh1vyJEqJ4c/iHqqAskYuUSUy6eEjop8BiZMuHiS6VoqBagLWr1Hd2NiTSZR4LcLHTU6I8L
RkVHVLS3ra0k49WUreDXRQrKrCgvT1Ei+4LdV04JWdbk9TqsQdyt7jzV3ELy1/2bVUcG9ALGXeHH
+qRNa60nDS6yh1uxb+E/fThPEr/UtIE53irVOXKsJocAAQLhwSHSbdPjszTve7d2c5cWG9PkR9F6
c6OxNiDcORo9StMDs/2+DPGTb4txiD/KtDVer1am+Kf2b61l8+a7jRWRbFAia1osj1w16BwF8cmf
7Tq03awU7FA43okNEGq3mJmd+c9iAXtTHZ0oTH9e/5mlGtWKBw9gLh+iCE4tv2ssAugG3p4kxJrE
2WqCK9GdVDFc9QYK5vyNgAhIFyUZYbiEyRkITFPGpcML5+hDE6ZDXPAMsKVZfNXbELv36OUnF2Wr
QkD73OEsmo4Q1vreLvd0eIzdyDLQp8cuCGlbgtXnOdRUVAPR/zgF4mMEKjdvMglFzaS9/XKAYK3p
B7DXhkC4LoRbMUk6geJH7c/bqmvC2Jsv00ZuQLbjQ16vJl23GKGRonFSpHJfInlUoB0jDnGZTLVK
HglRugDfnfK+uZAjLG5gQbqsnloXXypQ2jGV3p13YlP+ujQeXWzqvHpQ0lBcyslZKQWsJv4FILR+
UbiD9+b3BBqmXDcVRvhUSWDGvQISDjbFElJHRGD5BUMdjV4Rmf+DqznmMLB/4EVnxJ38rObVBz3Q
uPkmyxjOUvW1MDxq37+9iUbnd1+K+Qf2WHs9s+16Tc6f7i3zsVNH6R0n13yBR8slC2YEy4WSrdKL
dD1OUsHw/0JXW6vjH25DDpEuHnSNOco7B+SgciFL7wUtiG9h9gQVEvwkyzrVzIv59diQlxgV444u
+ri15prelSu/F6hO8r3tQPCJi9q5tB41G33BF1SpYeU2xkLmHT2+53dfdo4PKzERdlqkGs/9Y5iu
hHiWbCBU4bhY7vhuKinr+L9wY4Yw0C7DB1S7DBxJjCnGVbW1R+Vgn7xU7R12Sj0n8d0IZUGg7Q3y
xK4xd8tBGsPdDfRlJh9ywh9lZLhhZTPYt/AA1f3NWKEOiGD4xz2TYUwn99nIAP2zgdKaYKmKK7Tl
6UOnrndgRUjXUY8LbM0LBKfsYgMkkwpk6woX/hHcAUO8KIkF1GdmwnShtgnFiz+2dDjyE4CHE98C
jWVDDLwks+iVGFzch6UIEcuNpsoLvWQzxwfuSqsSigN4WsavzIkQGRiBugYcFXK73ItjFcewGra4
cIhSwnI+kbr+zVxg98ytr2nzodpzCDQ2e6owBQw7ZU152OMdAcK8ZwZhLU6DBcd46qVynQHDnHTl
p09ITjz6IFBdajKm6MHFshtFVJ7FG2unLR+u8+7GHydUaD1BD7wlK1ozPNJg9whLVahnyMFxm+qZ
Qt47CHpqSk8XNCbVP8Dt9w53ZMcrwGfGYva5DKjOXObyzo9cOMe+N9uIudJG0Yp1oJRXRGjfb/VI
8f2U/UXjH3pR7Ox//RqWDY/VAb5gbma4YfLXWkQxxc4VS4l6RMooJvr3LuvyFVk/VHja1P+DasQo
r7k580Eh8tINgQpMN79wbRB/Y/XyQNIcME0CxHtz61TxedlGohoKPqxYQte5a/Z1b9AfSr7cbqqM
HdmTrQUjOqFdKwwVbB/7yBuIL1+uledz9cdDZCRJBOYEWlbin745g2d6wqRrdLftY3bFf0LSCMxR
RGUM1nT4xqx5n7niPns9/1YY9DTpXXGKx5pMz3vkas2Ep5n+WnqC+c0uA4Xr3NtIwIm2MRIh3MPU
3+DuB0edf7DwK9iK8fDyu9Gt5p+Ydld8TH8WfdYv/Pqq/Gi3ZMu8qZTLCDc8FTklC0wVcJz8GgtE
pxa0oIGKFQzk31Ztgs2EyS7ZVATh8oVHH2lpbjYIxLcv8xE7ytIDW2PFiUrz7elryY1ER3VxktJ1
fAg58T+QCpZrsLywCjzRBQ/oEyZrHK7qIYqdmWSGOuronFpY9oYR+8fUiGtNRNyRPOH/sdvXRfHT
QF5oeCEfu1gbIJvq6BF241iAY1r+cx63GxikiZ5gH8yvUOLlQT0C32NiO6HMmReDVNjxAOLujDBz
LZXE6T1vkQOMVmL5ttW7+hFJzcwpSOzkv4//bgQy6uuWCTU9RNyLlBkMZPJzAY8LeEGEg1sc5lik
0X4W03b7/aJ0bfOo+9CiQRO8HfniLFMsRrkdlFbR333nVa7/Ms+LBQp1aul/027sCfQl8ibW8ruN
Vk3p+IHDoM1N+NQvoAL8N4uAzsXy3xQ+2BQbK5qrvb1Fbes05dfZfNwCm75zXnNSNUmOaW7Tzqrx
lcDL8gnbOV09Z4d0NPF6JFycBSJho57NEquVaK+8EGdBAdnicO/RHpXGWNj8ru0V4WsddxVc8BmV
dq4FccwbfBTHlQHpp6J0v3PJrG9R6xbF8rlBdV7YmMCuQzy0Pqf2H+BmmcjKWYZPpYbqZverIbf/
NIM6IRe3Z9Pr1tjfA9KmLcHlpLobB2gQpV+YjoeHSDozezi890udJDXn2CHATZXG+GBubgPI66TA
72wwCdO2nXWyXlHzwP+INiDUxKXaM3V4ZdCs940f71d+sO6rnaV/etkDbBGNYoaJ1CO/v+3JHX61
vNpvYlGivzBpUuhLhI0MZMu7f7caqSmoEe2Nwe3y1LI3zOBPzEilFTa4SUsTILVveZjrCSWs9FdY
1laziNGJEzRvHYsvpYRcB95W4SZdaUsdaC7NDOE50odBXD6kBQa/rysCV2UIAk4tC63oAh8pKxKJ
ZNbEUTynm6uKkZMRLejbesLfWD4qMIILEMBAdTFrQdW9uyqSy51ZbtP2IZI4c4IqvBVsKyTUOIty
VpBYlKZGsLwfy3SL6ehDc303mrFNUBhQBD6QEpOjuVwoskNjpwEplZ7oOW/ygxIwKR8jG/vHWgrK
dN7Vw0puL0m0XVXB8nMr7hZqv1W2Y5z4tSw7GAXIQZDcj9s9Ft/Klg1fHBoXcZ0oas9GqQNyLI5j
UjPBo+EicpkLbTHGt2SAyuPmXknmMcV38feIVkOfqypcYPeic8O49xBzJqsDiFS9BI1awy+3I3VJ
kfgTS86p3t0jnHm42/ObVmjMMF2s5qPOQAr2k0dqubUm6J4EX0ydnLZX7wTxtvG7niZDSZ9CJ/E+
JA8sznqLtmbNtUSNR7ldQ7AfTgct0+QZQa+dwXkIwhUIjX3CyFbr5ObIelNoSoWh7do/4DdKseHW
1hiPrQX1PhzgxDqnL0dKuhA8oZdFfveW4BlZAPZaIwNLpWwWoGkW7BMjEj8tXp+Rm43xiBruJ98H
NlnOkhYx6sW4+T2WSe+DrwrMkekn+NV8R4l7Qn3PYSB+Nx7P66G1maITn1D6Z2jhY2Nf8M91zwGy
54puE8Qs9UMKQg+TSXLQg9E/9rv6J+5X7kQWVpcHzjDGbN8sPAoF5mgWnhog2D6fWzgjs5ufkjr+
S6hHlX+7YbLz+lTt9DPyb+IQZLgqjwig9Xku776Gdb9ZTbtHbP5b7Bp8EZTy1tvbiCbaxEiUXFyI
sQ7aQJXBfYIuIXLPtL+zZksrXN+RLlyOb3sp1/2YM8a7z8Kh2xOKuufdPfV3/tyDJ8Brt7pAvAKY
B3ZFkfVIClazJX+/7Wr0yb+J4l2S+BNl634WYboP0yOen5vAcfRQJLNnelz1O4b3UGxryCTPAPsZ
NS2wmvYiogaPpt3gvuRfNifDiTyD8GRdY6KbMCjOjaJT4al3o2FLv+rjQWuFFl9ng5h5FgCTFkU4
dxQFxzdA9xy7jM5wHXq7xCg7k0fe7gVvjJ9COElnXf4Gpj4sIEgB8TjsgeSFNbdBtevJWFyB15ac
bLBEGoLvGx/0nUoEiSWntid9la9EMW2FaZUVFo9SFBLd48JTgisprrQY4nE4NvNIv9UrEz47rDCM
u+DKmRhGb9PTTI9aQaboeJrHACS5vV//NpHGJHrmhb5TkMHD0IZCXM1ggMt5U7jfo7hOyCPGaR5B
epfstUKUSA9/MJdOmq9nVOcxj/G1vci2wtVSIz+kqyv79zd+CH1nRN6LZYO6TEMIfzh6QRdGIScl
Pc9vZuTpWxdbyGBhUQAcS67Srdc22WCHCeK5tH6527Y13TyhwPYcMA2gkHEcfdARR1xdd38wp3pN
tws+LxgG+Hub8sGp88jPOiQRhl9BVEo0S9YugaDOngDEj8zv9KYQmMpJhFQXpGIgIH2H55dZHQXQ
xhXj9Eq3/9oSrtCD5StdOBgloqtEXTBRtTTqe70ntt+V60xErD0QdOjA8nhj2ck8ZW2q83pCmWdu
OAkE0nYRKnL4zfU9h2XTEdxyq7P0mtXQ5U7EFAzyHYds3F24Ldd3lxS4OOMMi7QdkjJ/fWHD9Zua
6SJrVopiq7rfzPr/xQCrpx5uGy9IM1xjP9Z73CxaUB6dRlvmWKdJneiX+pkgMZTp//Zeg5akq8Dc
ygcBXgQH0FaKG31KFb8CcsnPLfTk8JiY06RVgdnl9i6DUR9X8uTqhnlCuw0GSDR6l845nb2V/QIx
IPSRB0gzQOFv3uzmVyUBYTbp0LJlKpUVhCbB/81bUStubO5XKzadWr+cm7JvJMcBrWokyLc/QTAi
CJWKiNiWXIiSUm0v3XnwkJ0/cEbqb9nRdk8S9oCsGt5JyWdBiSBiqBOQS+qYpBFXileP4pVute/l
85teVUp7tLkbTxYkwrFycgsCn7Csv23a+jcnguiDI70Ci8r5ntwv3WZau9xueguGHxpNa7gY2B8p
u4y9KtAQmPSB3d6mvTSPB+Mhtttzz++/2G4TqDCYFfyjuif85Tfai9f9GxVtn8bxtSWhta9c3bty
93K9IPsNgaqyJEvgilWSwlDtA/B1a4smD90gZ5+HGIXFaddE9dao1so59DU5qPYBENBJ0yXvEdZ2
CZ9L7w499aw68WZIfVB7vrxSVIslB+2ypgJ3g8jP68g7bLuY/k0Bq5UFw5VJ3CIcvXMSbpXiu+zX
7sOvbevpXo5b5nZIJ13mYjR2XS8oxLu33dWZTcJBu6BVuGPT8xjRp5f+X6lEWVGkfldw0d2Bs/tw
w0vDoHPGXP+F9Iyxj/NYdY4noQ2jrSSUJEV6XtsLll9NHj9v+guso2kqs00lQmFqBQqNybwhj0jx
vIbA+pYEbhTSC7fCmRlPl+xWTWPNMyaIEXn+Cg7AcQe9gCmfKq1zAxo0vTTTNThE9Y62ftPgdTSD
H10/4EqSbzqxWnHv/kZdcbdzmYJaEoiz0Za5LAcvwqbL35WoBhV/70AyN3GV9RXyfF8RYe/XyYzD
s+yFyf5BQssYuHyGPDBJhis1TbSDlxwHyadPjY0tTvuz65mfAXdkbKrjJGF8JbamZq5PByzDltkU
K50ZzTOH/Fxi5gMbkHbVYJXY8zfPrmaA5vzJIsCwM9OSr6NQLSspumYhVOpykSBwb2iDLAh2VObC
YRhqMXgSWftvdNSw24PPsdZHape+qPfKCOGPKA3layEmdhJa+FdsYMRb4GETfI+U15z7Rap82918
RFl8y2WnFpsAlya0tbiZxSg4QPi8qTGghuA/fBJdlNaNLjAdPVBYKgttcfPli88mjSKRLRuYck7f
Bu1cA0twhEOr4G367wd3/eWluDEBuO/hEu1rM80rsBdWvpRjC6xFVlxhLzyr6Y3ubco+2f3IpJf6
oVjDpiXsJeoa1WroOaVOU3gZWxbM2C+OiFDz6ol5WSeN7+XqySUFHUGrtNxHVnwl1WBPgQSfjc9g
o34K+w9b9lqiRUWuPwAqFjjULeI9tI13S1HcaiJrnz6pH2hekTft38ysHTukPoxGuXiSDqXPIDZ4
hMRKAKsgtCoYY40sgmNCFWkj8R7kaOz5p9Tv/W++wVgegvY8l4E9ew9uKb9LNJ2g8nmEE275x2lq
0CRbH8wd/DlItME5i35S56dtUHLM9f0u56je2elo4wHb+j9ssNB8NhDKfvBstvDwBeDvWq9e5/hR
8zU0gOTTt7kbd4xdzFUG4m7pwX0VlOGbL2UAQfNbsP9mYJxjblRj+juMVqO79XboF7Ou0QWBDA96
B10dWPo5QZNUnFWT88NqZUScvS35LRW2YWT+LNA1iClMUR8bFsDgSxChN8fn3Z/jQzV/h3l1q5DH
YdfCiLfOT5Kny003f7veanLjRsBYWzuPKcOUsFykmHmdN6eZh62jYufzkIzILUz3iHQ/EwislV+d
8zjPZTRd0MPGCbH73ZcTCbq8mFX7/b0ruw+YU+pGExsw1dPtsxb02Ar7DqFuw6Vml2ABqUnWIql0
TWbi+JS5EEp9OkzFWY621qDT1zxzDMIGYXD+YdTYaj5pj3Iho+DOYXCjGYxB1p5irNYhIfemTO79
VV7Ph6tDe/9msXElzBVH7UglJpMuNJLGEc1GNBOuZmhY5iwhh9e58cTc7WNr3U7Nu5ICNputq7eO
WXtTIjo0y7WJGE88h/XkZQCI5Dtdr9ffss/WxHpcHpvchWhSRjFKL/JsrOhSVfQ+uHUQYZIPTdsg
y72sj+WFbDYzQbDVC4WN1Zj9lbPGTovKv+bEzOaR0CpY8HlIwPvJOiBI7sGLmRGgxhDUogL9Z9dh
Lag67KwNGf3fq+F/Sq4MVtAckiThIryDkEHC9XBrvCly8qPod3Yb962iqXxRCSDoP3n5Fj1n1TZO
LrwJrAcF6Nu2L+GzcBvyY7/M0xuv0dhWOoYDkKnovSHiZKNFgUOzkEuhilIpzmzwdHaqYp6MCjx3
vJJV36LKPCFIOTDI38/Bx4udLTJRTE+T8SfWpDEdOzgkjRl1zOsdXWShgHIt9T7FQWUA9uqu0izT
wO35SuPXiBnoSTo5sxhj07W4OgRD+Tn69kHFczA8yiQAAi31sNYmBBy1RTiqDnG9Xq9672B0XfnL
LPHjGypakdUgXRasEvCiByBcpFn1pM3VXPCgVQaHrzvNXJhN9LOxjRBa57yA22HJ4G9S7EutxVtz
XTTJCXc5DJ6dPhMJHeRSy/meKlGEmg2N8xAWBtWZ9PULWRefRrvGFWat6XDVMvHGldxnG9elZ10o
AAwUP9RQ+I751WMSdXaTQzwNJBnwfBZ6YvT83d+yb2iqVWOZ0XcOU4u9tmD56o+sYooaur061CBz
MGc1MjwBL386+e7E978jpPzij6bNGwCcloRQ1y6vOFgT3s0mLHUKKrYqPqseSh098W0yY/K2cztP
+rG1EWuoXTVDv+Mz1vykdTzeMfsXzaJsQDaSwgQonc+4Q2kuD6czR+ITTjGne7RABqrt6c8xY7cV
rrqhECvCmbWJk/FPW0r93MikNuyuN5o7AX+sH871UmlXto3TmrG9LOrb3IKaO3gf6MRgs2zdHWzQ
xxkb48D/gA0RHwvsDe++fSAsrqs18+4NAxVNZskI1MIE96rVRYbcaJrHElutO2ryNWwaYRDApy/k
r1wA9wQgVhyD6VZrgXG5hASdxf2F+3+eFWyyfuIXx9hVUZcSWD5NjAzyGtEx8DqbrBcu6xYBnlWU
ZojjI6DRj+8tQlPL9oISdlWIKNhHUdFEllpoHEXBYQhzuwDksmE+LRN0WGiSf1A3/rcb0hjk+b56
QRi03R9dX+F4/8XD4LNJGRMXeqDpIfKe1p+lQgy5NmTjZzXenYpPd4HQiotlApdY3H9+hTR4hczu
kOjv0V4I6Lr6JpVkwlLUPDIXbKoggNYGTbgQO8I7ZeVM7qBfTBcHKqFkch83yUE4ul31iBCltrZr
R3oWDcq/vZ1lSNqipuRe8Hcxf0oyBpcTcdJJcqY1DQQ8/q5FalhYCTDOUPIatMIaoADJv679b7lG
Iv7ghbfqwBtRnTfaQqxElY5OUFnnoJ+ZNLyIvDQJZDqLGkNkxe890rPWi8Ntj4MqNFedJHzz/DiW
KCe9tAQTRtROMuMFBc+pOpheHJhFveeVrWfxVzrXao3Lb2adrKiQshmaKkPyGpGJtRVp6RcwxQtq
0qKz1hm+XAbw63Ygjwcw4AZc6bIrravRw2FfA6aybPw9INWi3tV3PFClsrQRx1SE6MJokN8YXC1N
F0KQou7JMDrtYmUBRRJzHRE7Hzyi6ytZHYPNiTTnzWMlavgegIILI0jc7cfMTso6kS469KB+Hq2p
AerVEJQo31QACYR43vCFBJGiqxA3CqbTv4VwqN+/FexweY9UA9FsR0OHEZ42/iePgG1OGD+4v7je
Wa0l23KOm7bwgVho1dVq/E2n8Mz95eIqGaq/ivUTFal+tR/gOvPr/tQcQY3pQns4ALuk9vDZp+57
JnIpdNPU2qNxgNvbd8hNr19ew2035rasEMffZw3uxOlCvNDNIbjbnRZ/MLMph3LGvQG0xDxFlT1C
+acXs/leo2hEdt4ukwz+AQxo8B0OdV9rGlsi8srMpZ74qrHDUUlogkZvqETyGrDud6otuT6CaNpl
m55Cv8WtQC0Rrwy9OuvSwIoPoUdAq6ZtjLug0JVfJiur4VJ3vbE8rgNRzH8cNZiKPOhtZoO8DxwA
7MVkI1y1emBsmjfSkoHodPvkvBAwCQ6kHAKRDOtQOJd7ZfHMygd2/2hSyner4A7q8c0OtrSeZhZG
z3iV89jlpC3uOp5CvFyMTAX4Z437ckieipV4SYGCy4y/qWhMI9seeuVTaeBalVI+9Xgl2CkBVjn8
uATvIJa9kdm6gSZhnwvTUnQfe1mp3CtoTJ9XlLvqgGOrXOxQ+hzved0X7evInnnKGlUBApZCh0oG
UCDRu2hVMW0QU8aQQlhXnZDA0Ep7jY2b5OX6JPO9wJEAg5inv4uyEYaLl6nd400D65vOqhBFAoZI
FlEotvde1XFxGZOddq6fdEbcwMonxUIoWg4LoP04OlLengFWjVF2+bnHM+QRSziWl3DKigBZx/Xp
as0tH+A0fTEjRGVw3vFBWuw+24WGPJV54N9Le5FbdN+7NnmdyI4EHzwxqM8BLDLgS8uuiYdTnaGD
6XyM/0BygsJ6vhF/AqwlFmZHgjOzkKgNE5hfceJTb5UtEHuSX5MMCHJNgQmwRc2gfKzVs0egu0f4
uexriw8ZlDjaAarHnJBZDAg3C8EHyul1As3mzB/5URM4wQPXtccbHEFqJf3WfNPLlFwyOA0DGFQ6
2hYtDQ32BmoSf/mFWLjoANKuAQlDbXYYqO76rUutjvfWOy2S9r02ZXfUIS3OzWKu7jlLjDmwZ4bg
BYqj6Dv4sAH0Dmi4Pq6wRJhoAh9XIcr6pNskK3BojCEmw/caXMWnyOoIe1Srn1bGhKUniPQaqW0J
VpZNUYM8qrDVBMGmCcGmhrBakHzvteKxrRkI/a/o2We/vuJ8d/kdfy5zuBGS0oOEGGDh6EJdS/rj
mDrICz+/eBtF2iODBFbsrFN50nxspBZDpCaW3dwLGDbIh09ZanmlwAGUqcXn0xupHewOFBCGn7eS
ffnVSovO4DFduFgqlBIewtZdFN4vjfodkfsqM4asvdR2RoxqaxKHySiaPptdF0SWDGq5SGhn2Git
odVTv+HD1dgQmW9KqzhHLFwa+aX+zBJfD9Zqw5kyn1r4E+uyulVe9YsRsZMiPgwtYzbL64QtHWgK
sJW2NMzPA8hMGOtDx5SPG4pSZWNml6vZhrfM+4ASkt2qMDk7uzNtNWmsFS2cFNkiQrs7pdU2rk3i
yZNEw+ob4Yt8Q02k1VZGhZDZ3zUxNoMKENtnpvwFBeGw6GYYyUkGE5czlrEl2t6doD72gurRcJLZ
uvxmzwHPRV3kDgqxA/3sEclTEstqCfDiTv5+wq05ITfY/OkaWn+sklFaw/p0CPECb3/fqN0kxEms
6IBLLuU4cBanicT3A5F0y5Og+q7Yz+jREZYvH0art/qSyzBIsxJGGSjh0ybVe0ypZTqmaprornzU
/01qO5FhERMcADzSTEbTDvSftlSp+jF5f4KKeSqLwnDeQlrBqJ2EACQ0jauUWydS3UBuij5xAhBQ
fA6Bu1kqiNT+HXIemzwUS92zPdTPAizSZ37Zbu/ZeEfmej3i8Wujxtk7akhSgODXZ+WberoRsJSr
N7v2f42IdzNaJlz5njhEFq5my0xzSc5I9gR0A9Fwx1S6LrpqgObs135wViBAt1zVlFUBC+Wr30Nx
ZlrWSurAKKrTzngorvOuEXljMaDOOksyjQY+r5kCo7YJtHBf0EuSJQ4PxL8DQb20hGCvI41ZFi5M
kLdatpHK4DDlelSPWZvN74apxv7Y4X2Gq4zkqRJ8yDgvA+pqdy9fCbdJrS1/q4C+22niuotqCond
ZLxo7DGlJMpFFSRzTAPdoJoSk6d+xn9C1a1KHFQYX/N/0W/votk9bu5ribj5wKK6s5abY7zi+2NE
i9XHsXx/0XLIsZePHbA3dGQj3mocHFPX8NLEMZX/aVUUhnxt9ZIEJ0DAyghFVoW/7auxdiXCPYTz
RWLvguC7M7XghARdcc7AkjgHstjAD5pH32SslIhVrWeL6+sEQ6IZz4FqDPvdJzAezG1lmtjQPehz
oUTnLdpOGFn2K5kHd+yLo5fW5zjXOM502yvdbEDlQKYiBeGpVG50BN7MA5vD7+Dp/ah+K2VPyTwN
7o7ybxMImHCbqpMK9En94ACclwiB4/z0DdKG6Xe1Jm0Uswxgs0gIGb2jnjIBe7m13AAF+SJs7nwz
oBkvjTUqWN4bjRf8P4pj2Rari5ibRFgUxj+TI5rtLQdaU+EK2wYFQwnvj68JICcJqCA8tCfjfgpT
sQ6riGvf8c7QJofGQ3S/YkriI8/pf3W3xGkMRk9a0W9Oi57VIqziujPTyinBadWJ2LxiA+zPdhSh
D66T/fqyJxKEa0R2JjDdPXKgTjIL5dgGy9sD+6JlHLvZ3zSyksxiWFK0V9Z1uxYSRQt/ewionPTb
GhQm7x3XmEdOzs11fJJQ4TdRbVW5L+J+JaW3/0Uq2e+JY2Sr0K8NP93ga6eLNO9ixX7JK1x3gmku
2AuHtpAh0rKUtJ65O72j6qbeJzu+DfkIpS+IzSEaMm5PY0bifesoxG+BOUg1bqVUE81HMsfx/C9A
bN6L8H26VGCW3iQeVaYcCNg3BxF9R3mYFcui3yzITDc2uzkcpy5IzC73Q5Q1hwMRU4zyjPbB0N4I
QAuHyrP7/E7j+t+DBaD7Bg6BWsefCQSsu52IjCyu2TTXO9s9+cnrdd32MqHYAtXHLk1z0k9GiI+n
IVtSU2fpHAGKXMY3V65Wj8Gtecq+DHwKl03Ev5kzgBQIPSUaWDW8NrLilo51sDtyGysiVY/K64P+
nkGrlJYBBDpSGHilz5pGt1qV/rxwnNHgaDEr5jpY/pVu3L0NHhP7Vp69Iiy19RLGx1T/crGfYT8j
qmyakurau/usLXu82NbZrsVN3q5mnaJwckrrnYwPmNj389zlbKg7eoMRFcZzB5eNT1FtOGzKtnxw
52AgW3HS8if6miZRqBa7g6xT/8m8gvHdoFzZ4CHRjoym0U4/IOVDm/9h8l9sqeiqcdny2YfzCtXg
DMCEhKAeZ1ob77RT6jiMrMfxriemDoBMwn4NrECD1I+K4vuHK0muWZm3d8JxtjI9mbwjxx0esy3s
rdtEJSZMajVqPNp67xC6vlh8ZrZZPPjseB9/3Kt+UIw06HMp+htOaWcxgg+qInGiRoMHsCTHx0oV
sPqu/z+eQ6rKxb4vOigoeupnhoUX3t/8olCyg8E0w6UgbQ8CAz5jXTYbwxNYr8JVocnlkLr4DWBo
uo2HpA+J0Ux9FZW9NwJAqDtJzeobot4oWuBDeF0ltQuDLB7kn0Y4GV6BHeGEJ9DUK6sueERJZHHE
mQLfq0Dhg/ncV0p6owAYmziN3/HCneN4/Yv3tgc5+BzX8yKc4GPsf0RLVG1f/G7lSyggFFnYlv39
s1Zo6nSM22SNb+JlYrWRV3xoawsF0JUEkKIG37Vcde4Y/8EKl32DLNk+okFvwvyx4zQBgAdD8fbb
DS2Omvjo7DLCdIJ8qwqh1U+CPmqGABg/B+iud/E9vQiB0TI5ZzgLvYFgBzPncSoWFThkkc6nI2yl
qVjZ2LEv417olhdMiCX3MsDo/J5wLdX8A/F/0rI6iq4rIfwYw1AYTrDL4ug3kc/dsAhakiqmELQx
ZmgrCwGEQKCAoGdWVQ5tgg0yjqLSb7tZVqcFzyU/8jNV03j0e3VinSWopPrRkWaXC7A4k1EH/+Tm
+Q4kLbuj+vYBoaM5Qk5bI7FkZW2QDHPjBLYHcI3KsRfZQz88VJcaZ2ddQkcPGn+vJ3ozSmrQKFll
jsMqWEVYej1Nn0jDllUrk7X5UqF4ui7wko1Rket/F3ryIj9lH1BKiVEATnrxNCWbv77LUfqD46mI
9x2+waDoLhmrmQeeOjDZE9VHOqSXOrAFLzT1ZKAFPONvIhnrSa7NijtlQlbF6aBOHG4oYb5VjlEO
DfvouBfwYu0cPWsCfFq1eM9wn6dYxyoN2oXY6jj3NwIUttiL6MzICuqNTlFpbjb47VQrDBN8c2Qn
O0roMf+rrP03KO8E3psMZJA91U8SoVbMcVOCXyAmb3ek9bbUFlSE01qFp/MpZusNB6DvnIAiZAD7
nGZJO/J4OL9QwwpNie+/4ewGkzhRpnfSDMQ2lUurGezxuwf6oCEmgmK3N7y79PJ4U309u+JQE19f
Guo60qKBgPc1pLd5u+AezjZnXZnLUZKfJ98yAMXPjTOB2ResfjzL9YB/oYZGZm6G20NodnGIJppa
UqRlajIs71tSTwNtQ5joB0LlDJcSZJpLNn6wq6h3pHZEOaWoLhQnRuoIDppxaQWEFTLHJ4muJdSX
/2ZZkBEYEmQjFG8Ho4ptsR24BWHIac+ZlbrKO7kMcBEe+JHmttGO3QPdKkQAqwo1VtWi3wRm4FVs
22TkOLtu8EKckk+J2fObkKaW+ltMiNedZWWNnk9ED2TK/Ze85e48SEjbfU0saJ4Qd38i3a8hPC7L
NUg7eiiH7CKLoK9sOK9kjVBrGtMto0U2vVAf68ew/dClBWytUWkdKgsp4SYO2gPqvCtd9AW81B/x
NGU7gUKWhefnk5jcXuq70Y1k2QYdnpzAs+Sefnsnm7z2nzmqN1YNbXxSZ2DrQK3LWMowsupStZlU
PR0o0L6d6Xu99ci4+uUzlaE55q3wNKrafDlgKu7wkFQgokwCc3CHkcfc1C+dK1ivOCL7S8lMjf7J
5wYt3opSz5SrYb4iyhfjV/6tX3gvV4eylajVpNXj5VRrBv6asehhBRiZzecmuyodrNxs+sDivx++
77GAks0Ns2uSF0X/J5FP5J0bTZzLUtUG6H0QZFU3bwvuD9s/qsqRrvIGdcf5wT/dm2nTP64v39qk
/KKxWP4NFmdPdsaXnUVlrOBsh8I/Q2K6P9J4/CUca2orzD53dGY5A6YeXe2yEGHcPAzkcxoi52ef
87SaH8l4/C/CjOMEoirmwyosX4SI6F/bSUdFQFUt9ja6foFfkc3G+oSXGQ1Q7g86twvvmN8LjxWS
W4FnfRUCRVGPVHdwWrsg0p7idImVJixzg/mC+S34PVJdD9y1tkDS6ltYHnLkyya9sMKLeX4rbwuz
lWlzwJn68H83BZwF18B7isp6+KReVaeTXMSxAAJQ7/sAuLcnOgf2VUbSXLjfevmy/CzMaGIf0VP9
T9xgVPYVjaiQKGQnlBuf9i3KKqDkBdkAxvbxyGHVvFDCCGx3UK/N1uVQ9y6kIv1LVFp8S1aZ+aRm
nGgIUGh0eRctK5WKrTLwY5X+kmKXwMFimk/BTAX3tdAOoGZl7ZW6Ys+6ydAyQeyu12VLfDd3pzjR
n+FnBvYU6+jvDF9EDY91oqICwnYVv6RxN0V+kBBsGcFOIg9JZH70OFozObKO8CcS+MZ1ZiHA5K+D
kkRUbwFOLpEiCNk/s9aEXSvtqtuIXVLKyDpNIus/6T1V/L9J4bZOSWrwiUY9een9gO7atruUH294
9jzYIhWmVEXZl8fvZZvlCU1K9Z80PTUKE2o2sYjnR24pksdN98M5zPpRs7w1CBz7aExKfXumVKwx
emF2lqAYfx4/yxSWZn77yBVBP+7hUrSCQ5hf69adEp7vJNNVw7OpsKdG8Chy7v5L+2RLF0RdWjdT
Ics1RpokiqKnRMaPB0s/+UINClrWCqarQXdSxdq31EVhfPEquPJyQfWW5UW0kgWdYIRwuxL/vVDG
ho0To1VqknQYzbdVurHkd1N1yoQz/o7bxMvMYnhhwtEXe25iUZ5KldCBr+a/7vZuuYANfaIo8jht
lNTlQlteeQtWRfIQySeI69VNyjJ1siDPZ2G7F8FVqDDkEQTNqqvF77lwu9N9JTel5rnFS6+0RnDC
RkffvyF7pSjpRIAbLupxzLEEqFmqKAAkF6062whtNLEP1+9CKj3v5QplXI+/41bHblbSnz56l9Kh
y+p4s2IHo7WtufxsS55KYFmcCOIG2EiSBkw/Kasmhs7gANZYNZ27rzrCAXDRjaSWnUUyvy0CpUYP
mWMheVQpkyPvCVM5YNDLNdpjlDibYyAEhCNuaQ/UPg8iU7xvBWej5qUMgL+YfuEThzSwefs/LhsG
mJDz+7D0vGl5iZ+32creW5WV+WQf+ksNTuGsdahwQ743Pa1sOmLTOK4EskWmWoXg0MAG2AKfFoWc
B+5EYIe6G85NRI0xdL1apfOB9MgF+ksslfugngHKyH/1rBKbhZzpbD57E+xUyPB2fT27vNt5TW0M
oKmKGXxPOgxrAqLXCbT4Nc0R+2ap17NHGfg0jr6jUu+yAOQilcecgsqPhTddj3f9PVIwHADG8pBu
7G4WAL5RoKhNRq+W/49bUGoxOXZR3EDaSGtxdXuxm7S6qyfXxYOQpKgcN90VXRXQ8WbTB5piVqS4
BEGUjxNhR5Rql8m4EJeUnM3HXsQ0pvyEWeOO7M8r+6MfNVc8fk/Aj/iABSTvPbrdaZOAvN+OH5Mj
I+OPOreWlji/aIDxOSha2eQGO/WxrpN4xiQqjkHbX2L47GbQzTfDfPQlNf4kdDubiBKADF2YWeSY
JBr7UgeZTk2g8PvLDVAyNqJdyYLpiz5C5ALlforFg0Ii/aHNofHyclSRU0xAquLm0gYVi6Tf4PFR
7f9s9tX5rc/tkMuKxKPzyFMDwE23f3CwO8oiB3Vy3rpdt3+j3sny9d65PKoik4/Jd5LgKiGD+JKG
JNpStgwiL7c0AstuLTHQxPRMYId+0uSRWzD4+DHSHNhNsvqzcKuPuwT0b+XGV8YLGm7eeVlFx2qu
iKCxw1THzF+xdE/9ePd36Xw3S4RngM1nhxBkuGWuoTXyi7vEC03J5oktZrdOQV8xwgpQ3TBOFOxg
QWKp7pbTxupArGf4V/xD6PtKjNRDJvrexMrJA3MlYXqEbndiue63WBO6ZAdqe/sKK7v7HxhiFoTH
fvsFecss7vEQle5lMRhNrVS/GpwxztvCrJF98ySWYq/wgrdwzcDU+aeFVMEput0rN2YFxguQAMSB
yunNbrFKZjac7iKLJZXT3xQQPByuzciF+8YAczZjqb8g9u4Ut/y5BhE3eotue7jiShPbE4J9mQYt
r92PxvXy7ugZL/KyXQGhsbrqgxTKyzV13BRgy/mqhvLzKXYhxfA9ryf1auJp2dc7Gkq+MqxaAp2C
Jg5+Z/NCjnaxCT9ljA9XSfpih1aGZfxMDcrwRvkiFLcLuHjV0NjTU+yc9qMMpJQi44uXly2cjR4b
3BVw8SsqyYdeb0vk0w6scYN1onwGwuQEBg16xl+UctHfmCsGDr7D1IrrzmPopkHfsb5AOE1o1XVs
R2+r14qg44q60qMTQPmRhe0Xy6EN/BQX3jHIkqGmeV2IJ4QHTb7vXorDNjI2Owzee6lxKxy6C+8L
BCov1BU2zFy/BnHoCkCqnvVfIxXk6igxH9b3VHpemNRYzwQqwI+S6Wyb45iAhjoPrEPoCuN6uQgJ
VHau62LeZbKIkdsEnY2H+7ImLl/DpsLLe58UH8MkGnOWBCOtguMw7J/jsxPgwb09mQfG2W0X3qn2
xNsj/Y5EPv1S8gbwVANsES/ENBKRjACu/v19kWMXBo5tVs5mbyHaKrj+7kPjst8TiT4t3UAIHuDE
j+B9m7BB89Q8IJFleZ7JXybmPWEabu2FAz+X1O9wb8B8LsHwBden5cIJLzoJnjk0o0xHoPWbbExD
SEEZf2O/3AbeK2yfKX3c2/QRZNYGBKjt8wZryHT1NgRc3tR/i6uooJfEhe/XfRiFirDvjnpyVX9o
Dujr1FHivx2dr1XwJeYO7mkvCY2P4EMN4b/cEopSgoqE+f4dnPEuoML0B56ncQkQlLSh1aSy/+WR
72XPNXD81plcrfYTkB6F1aVaulmJncgLdaRoQ4btL+dWrQtuCDFFOJeiygoCwPCAnmrBoL09klyf
TPEiKxHOsoPkFSWpGbrMdLFHGn5gl3F0sJcvF5qaNBih+zwsycnY/f6lsU/vrgBbssKtWY1KakPC
yDxAnJyZABujKu6XUyoZA3Uhnjmi4Gw0h3gPV3tdJHAcrCaLI3xnyuLeOokMNWX/NXIMNDmXIClH
Ms3Qyi2UtFICZzeBS7VIJRU1XiKJT0G24ETUQMs7cYS/n1W3Jk9wXESGlSFV950VyNiOGx3TmBzv
5kfLTDxYceqIPPY4/sTAlWu2D7mZYwlOiRhmhGDhEKDK3dmEemBE3UzbrIxR56LuDPeAea1dLaIV
VCwru+4B80xMe4fVjPh8sGEwuszll1LceBSAY5CU4XtZcozRXt7oWbJktCqWeIZX8PGr1mXLcNI2
OqX9ln4EUgRenkM77EeDX/hXEJd2pCVa4VcYRLgRx5UI4J5UmSr6X/WY9nGUONuC98IXx0bDQ/Pc
2ZcHUzM7H5Ks9uXRcfseBqyRDUPPdQLeeJX35pk/lgk8mTTelmlBny1IHZLsCdMSXrWOyT34ZTCC
bdz27BayUBmcd+wWfERWUOlpyEE0SOUGT4m1R/Hcle752wrtyOdy4TgqBxhS5TZt/6CG5b2BQdJZ
qDPIJUFf1n6+SoE1CFWW5wwiEh9EsYcelV+NIPliFzXiT9selrqU7R9dEY5kaAx2imESknnoatps
F22vK3nGnN4zdLITKZ1ETsTG3s+EuaQZJaRStn/p7StfNxgFOCSCkrYQh6jNGpVk0ckEu4MxBkS4
jT4IOWFwyst6VK7+fYJAsQFxeYiMKC4rGzpRE6+C5+lNsKo90LrcRddAiCeo+ZcB9kfWQGE+tV+k
tYMOTu4EsKDK0oZkXAjw0CluDFrgqMRB8UL5pzS1WVfUVhPX8d0j9D4+xR1UHpy7p8MDz+A54LgW
cpPi91Sl5zOqbtC8nu5VbmHRmTB+0aQj6iScJE8h7h7d/4N7GIm3wyYhIqjb/CHiIaZdujz9SiiX
rP9W06QidbbEMEmhI1Ky8ZjhL8WlaqqinbGmB0Uz+ckkTn2lCgXjSvYRI3/jro02eOTiHf9qKFgu
0PuhlfbPeuhaCOxZ2iEK6yqKdypQ63xXAt9FsUi8SbPj9n4Mb1ilO59V7E+rkU3usXh2Pz4Iz3PG
GkleFXnUPqbq8EdDdwGWn1rKg1wmf3PHKamOR4dSHaAnxNGzerzD6RL9PdR8tp2wlvSrMwB3XW5C
51r+jIUyHMItREG19HRZ4ZfwWpuKuWb9u7TwNvWxGmpjCzPs6H5BJGpW9OFM3jNB1Xb23Aw2gEQw
WXWuTn/sis/zNQ4PWxroqsrL3SFjEqmCKSB2Q/13lPK3YeAjrdFJb4XnE2LzM2fwMosCLxt42hkq
Ply5xy/tffscY6eBP5yQ2kvbsAsMRECo+MjaHtho/5Mn/0hz+jlnsaxNm7hyXn39x4R6BHfqPBJZ
g945+XKIGx7c0ESL2on4UC/lSxr9CzYHoWTjKpyiT2Sqo6W++f0rPxAFL2ZvkT9hFrdg+jd251LZ
FqzAquQgjbFiF5sR2WRV4sD+27C0sXgG/QtI+2b1RWu0EgYaT8L3S9jMNNdsBh+qpk+YJBlo8E6D
Pba7fOJDg1tuIJqX9RzbqFJK7rWrMzdqKcwIH0kzxj+Gh7KuNo78P1Skri73nWqXk+ae8K42f0ZN
J88t94hg0Trq6q/o16e3IHWn0Q8DYWKe88OSEfjMVdTZW6M2fVp5i389bNw3VGZmN2l0KwtknYsI
adcFyHzcY+8CsgVE5vw8XFqbxKPv0iN/Z3EKPiWlUM8ONHajpD/KPrnDwSPK0ULHH7xIsvxOMO9Q
JXnn4zWefNqqKRAcGoMmnSMtQ4sjURpnj1P90vhEZ6MJpCgkOXzbmZOj3UQ5KRtpoEZS87Sdc5ng
2kUOBnsD6OeuSl3tKtkqfoCylj8tc76/Ddyn6+plPIclm94lAiG5BapCoPRHPjVSkPP9hsFu3CD3
Z+yw624RQx7JxuIBK5tul/8KH8dK/dLFqdOTmjDW/zbaELOwNQxb0M0r1v9TjzYsQ+dXjRzoHL+p
SVsdjtIS2XVxMNSrTjZ29CI/rK3+RR1xDwLVvp9NqA0n5Y0pXg5uocLkU/Y6Od68y6fqpT2pbJzJ
QpfrpXWXyZuaHocP87pgh/Mvj0foSjbIJGtl03A5c7BOFvHpOww2aVdoM1hKsV8sMe2FagQPfGQ6
+QdGL+iL9pJcGMQJiicWoK6LBt7jYZ5r9lkouemAA8KeZ/Pk1dzaqpL+GGfj0poFXKX66bjHc3t9
oiOpwxrMKGzIEBLUqMozCkGx/75IwBf+8BnQDsOyEi3gvUjbdkQA033ChXRPplvEqMbAtuhPjMvP
QT8EYbpO+H4zReQesmTHGJ5ENlHw91PWk+rJJTYlti2U4Enc8Jbx6KZ+Z+E/yFDTPxmk/6x/jHf7
DlIxfQX3aaYjNrM0g/Pbj3WHZk27KPXvJX799l6gwMIlWrneX3KiuhuCq9ycf0hOriq6+ZazUwfL
3Ff0KqC8kHrktZ84eSUyvWc8CEyUrDEJ5KAazjI47bcb2vXz8WdrRqvd+aLNrHR6pYAug//tXp8d
95SDVSVClJ/yo06sm/jmAP1NZGoeAsnrncdMB9suHee+M3GApzhcegfeXR5K5N3Fe/BK+ak6W8Q7
/ZjQ9cH9D6h/hQrtiBZbqXgdemZjd+ABM5G+QLcKlTnxgb2eA63B8G1BedyiC/atEm+4G0XTY8T6
seiaxgbLNM/jhHyzm2e9Wf6SAxXb37xN5yMO2ICSvAFa9ijBqhNHRGO50VX6iY0dyusq9gjH/qWX
+DnhC4sBNe5h/IaOpVVJZGB2RZj7IHbKVRBmaVcvgCRe/lM3pe/OfyHMoZrN79pU30SEab15skVa
CAQR3k832D34ZmKCX3qpRiNUYXHUkOTOQJVi2HNObQi2WEei5+naDjYNHA0aWxCvmENl3ji1TGi9
myDlpT01qZenzZJCvlip4COXf5Ltb4ZLD36XI/JKuXjy4bZK7dy3/zQbpEyORqVaas4FQgnyeIX+
5MFnIIZzHyNwpPp1nsLA4SHU4K++jadYlw1XVu9gqGNbkepQ5hA4TXs4jPRJPNDb7gQS+VMejIM8
R8CBrsyxF7Ff6FHxOS2MwDlkiDviI/ITLtfiO7L52e6IWyFYIOQlSSx6LIWDa2e4yLK1D+e8NIpM
rrm2bMLkbPostuchqJhyGJSdTZL/oNRck42/2WmxxbGIoLvO5hSs3RSif9jwVimcUnlUW0sFnxEd
TjdWAblxvBYc+gSV9FoY/y/qUeNNJ527H97JIyZsE8Y1mrf8Pa7ZrAD3f0LJuadQoDlj74w1qwlK
9HQl5f2lz5p52i3VGrU7p36646958N9am8n/Ar+i1LJVRjEAOM5sT8isI2TEZDuijlayTaaIfnCb
s4SYxJO/cMJZFxK8Y37akrfj91bxFdB99UXrxGsryrFir2UXwQojnRFwQlQFyMEQpv2gIwFSM1Xn
4y0OJoSs/WxUEe2gqRfTHoBN2RLftiNCjoRV6dL8DDGjBXWjcpDIVAQs2FfXNjL/RjI4iE/iA2g9
qvBA+SRRZewDI4+VDYWvBWbp4znpPCrwhzTCBDLZP0NpzC8hv+Wa/eAsGBRGOyLvRRSHdjxDxODe
u/aLZE4TGhnENe9qX053/2VhLPd7pbpZYqHNFysitc+uQjSucKnQjynCwyipPL2koPZyyuKYekOT
HwO8RfEoS3OvZt2zxgjx7CmMZRGX0S5BQ8u9xL69OdkmXE8dSr1e92OcrFfzgkFewe7rl87KY9sK
tug+x8C696ZbC9Mp7O6+6w+W8eRhe1PF+QdZIXW71pK7YYhZyXobFVP3QO5Wdh8ykwWd6XEHVPki
5AbZD8c0Z9+tgm4lk14TGkIBn88H2MkBvA9FKnYRUzJeQANVZ61Y9BX7yS5bRqlSLB74IXeo2+Ig
/BptjWJdtenLINevtp7IRp+MpsbPTZX51eBdV8sW6c7Dep9vNd0fYEQO78R5vtqoVNgYsFz4PbYp
6pbmzKSd+IbWfklwaHZt0SiFfX4zNN11181F+97Tx4UT26XpA/cOe3IEJ+K7TnsO+aQ8+htlKQmt
xTJqvEzs/ve5ieHQNPTMgF9wOyD5oNbOOtvaxaggtsuCm6OJ0NVNIgfImmCTJ5tBe76kiadtxgOY
UMVQKVTuArtp7CHPHJgkRfHS/WmsSkPPb+irrIy7JKvySSfjoBzT4NLheR2miPVxYsQwhF6AB1pF
cQZxoY/V8owx+U7ImOMfa22vNIzG0/CQG4AKePtDK4SJ5VYcMn4VVqtlyV4I5FV4YOd7sE+vmYCW
lOverniMlOkyOkQ5xaWw2ZHw19UNUCgRSuu80UwOeJvyTq6YrXA57C4jdVNZBe/twKzDtB3u5ZDa
/Mu2IV6SM4fRfTqGgxW/TDSXrbZC2Hegf0Bjyzsbduo9ohxUDxo7hKNE0+YF2gF94y0QXFh+icgi
r5OWUhwwLsAW3a4eEEKiTmIXAqjgQSlKhBFzDcK4Yw4MHSX0yDSLhjWSCabK5uINxjMH3BCmrTiA
kFaLAMl0QEl3HvOF70zzp2x7uHj7O2iGatkf22zalEHtPkZavULm9v/9IVyaurUEUzbpyqa86E0Y
objh9opsX4nfiZxZTFVZcRJ8yv0OaXr374rIAjZju8SLkRNT0cMTP30IcomiJh1IvSu54aowxKmQ
1p3R9HVfiE9rKgoV0+AYe8s6tEXH8wHc8GxUF8tFBq+j94Jpu+CaUcoXxYTNx8QBGJuKNXc/NIIM
BV+dIH6VjK8AKCb3zWZx35kte2U+ymr8C1Srnovov0ymwxIYyEoJsDO+WLrDJxCgr+FJM4WLPxmh
LJl1LyMlTom63TkJ1/ZTuof4JIyyEE3WtS/8grmrVVoilkf/xmz4BzYRjOR909859t+4WQoZ5vsc
QP1/eAxdvLCOL57NSNTJ35cWsK7rIwsLMGHSpqdnuFu1tPwfS4GwmHS66dux3+scRlX/Bkz0zQoV
yjEE6NODJrzntPkL6ZxbqejE8wCJO62s5y6dsiKN6PJ0iL209VMV+Gif6UcLiJR3sZlIWHtbW17I
GfFJ2RRK6tinS1OtecjPFaqmv5TC9bG1XBFMu91vglH2xPer2QnWYaHTL1bNreXmGiW9XUu2cv2/
I/QfH4c3PepGIUTIdFqYzDxMqpLYAKvsFdlgpG6xPWtnyDsNlMQ73V7aP8FgtaYlWvb7Ph3sJ01g
fxxuSdP4uEmp+zaVr3+tJn9f3Uso544jbK9Gr6qE9LjezRFT8hr8fw9aVlO2ho+YDYWIGG581GFq
mnRKL2eJIePrNTAGJc7xSFrQIz2vJgBPXuZZNu3kc9ZcTUVgFYN4iUrZSpQUOhZRWbWL/plAuwhi
EQVq58Op9TOXsONig7XdPaNgWvqWk3g19NE1wORAb4CPXeph8RhO2DZYW1F1Dh3UrC82eNg+1L2S
u0DeJK45CxYr0fNEAMmcEJsYNLPOLQnT8B2aZD63Hjg0pf9dwFt2j/6ndzqUvNkJ8Lrnc4/J+tyJ
9LYHumyemOev1l4gJcKCNmobMipjXl+0IvLP48LdHlSVCqTSzgbKcl/q3g3D7QWqtnF7xhd/Hs7Y
EbKBHG+X2rVDtqwppFCmdhWZtuXHT77zSeyPt4r30eYTzH/UYNRriIFIab9tfcJWmmVTZQN7bBXp
7abGsJ6amdfNozJMcrphmDEntvWjn0f8DKEZ3dfF4flO1MmZdILNqZhQDZVeuPka4x18xWiHk+s1
ZlyiVwTaynA0rOOtHOHv9pp9nGeiZ+zmyAmIShQyUBD8+G7x7BICQN/bFLTuXRvO68UeU+4WGO0r
uf5gkaLeRhLWuzXDvlMjulDs7Sc/erdQG/2/hqf0ba1aZCZ2KLG2JVkzEKOXErMcCqhFN5Smylgz
lYqOY21bInsJU1GiKgNrQDbNFfyhgGHYR3ZpASn9L5HHq+qJAQPH9QORDA15RnY5jsytXeCBhxXw
Eq6eLhPAJ3q48Axtz5MYF8HcoLU+t0XEHgzrKhOudo1gOees71uadEm84fwzdHYwRQWhcMKhVaTu
N7plCGGMgUUkpqbPGrsJRY3Fitasudxp2TIkPDOLXeNFhpkrv9G68+r+rqBX2vRSfCtGm8t/b0bT
wZVoiiI2sOU8ZFp0wseWxXb4xXOKhMtHYtGyX1MKLKpuWdATiT1Or2lU9BdtvU0u8BV/Fyz02EhK
gk77Sua1oeU91DUFgmP1FUnoIUkhVNuNMr/CsQ/HZH5ExUQ4v6Ns0opF1DyK5nTjjuZu6D3kG+F2
tf4OWnGQ1PsRqT1YzXR7/Ciqm1MMmIS77J/aFwueNMyuymIVRRR6BGr110NvS0qfgwa755qxQLwG
0Tdbp233blMiarg6xkzYpBBwUEoUPSS9h/xXsIuTUN+Pw5egl4XVRhkSXJVSJomtncuSIKmibg2f
L0zY+zNkx1/L+oQNMgas6s14dzOdCteokNttJIjyD0z7MuYKk1QzhIcRnivEg4hokPnC+b10gPHJ
zUEiKXPxZYc5lNXyKGTGEqtLD5zDViuMZMl8zVg5aEqWXKBGQbqqp1kkVS9yMUmo6mWiIig2hd8n
E67Qhz4z/7OvxefyPQz3cedAfPm2bzR/bkhbV6xzmXapn/O3Yn8qmXElNLwfRR43uqhtKpFDUhH0
Hp8jT98SeHotfjkHdtmHQoaE883NVRxVKjPkvWm2ZynvbmVGQGJVKVg2AvJAHvVSS1xuyqdUBtuG
aDOJuDuCEF/cUuGQGoOpfsbL+O0bOnjNN3Xr+6G/ndfqxldPS1Xlg3ko/PWHy70utRk+I5V7gG7d
cO3nnfI0eocRJhbkFyLSbpctBcM33thFMoHSMaM4Qsnmh0gYOMNj+qUMVvZTJ8T01M0ASKNlaBq7
Yw3Ia3CIXkL+Vkbpdx0yTNyJE/BP2BKh4lgBTb//5O+X1Nb9dbqST8PmE8oPnZKiPAkxGVi0w8Am
sCmervyHyrwPqJ5VTli+LpEPahlbcGTEgMt8YMj2p75Eo85YNrNSaA6PCYcPaayXH2Y2Yadm09ZW
rMESGh/6a9j8eEv9L77UIdPA86yeiFIeKW8IglAJVLi41xObe+vlzWfPau/M2dabG1t5y7VF9CDU
065YXI91KY+G9rMOkcxBguRANgVU+nZydNqQnKdOTNIHqR95CKsR/twAZpymMbQWkfs9WFKhDlLX
8KWmIuL/tZ1dm+0gBojZcBxSNqJ6umTNmsXX1JkpF+dcYKEsf5VULBKBXFkWRdxwlg+uOmVQlpT8
6UbZtwXUcSnhGUTktjx820pdTh4CfyuZ3+XycFzwTosCRk7FMhmmOz6dbBZrlhCAIXjBcn5uoA+y
l9TfHXIdXXP/qRw60xO/SPGpiCAT3GT0vrgjMOxf/P4O+gsQjXh+CeaSRYjeLkadD5aEsAQykSLk
7TPzg0SFa0yuqCd9Fo2ZzdshzkupwFG+0+c9B+YkcbZi1TrVqHk9mxzlY+xIfr4Onqqv3fp2b04I
pHdM0Sx5dwHAucCUWKC7gyln2GmNwR7Yl5JEKFtKF0p4uGVgmU6rzRlA6DGfroIQvmrBkViJ62K6
9KmRNQo7Ph6924utWORHUstjKz39+7RluBkc5dMf7oQIyOVJbJbU3cfvIiOcyeFQyDAq+mXXQ2zH
j9+UFMSI28w2xcpXx1/CdQIDBewOQe+LAA+OK3TTkut/imgdnKprHAcyLYo7+muUpd4aGkWL0Vzy
enfdZVM3/Qovbqa+8HgIeC+uRr3e7Nk9Qb4irIiVH8tbrA47UKhDZyURZEuu3DjRofMhLw4y6lTq
Y3QMxSSj5b9d0de4yzmWRC2YRXh2LYbmymAFJ/Y+9psoLI/fjg6Y1Iv9EJN/kgK4CtwM+GWq2G2g
W3jRQOGpRGba6EwYVSQ38X52zK9GD7B0pXvo4Nch2cTdB5vXN4tiF0hRb6wef/pyxiVzzigKLoUn
TEjve2sLmPSS+3D8mWnLZAo8JDUi6nmBSW3qtPr7E/+utH9K9CNgP8R2eHZPU1wjsjh76iuVA+Ql
Z096elewcXlNdBD4hNU2MaKELJYYwF8AC6LRmOzQoXsa3B0RtEtqmNAmbSeC3U/8krmmIpg+ivdb
Tfds9pl62gufmIXJ9zKpBG6zfLBVZ010VvDQIP2dOD7MpFR+xpB9/WXHkLyyDk5/YasJkOoTA2LI
HnE7O1amevfDnxQsVtzYPoUyu7zwhd9zopf3B+RB0ARMa5vXVkGGMx3jem+Ri4oMbnhjrPUv4P5A
+T6XntwMFXmSWkT2kc8c5tneTaFs6ELqMb45y5ULHCdAG3jiqG0qW1ERK6+dgBBJAQy4DY4xwHqI
fYir4wVWehPqOKVYpdSIl7hZNHRVgI3iZqdigxBNr7XQVqSYLpMVFgxPlnB/5pqk21PVjOfLiSxB
E+qT/3i/cUWr9EvdKs5rbwwXS2nRao1aeJeHHaaE/uQ/MOZZdmJ645NlR3GDkogTTf+rz+uOCoCC
mg3QHiFdg4Mp5F2rCOAfONAYzPqROI1WmvU3hO96xWjfyo46dVgzVkMHD7PV9v9jAsoc0um9eapX
kfgntg47BPMk8BhWA3YSOKK8HjK+7L8MTaUlH+A6wcaA0kLFWeMBT0KkY1Bjry4hImMN3uak0RbD
i9aOjbBgPwki6QMfiRHYJRjEhF19YPPNb2ad9vUyCuTWlI000SVIQv0cqpjp8hrODvzYmbG/R4ke
q+r040ghTGoF3HNelLejYBFvbrwnf1BqNRYjrdIjRIViy2jtmGgqc+amNw4CEdFqPRoGO4vHd0cm
6nKm3ODqt/SEuK85lGqVbRbMbfTsIIVobiEd4/nRNPrsE82MMqYadp0YKpjlMoNXhkIZWO9ZLkYk
uTm1wZANcEvOGRQPP6/mC6r6vxyWt6OtC3DnEIeBl++DO5EaKk1sjsKsvQxQPbBDOv3soTklQPHH
vGYT6r5B4JlfnCY+2O1rj9bOmVnzoVhzoew9rHtICTgYl/HRgSNjmKXEbyeVygFqXbWX0wgMP7IO
z4cXVJ4oVqtyRsChNmg4t6VH4CtwBNTNEYw9kDsUtAkJc3CpiLPrXsVxxqjLVQ9V4WBUZHOp0Asm
x+uiRErMYgEL/vi5vd1477sAydMKKKiSGLNV1LDuz+BcSJwqwpfQvOp+jsOT2GOupbEJoj9v/caq
Tpqb5cqYm5ZrDli3986cavSucTS3zoObxrdgSGn7f1seTSAMUVH7vjam82qKzuRLF8rBnBSGRQBu
rIDuwsdBVYTlSrkaIXA7Gi4/jsEevTruxFdyjiMow02RTlk6RJEmOIvD3KdmFFkZq3tirmF8qo1W
fHtqcQsOBu6Y47ltocPG4aCLDMUBGOfXoms/YmocbE7Icokc7fBSTcPiuMMTnSdPWQjgWHWz8uxX
Wfe48jyIQSCrdvJMHVtgJ7p9FM0KQWjmpcfJbwnyaahG4NtymsQ/qm/878eLly2aUQAikKO8HsSQ
vmi54C3NtQ2lmmTrgYgKHRqvw69uyGEbUOqYn9VB4sNQB61Pb3G56PZL1IubQNyRkKQ4ZckrlVxY
orGAk80Zsnlhs3AGpYL4mrJXs6UfPvV+2Hl7ZJqf74y+iy+DjH/QxJayRi2YIZ2VZg1l8yeLOK9R
2eFhAJrqq0pnKgnuZ35vKZMRlQHDuR6WmAKALLqiSXUtCqeZ9g5NnpDOMqiwvY1YuaUBV4rLxUyM
PqdvbXOGgJBbGqlQE0qTnWsTUCSwG5piNOKywrLNp07XlC0LrwS7zZrvvWe1AYDU2d1ExLXjJLAU
PvKp3yukBjUwZ0BhLXZSBTNxuDMnQGeCvNahUVKp95N4AE7KErdGidhycQrKTFELG67dYRYbWZUs
EMPOc7WrMkaWj04BkqjFagIh8zAb/Yvb8QibGRonmysazv6Xho9yvVF9D2u+TwQnr5rMNo1wqBzZ
Ooj5vqlF2rjo4XjYylBUAPyJF0RNa70twijE0lZyoHz4jqikAnsogzIeT0qKITSE8Ly60PQt6AgK
dQ3JGTcriRcg76GC5kgXdywAZKfknoACnrZJ2/50sv8+jraMmtMg7klotckvLpXkgFP0KGKKzyn8
wzbKzv9AC8Jq3ZqonNnne+RWR/oAEM9ssCkxy1+MnzddY8RGpWozeoMHdrvXNAuLhrZ4e4yP1MNY
JHuoIS1pw4BbSxWrI4KKIFm+B1foisOk0WKUNjzl+NAf/F5OSLuFIZr1otUVKaNoBAxRXJy/bxbJ
+cZwoH26lR2C1VGiIZIKbF3Yi13ogcXHhk4hbeXC1bd/oVzXAm8/yUwLlmuDruZ4OOzr/ecAHil6
9nMvRehzTmHrdKX7vNnBIaNT10Ojyfj6ymRrTCMj8h6ibwFL5lCMFbN4hQL5lqNPw/a883HtsxCD
Dp0a3wCfwnvwgi5mlOXjoLI7HMHVE2A9s91qGXL/yQxZSRL7i5pirPySbzqR6RxNjq0eoSKwjPm8
cfJq//JiyYRRW/xEGQbUV3iWOEbafV7/U/BLPu7F4r3OWbuabLotyIX3CvAgY/2TQFPGZLWq3HSO
j12Dz/9ZjIvPVTQC2e9fG8PQcgmLej/9Ej6kooHBB54HYCqah4iOQ46afCkqwqVpB1MnI5Gc2prN
+dtH1po+HELz3yJH/clDS39CEKRofxzSaLYN3FktbdKJMCVPkA09uH5NMhY74c9W0qzduaD/KQrk
2Eb0Jp1XyrEPq7GVFiFONpsQjECn0pikUxUzYrOVz/+rOHgVjbgIZiWkN5xKaekksYTlT+iscTEX
ImTEDrY4UndE9x5eUjFWReigwuD/UdLzRVlWEkCMX4NIeaLhwVZdhMfFKWBwFcGT6qmvUpaLvQSE
+plFm9exHdOireNO6qZiuY3F9s94F2SfckG9ZxBtIOC1EVRMODIxUDxsVb9XBEbzZjx+Za7F4zHG
8XmPvPrPorTpvaUTe5M172CsucU/P8q+KNptZ16/vWv/AYHBFky1Wnu2tSNQR8tMVvlP8YfN6mhM
ShjVKjthml5t7/qutI4MIO7QDet2dUTI+ul/PYquPKl1MA8uqcq/e8lbKjSP4BGJnF/VmrCiB9la
Go4La2fNp5wLUETTzoYph5Vp5kzY6VkcQoWKtm8CABSZk1H/oSx5biVJd+YWEgSM3QvNkpk+SWJO
9LuBJRo+y79LBsdvoT+iDf65158/suThIClyZbv2x2ZNzrePIMS3Y3PsENfqyPscAA6eMuvntRir
9aUF3UBRzse79rGPpaBieqZorzdfCQRl1lIe8fWSeZK+OOQE2POMd7bbOJ3Mb0MKCbGxBzW45UMf
GNyPxjYaGON25yetntI14UiB5E6WCJOFJmy2nPaqIviyBYyLkeI+EYN5xDCJqZBLdfu7QMv1JeKZ
78RGL0h3CI1SUBiPPi57DIX4Fxg54qyDHW+DdeYInnmMHlhAAWZtF65sWWqzADbVU7eKqN4xkn79
9vbQ7c8Owy0guVt8jbPoapc+CZBFNE77ERLt0atkD+nNajDvfDr2rvCRTVNpOyOSkaDq7h5VRIgl
LSKhSxfyeJVHwEPkXboMeyjLQE7JUm0mW0lw/xDbE/by5/MUl6zrb3fqpR8Nsv+dxYT+B773Z6YU
jWYtnP2/g/llIG6wtEUobAYkdhUJBPDVurvjJNEkSHsC7X8/E0JdkNGaKLzsBVwughvW/P/k8J0l
3Nao6BhnE87ol5WnRJXlJFwwFifi7hOxtxKco2kPbIefxobSHFQ02+5PS2m3oQnfVqkrPd5051ax
Dw1CInlplSTrPtn3GPoPUg2mP3F6blL+fy+uHkXRrhsgrjKTn4Bu0kfrZyg3ZmTa4Un3h4pbUXY+
AFhOzJbUfQal5FoucMJHpDIQe1dZ9sD3BWYFMAYJOp3ptqTZYq2XBC9iRir0FgRufyVr+d0qjv8J
CK3NcIyaCovxo/83sgzdzzsSBSWiYYuFDsmif0GpJSKaLh3uFSGTmSJ3CN0V1iqUDKDYRxKo8MuF
qR4NVYyH5yblJRHBsBeaxm74htlBxPP42lXYn2RxAlhttqVTgzJo90lKss1AYjyPah9iCbMAgYVK
2zWybrqBHk+T+JR7gweaGEuq5TtVQJzifEuvlV5TjRo1Z/CqiyaE+iERNMGJEGj2gM/p718Z3BRO
AFkSt12fWS/tziK6KACLYtEU0O8izr20tY2cZLxvl1l4OFNMN49ipML1XxxSI/l87tAaCtrIul7x
v9hA83O43WLWWCQE22Qv8qEoU5rRzyEykXa1f4rws3v1DtnDPLZGoT1E43ouB4o5ELj6JT0AWqV1
n1OaH20cb4Jf5gbh0BVOrBfYfo0DWrRgSQ8uHUrwbTNYZ1mgF4oQNN7RN7Ya6jD3vXwwkSjtekU3
zZEDZW8/uvuGCwpdIOyI5TVS5D7AMq0hNXlIYnGDNaX/T4tBSZbj7u1qBjeUghyCQbrWm0XNSjxG
R6vJlyS5ynS5r7Uf2RejIAFTGDGiPtsBAACNq8aCORttGwRbHJnOxv87o1hhu+QyGoa7Dj6h7Ld9
cLQMZSyB/Ldh8PVam67lYTEiBqX5AW4v68DYUFzorOKa1pBGacjZCs861FKmlAHsEe27jje9800h
jjW1BwU9Ip/z7q2xKRpjA9rGz+7I1B8XLJXrR5pLPIW3+IGwz7ygA0vaPzmfhDrWEEWzHADGoFBp
aV5Idqmnti0MJ/RYVazUVFP8+R0DF1mw1g+jIBk7fb661mDP4YN/mfoptP7wOXEHqPmw4DB0Zz9Z
1T1eqn6s1Voxpz+V/Qjsdm/MbSNdPg4UOje0IeygTXoTBKaLtYTQ1AyzkWshhwXPPlrgOSeE6P12
aUgYFQH/na9q28QJNIart7nGrsrbpHNmhOOkdu/q1y/kSBkoKIfaFPaFWEKzVUWAOG3yjoxW138b
tEUFWrNDTJsLJcJHZwIr3C2zon5TKKwcMznpO2yb2mnA1yY2zbpcFG6mHLNbL3RJrNqC56inB7Ji
dOLFSOHhM98LH/BtsHYvexgkzEj4Lonsa9p6wWXZGf6tAJxbFCh0zwjxd5WuYz3arExnlnO6I/VW
MSjvQmW6r0+1UCBzcBSXbo97HBkDm1foFqSyVGsVGvYQI+sntEpuu6LuaFY1rdy/43ZSg7OqpTQi
Aab/Mw/K3I+Rau/5gk8CePF4fGFpKMVg3KomTQbk+AelpmT52u60pNIZQwRxlrvKIrX4lF1F7INh
fqKVNUIF+7VE7tnuFZfLIi2PKXSvJz6E9RnAP3XKrw31p/meKhmOVgpt1CzOaW7axD73hlV4MURr
XUqVCP5oNR8F0xZpgGZxYmLjxjZi4Hf4jn03bYbmtdbW8segkvOlwalhbFoRv2eWXGtgOctCZQD1
aNX0tnDmskiOqHS769SWxzuaManYoBkOw11neFuySa9esXF5+zUHNTKMQybCwYHO8iHjiiR7Tffb
g80CuV6+qJ1CB6R1O44axL1zyRjjgKE+dZAETYH0s8OKrwv9r06Au6X2f8IEqd2fp8nYxQhVD2YQ
V0FwFgMMMnquCEL7ad/3VLtPIvm+eCsE50GhfpGje3mtTlaHE0QXvs0Zr4clFXMd/rg+/ffKG2vo
6UU59v2zBYpYC8fMrQnQY0B4Mk29QlEHT3yah9CuOTwmYQM6fx0YZg+xXcQMfWYXsSJ3ynnpK1Q/
oHJTfSXAW4P+kp3dZtHJjHVltSg5a7Gfk2DdBf829sTBgAL3U0h85I7TYYFUvTpD5t7thbQbThpt
mTbGZP7v/XlJYuD2c4cMQyhioVhlh+qNIMVtEu02G30iZGLsPqHjAVvdRqROIblnwAuQDWQvIIUI
SJuFI6xvuDNxLuXFCOlrikdG47EEP8ueUeeS/bVQg6fMAJDHTZ593kfA2hlY+e/wiPLMeL9z3TWl
oD8V38S9Rb7dr9McNgjlz2P0m3ZUvMGXBR986vE0ZtwmRte3b/xZHxNqBsp9sJfM9RInj3jSzvj+
SZNqHc+wW6uUXMUGyO2TDLqzcaIu/fZxSTCW3BRaJdPkhaqX4Zw6qxS4iUDnGSj9JCsnyOpF7Yut
sjQ6WuPN9l6n6uKh5m5MozWGhsmToQUMy3jJfxiAlAla+pdwt75ckKjRuhWPjPC0qqV431us5FJZ
CtqFbonVDPLuQcNrn+pUoAlOQe66pDU3Q8+dN6J5OtjT/K5lKXJIGrJsLshRS6K0CkG474IOsQgx
Fb7GsMSpJUposmwX4MvAqNxvaVog4TN7TUrEQOMdbHlyj0U9shemAtI7Q8ShAcDjpu9Ve1fu4GFm
ZthnMhFFemeDbuhWonnvCGKR/HHpUNoPhiaXiCrniAbDGN4VuQDGnW84xOZ0n0ECI+OhCXVdOkn6
coMKby5Vv62AXu/TurHAKoKGJkA9SWxQhKjurP4CBhk+XrCUPCbbPHA0lUTpeu3Sr2keZvzkkwWS
wwQ3fnZUSUTw0p9DfBjNbLbk91Sf6BJcgay640vBFvzIENz32urOW/C2YS6g1KIOmvlbcY4kA3UL
z42MCxDnr0jRi83HB9qiYzJhE3A96Uih3zAW2hpXZdRqN3RQxh6gz6hAdNJGGExxLSy8x3UETfH4
R84hJgA3AMYdTKy7BXudG6Xx9rtO8kQb46eBIN8YhHD2usFStdsjrHUTxQCq72vM1RuR3bbMQHxT
oNUZ3k4yW9Ol0fCEnog7kd91Hiamw7gKYZ+oSNZuTjBBlTv8DQWwbIjv+BjW0Im5Uk9jE6/kgPS7
xVIJgS/JjaSBwDntxpNxnb1I2gEVaY5vProMrkgImN92+q0Q9lAh2+DaefrPjNkZQEpm3pMhMyby
gRkZqt39lFpqx53xgn3sdwXPb1XZPUFZ5YvXOwViSW7U7drP9/hudncTyUMHI8lAE/xnFWfVjF/M
YON22OUSJYweNy/t1T1m7eHMHUE+wXCilg5UYeqBYxGcNlJfDO48xrSa3a/glPUZO1wF8WK1ccnS
4UgK0csbG3li/smGKsoFYuXzodTJGfei7vAAttLIQMunI46MDiDaab6KLAObKTKqR14paUscwUsS
BC4zquNXZEykmkmzSwt0TNMkYjcPcE0tzC+tKflp0PwwYSKPakGlZidZCM15h1hJ/7QLHNEcUgW4
KkS0TQdoTncsQqT6EUvDqcVDDwRuuQOYMWMv98GIYzSyhfzSvOXU2FeFIww2i4rmpKsvzD/GC5Oz
9G2tOWy0F9mHkbPR4HsSrPWmuwVuQ1WAiJFweOo8xepP3tfnstv0MrkaQPbLHbyCc8hyeOSj5wyq
geguJQ9PfIOw1R8rWod/bHxzE9jQEFn8g1N+4u+UW2sso6fSu8Zn1NrBnaMvJ14LS+u/PMyMelya
6m6fKh7QRY2kpZb2rCanK2PS7jyEKsuJTaHvsuBlPKeBW08MeRwXKqBdsTKmK3loqbaF0gJQvevd
f97tOLsHqLk4yVq3aWYd6MstosRrGzH3neMZxm6VYzapFp3qNEHMpVJTLgAoOQHiYj2SBZw89cv6
7/vLiJG1c+6KoUcq0bo/m22/2QTM6/pFfoYsRE1IqSUnezBP4yMHxyTYvoXwGZg4AN+MF7/0nS/p
aBuF5pnGiGjNRGXxcgLCxsQDH/Ly9g7Els0KIC9lr9huSf4LzVIFw59XhpQrimifVzs06P2gIKOg
RtfWp/4MI1wMqXw3maiQgKaqh2JnWCm5NDqnqa3YH7d0TX1m9772xgcoAqadAEvAiefkAaTgxNO5
AxAjmO6WDZGdotN2ynENdG9ad1w4Zo1XOPODPGiuUpcNjcTHIIRFlbJiDCGR+GYaEda8WJW41+xr
QDegItQ8RAJWqqzw+cJxy6eGE0zkNILCuF/ArmQtpSvym2Xjm10ekh2get3XMvC0/E7c4z44TS2r
K1PJl3Bsz2d/I2MSkV/UAvCSdugKtdW7+F0Vjv9B0Gt2cd1KkI7eiPZAOxQMnWQ0eKnh1b3zIbfY
k4/OEPmFJ9iSOAcI6/mHX6uEceaWX/VzBajKQU0/HSg8TyjIrRNc7JdGVFYwzbQzWRQexfQjE8Vz
dwFzE0T+v5cyCiUojvwLyafzOpHVSNT6ZkA/6qLl2qoKE5Sr4uf80d62pmNiGkuJ8+jwR0JOXJxq
lR9ne9YpYIUp8Jn9KrKeCoBCmMe99troj6kiYkYaAKEOPAr5fxbDI9tvH3qZlaCcEsdRkGpGvOUk
hUBvveGCrIYeHLdkGTvID9vpURYgDksNPCT811iKloBgcWLH09gZ4nxGmJViecZrDZbBmQOT0rKC
92OtRHg+IuAYG0q0ud21j6HmVFLfWDPoHNi6aJgYsNkxccZSjibfW8W+1BCOYOiYuqhq+H+PkVWF
DKyzXEW6eIUkAxQUpTDA0KkYc7jIwcTk9KxMpL9ZbfPpAlJ14cWZ7vrENx+Jjd8O1qEG6aBiWDdT
ZBap6IRnjjCihW/grezxUQm1mB+mkBlpzNTh7wYVjbkEfxG+R8EA3bpOO219slGFeYO1Fu/Pu4nQ
Oj4h7Ji8HT2QM9Co4dsa82X4JKaYlmGy13GqVdzozxOe7nR5tg3pIbcUp26g80jL8lp+oAXmOO99
lyV+crdn84YS60XD2ff1RDzxVh1pW0fF2Sr8a7dBhDsDeJNyQWaRWQgIbMvxtGKNG4Ty8VYlktlQ
yZrqrQECDKBRJbNLySQnLTI9Jrnip+9KfYauO3S+JWyPg+gUX1omKm4K4mTPlh1OTxLvsFP34me2
dC38IDBIwfLGc82PwSIU9TvpdB5zScvVqoKBYMmZPWSHG75t+XAzrJrb2J9Mt98DcTAxxfxvTgkh
V690SxJT4YOB1CMJm6FPYtCdrXKmy3JjTmoky5pMnd/dQUY7fPCRKL6c+URys+3s+qtJrjBsAY2F
AE/AoFMMvrkwrlUsJajOxwU7pVkRv+uVV0q8virg+bAwjbV8FrWSvPBUFoEnzphE+ZS0rEikbw/g
MuCmwYZmht1Rkfu/iEzhzd2NWFMbK5EeTQH2ZPGHPsOql0bFXGwElE7ztK+qu/daqNirENBb8t11
e80dB7uAFG7iSBmBRrNxd+0Fd/9o8AHPiyHKpyR2GlRsaNrlQlWIyGX+qMnV39mzh2plMs2UzmU4
ma4ehplbqV5sCv7/D2p4YK4ODlrlRTglXMoLX3bGDc8+DIfFnt4T8r3IqhRpxZRRTVFjHRNuHh5w
a4IcgG+W+h2brA1eNBeStdpYGqXubtcs1dmr1jichjUxaf9eTG6muyMOwNuH2MNf6keN8FLbX0m3
9YOcupW/PPFo0E5vvmZ1iCoUDAYcZWtHIM0QEosH5n0K1BC/NekbJ8lvRg8NaztpP9LjA/Xm+y9+
F6z0FM6kpPJ5d8Vc0Ni5Os5F+51wAAX5139Dyb7A6XaMd6dJLCEkEekpeH1Yv0jBrLacaFjbtr8z
WE4LHUfeAMNEo/GDQpZyFLdScJYBoEbpDJWgJ9gKrPyrFvU/cZ+gVwQyyqZuMrJj2FIV/WWyA9b4
X3n0+I2Kzmi6VNPQzWD+er1rseJpZHMkrHwlA6gH1xzDSF+uHizS2+lwLSEsacu2P0qeL3la7K4m
5PuUVvTWVpBay80aGv1czGix3zalCTajF8+8YCZEY3WRCGmeO1V8AXx1UxMNjHobQW5uZT+DSWJA
P7TtbT46GpX9VIeuar9UifsCgnEtadf2MKL4FTVdIYHh4lbWJcFHRXjv/8MCdUCsFnivNvlJ/Q6G
WPQ5MN2XdK1vtFWJklf6iXNiVwoM4lt33ICntHqBm0e6kGEOLkN2l/zC8j0nA74wlIo/G1TN48Ei
tPgyE8SQbLDm7DDFzh9fa3HsVvJa2fRcqOurRX4PLF0mnwWJFPemDeNZ4jiIIeSn1cpFjG2tjA8u
VpSL4ozAZDErcPLtyeA3MPg/LsJLAx5I8TxQPGo5m4QT55jdaD0aUEdx3RIkyTHGuhe2Sn8ZIjRH
ZE0vL68fOVEghdmhV86THeYKKaFIuG2C+UCSv3RshRnJI+vMPTIdCHACW8wtep38Ahp3KphlJrap
p8VbxxfNXF4fiCQwuJ7LjA+Fgv+NNdYICDrVBL1YVIgovMd2z65mPubjWp99CWU5ftP/lkT7KjE5
SF2kcGYCnsEgFNngD2Uxdx/neAknS0tM2hJn5IdKejEo9cN0XdMG8VI+KcLcCg6BAv3HRFAr/FJ1
w+wzFqKDuUP7WnEiBIkRXqxaf3mcfgQMWZWyYHmcEQoj9Bxgrix0YMWpQfPhoCFurNVjYigHL6gd
UFK4T34G+0tbsvV0KObphnM3fRJGyKOizjgilmp9Jt0lGAo4jgSRximqeCLgHSYvXyfAPbXuldGj
Etkn9dd8gDOENXTiIm0b/ddEOVQxH7R6qeVyjVZWpNOQ7LUIApTwc7Te+MpIBkMwlQW4MG4Yit5b
3ONsZvaQbcoAy/VnWiksV8VtrJOPcbfU2P4c5IXIdQDs8SYGEAhPMnMcQ9KWVBFgM5rBuk6rxE2d
9qGc96Cywl/4nqsyPMINHvEAToaVAd7+FXL3G0lDbdmp4td4TGGCkA1QXMGVfU+ssSXCXseA3wDZ
pvTCO/tfdayqQyNnjVzkSGx8puvQOg9kt6HqB8tyMHWYni9r9G4h1wlrxJnPsjvi/5PRIUJ/zNOe
Ey+ygYlvvVjuBaTCL7gNzRxxxTKsuEVLfUHmlEk0OUoUM9DEY1WTQeYDa/V22xO+E6pqvgSLIGPt
KajrcgmQvrJwy5cs+sAB9ZBXwUw9bS54GE6zNK0WxFg4qApYGUtUysnMR2kIS0VIre77snvCa/7w
p+FdAy5FBU7JwjvBhlSRU87+tjeJLtNqclN+Tc9VmgkIU5EbZK1Bo1JRplaJOj0uiCtGUlKcIqyu
JSNtcYUdoOm8Ekbm2ZgmUbRDuOqDBIUNx18z69OSy/F6BDDqhXa6eZg+LstUkdI8Xp2Tr4jRhQZH
21oL28E0LoyA7s76ugOUBUHDVHtPxSKShYGh9Q6/M0ZwXVkF2PwrofRvXdniXQ1LeJTkZx3+EYLg
vlVhXY4N7W5UbO0DKQbP+sG9Iweptf0O052i+kH44pg5Cpk+tNbOqwvFSBS/GfnSItulg9fIjUax
RlfVEX3y2LTDIzO8V4IzUJzKleqY4Roq/zSGPAiWRdEnzd9KoBNuHclMubpfEKMwxMmSz7yBSK6I
miq1ymSZWK8zgRehONljicdEcDoniyBoSSFdLjL+c7fDOMgoYTZjdTxiNlV7MvNUCSZnrzcx8n/+
XJycbpdGlZUZc25BejFUOIWXgHTxVk8QBqpj9DX1rR6oh05c/mK05QfnA9/l79Ne80HHtzw9dgzv
1t30fX8EQ0f6XbjfHYrOS2nLKeBAYmUhYaABJT+O+zpwPsCTdyKNwMFhm6K3JVlQbyzZAakzBiSw
kzNLslOZMhsbU2EEq12HURfHoD/iN4eCQbry0BX/HXVz4f3N0eVrDqO9KExfjDf7UkmOH3fzaFjk
DgpfwHmvlVdWhs3W0UQ2frACwI4GyOPK4GcpDCpDnvnVke4df79J7ti/UxtNYbHGYDgFc1yKbhQ1
FDMsTd4DETWwHq+OrihufpaECR48YWwfwl0h9lLPqnhwbXkOzhLqAVmmg2nkPhyl28PgyAW09C5C
r/k+DaBPxpuX4JR3Te5a7+FZiCNW7zumvLEIU7WePCX/+jk+kN+IrAx9bdWbYGPgm1AhLUTUgG+z
Lh/2ey0zRd0ygbdC49NKb2Ybn0Gb5FOmG3opXf+mNWFl8GoQtFwk7IV6rBWg5U4Hx9AK7oa8eeVT
lDNG9FRBURsjUVfyNmME/fH9WC6rUdUEEY1/B7wC5yDsf7i94FcQn6gxkzFjK+NLVV4KHuKv+88L
qW/8LtYdDiZoqxHLufMZiKybZ+APSB2E1CmZMgUu/DvkzXK9NC415It4MSKzuxD6oC21xmdk8w9O
gIOljOM89PXVXtbbj1jtpllKHglZIZOe3pzvwCDUiHL2Tlq9pDbj6+DT2I9wgVMxFP+uFXVet48z
xBHXrxN3SrE4YTF+jVbqWRudsttiYMNoCzWKUbEHkGG4WZub7XA01rYtr7LQ4q6jrYMnnvkv+WI1
7LhKGq1yTAvE71qZ6TV7Opl68VcV8V1keKOqUVyeiuIOUJR5h1H7YwgL9eoBzCX8Riiju1cQOO+L
W6NH4UPeu7yTQ7zen/J0CZi5f9MlA26CMJo2VgRw4lFA/jvPst5+sQGBZBhT01dGpR+67gu5enA1
U68ZxuSNXwV9VpwXshhyiJ42FcLheHg5xEbLLN6S1QaDl2LA9QNz+lKfArcCDCjCrVRSYGXuHoWq
USIP4hLCw5bS7lMTWTev7yjFo1U3aeJM2UZ157lLiLXpD8FHmfBGumGBpmzsWma0befEydHAiDQr
1Oivk6yAVA+qgzRk4DgV8j8fXGmxg+6f005vvQJG6MQWRYR0XHY7G+RhQM4KeU2djsvY9Ygek3mW
FKvbEkWEz+V/fPw7seE/vb04AezWOwf4400+78cxBL3bzNQZkZ1/5eZLn4N1/dz1RZByIh5yuy5/
0HGj0czqwDGZl/UAlFtLlrRv5DcieAxOD5tlGA6oJXKtY+RvSan3XtpsZ6i5zFqvlMZCDDQ2TutT
6iHxdrzb8PC4dKHXP+Ue8+U0R6tf/r+foV4IplwyTLXkeywAoBKUGApeUX+wZzyxezMI156Z6pb3
m1DmCwEQhHyZ8gGuNsPzTIoBDdgAJr9LUaTxMjZazhdzHB7KJmTxv/QM+TRh1Yah1wqovzHx43o0
vMGxGPNPxwbSaG3ZiHGAHUuMkYRQuznkmcX2I5E32FXMoLfBM3oFoAh4sZFCikJOi4ho4gmxXo0i
cA9C1ZvcPqpGo/ZO2H9mNu2TijQwzr+jlvX8qowHZbeRhLug1CYE5L86jGHUG7RqjC2B2wGLJ+Qb
v/WA8lrwoItRU62wLsZlF6I+ivgo6XXev40iD1dP3oEUZ34widJZTx1lK7ube/fC3jfQrbnVb7Hj
y1cblGbK0ro/yq/CQz9vNpv4wNvwxNQcDfB5AXAehy/xTuBDF3nzVmlaVbSm2G9ZiTH23zGVv0S3
73QwtfI3R9i2E58rrmSRcy+BOYhU7w3302FgFs45z7xxJiOf+2snxo7sFqli9C1LreOnn12SGIrA
pR80sFcwLXfL/OM7NF+w3Ps6MtJnfF0EXT3fFg4qZHQXcIIakprSJnLU6GXRhLbREuJySPO00zgW
cPD6Ruelbzi1XCNUzbSbKwNG+D5Mq3zMaZ6Jjtm/ShRmmCzKcGguUhtynduZ+roVKOFiyUkQEv0X
46sIi+uONF1KhCMa4PtPP3FLJVN7cJ5bQ/XezBhq4477Ipc35kkHzDYpAPE7tmJeQMMtvMiU5S5F
5I65gYTl8TlsEP3VoNc7AGgcvvSLdpnRHC455ovoT79+piGbQCxcz5F7LoyDyOo9+CiJwrxhtPNl
K0fmmRajzsmRcKFb0URZ86wNzi9WUJZt+AbAOG5oHVAHwgs35Ap3sTB2Z8+wtjgDNJJ4LCZQ9RIS
NJo4EX0LvATMGVLnl0LNAqkvEmUNQxi3AoF/tZiJnyne0Uo4VyTPdRlYoJ4TZ1jSxz7hj+hmuy8I
4ZoKo8PRMVjTTRHB8zrNuY0z5s4DWJJ9GDfUe+QspeoEOIdJsi4R4/QRHVjQ+PM74C3EFfNkhKFr
taIgtA7xdjkkiaoxR/azeH9wMf6eqQk4tz0nwa/7Gf+9OpIDqpDoPeeIVs0XzNzSDl5L2+KNW7KU
JkQ7ihCKMSr1viWsmfP5Y3CpjloDYl+oQvoxiGjRdpyYlFlpg+9MxwEHXHvENs4d+gNEST4EUXAx
zLfX9MrVzORi5mv2e2zk3A7PLidzAfkHpf/vCG+fjalivPDnbLWJYswvVzdxBduzZaUMCn+KH33T
4kBOQ9GfvoyjFxt5d5KAEDOEjesX2NueGXjEib76u+ZMLENNKpuvVwKgc6HOnoJZP4XvK0Ko1jr7
XjvZRqz+3HDR+eJS4EXUYJdAYCHPABW7j4Q7exumLWjf4GFkyPy5KAXWjUlTDnBtc+qqtTKSXpqU
m4ZoP74+qJoB73qRivVsT95xcd9+JNZFZbHpchjiaOaFuggpFQJB99yJRB2i/M/TF2cmMz/nu9yd
np1IDjhpCyk57oNrEdhtO2WvAuBmaE1NRtTSW26/A4LMwMjQwQwkSVuEkN/eMMdr6so8k1dYKtXm
AQaRffjnQ5F1pKk8c2ZpvHoeJQrkTxe8AfORn390lEWspkoezIc4eSVnHT3pyQB8RlDR5vyFjvKc
UMDKvkrJpu/xU5xhyFpiVT00haK2VAnsUin9gaaFHryN/nAmia9GxdrP6Q1J80fkedZzdvQCV3za
NnWzae9En7y7SBZeujaN7Q///gnb9PTcQpdc5CIOLAm0Wrnem/bO07KWuWoExKPql/nWE2qARvfQ
veUVp5ThHQFvX8HHplL83J7a6ydammkaiUtSv9RZj4JH7a0n2QGQeo0PuD36r7JgNjQSohwxg5dn
ngn7he2ffSrobujYam2AWzCK+YIXSPa9cGXVPpwm9pAS7wDR/4XURa7Q0pcFbK6C0Ua8vRNmRoEe
Dq52DiNnwv6jUBytRyPpBhvdetU/KQ1K9+p4/lz4XMfidCfpGG3F0qBKcp23aIE58M6feiygIdvx
i3hCrldombn28h+MMsPXbrhJKh/ghyf6pkKARrhlKCHithQ83kJ8CR4UPIU7wBE1OLoR1XIc8Drl
cQ1GvtMHQukvi1vXtlLt88PAMuofTh9Zw1e4jZvwazSoqNjFXb+hjYw17odPrQSNgJuSJCidARQC
h2OIACzQ24OVq8TzUWKdixNnL99gfqywam1XAZsF68TxyvHd1rYvf/VpAfSiVs7RrchOlYUCZtBo
kTQ5iwRfT0y8NpgL/+W5PcDp3lSJAw3G0ij5u36q9cNZyIuureLIq11p+XKrpRcm8eMAQjVACDRM
PunTe7yBsHoevnSYW81sndefuSRe7cUvRHjw0pGxSHsTN6Gji/vzdsPpFGCuuWYIjHDUNvom38yq
7WY3eU6Z4iAHA/+Hjk53FAdDoB8wrbVLvUHBokZsw5SBzW/qdGWptvFUgsVGGAjNyD3I6vWcAkao
OxTe1VMpTO6HQtudW0Y/+PsA0+uihLZdRQ+CcIgOULx8ZQt4uMbZTz9CZ73tuXczE9aE/oMY2sYW
M/Fz5t53SU46qtCCZk+17kiopr6X5CAxvo6J63KXsh3WeJuEAGoLiS5F10dn1uoo3jAs1MtPLV7f
bO/UOhwmcWQ2IbmLr5aRu77MVwh7+hjBdzDAZkgrMNDA8HiCTpN77DpoykK6gHuHPEjX8etZRXKH
KiGmdEObtBkZ66pnBFNqelwhKfQejSuvIK0gSyGhggq7N1L3FiTnypa90gSAWfmiD6iu1VoRMM4o
12wUFRrOEzRpx8U1VGUKi0yntBam8DAfkPzcH7s0ceOtT7AKT0cgTJmvsxtNFvEbpfXhDO9VnGSG
o35F+n3b9TCwaNzL5uh8QILk8gIiByT8N40UQF3xkJ+sNv6lxsLCnzJjAM6L747iROm3Cn6OWPBO
259Era9KTtbMOlt2WLBSNT6aSraNIaSPs/lKa1+in6KM4PvHBGWS0+BNT/sjFL4fCe4YJEpFWOeG
nWNW8A4qUUCblmTdG67lSpIKEmrqsVL3PksZ07L4Vbhw0CFHooLw6feLlf7Zr/H3VFP0iM0gXiTV
mremATYoHbJpuryY0RwxfEWPJwiJBvx0u825gUcvqoANKuZxdm4t9ECl81K3YnPALvs7nrNgG5OF
LfOI4Ud5odzLAmvD/5ltYotZP0E7Cw87c/iAaZEgZEJiPHG8o9ZFj2tP+HyYyx6tAvim5s728Zhx
QajkmA0NVwWQrZ3JzOFqw7q3TGViW203m8hK71Bg40hl0XG4EibbuRsETuhoLS7a6RwL6AA//qVB
vaIow+zP9rSJXpxENIfZfHU5FuQ/7i5vjrhCsTIRx7kC44AudHoON47r2XjZ3uzIRu+NNVqCMlyM
PtwVBkuM4su7B9QJA1vdEETlpAtkSLAtoV5ITp2zbbgdh6iJjOT1ns5H5Nc93gXDXxeirJh6Iauf
ankO8XFldtTfUbKvxx9/lPZL30tWJ2Rwe6DiNSBLFsXjzttylUZYroSdoG4J3jlFLJvXEEJocZFb
0PdoBw1yqQhPYiXfVABmLz/SKagaWHajbFdhNJ7i7SoJtdhojYe7ME/u/UrZsP79XBQlmVF5yTzS
cmh/nAZnxHYZSDhYLqE8S4M80b1IWckeGgYlEg0Ti28cuSzOzCJLG8lRXnqgarYJtRhADGWs4sR7
NPvCx8KUizB/XfP+NHd8OG5J7v4dEmAS8oq4Q4ZZy/I7+nhN787XTMOI1i/qpA8K7WVpkqrnjnbT
kRKtkL/Wa1ufC/e9v8pwXBlfzGgIjRAtw0ZPSX9Rz+MR3HmjsNf/kM7b5l61X7SecMtsPCmkav1J
7NBB/KZngmHfCsjBcXaHcNgJ1Wwgpv9eCwo/qL41wB3JzYFvnqTGD0OdRASx49bKlwgUFzkGxenA
0+6cor6Ad/GZ5LX3ZZFJ5cKfDTpNeaGF3JdyECTXf/BwYidsuetWNaMTWUItrK8uh2uhunpHpkCg
qb1ThkMziSMc/A6DMzabdgNDco22iISKu1fA2ZJ5+aBlY7L1XnUUb2BBHZoC6J9pfTVms0lXmL0N
q73vYcbb0LDYYW7Le4tUr7ev9wv/nEwy7dcUO35QLNeNNvqf4IBusB4vZIORi9A36CcausyPo6dr
xemAaZH6a5KziYMh0RbF3nIanreiUBCRbQ2bhpGQusFSaFQVk2mw7RdsZfpSyKa9iV0GI6DE8Wb9
q2WvpoZgvyR0MAkf3cUmdZqfYQM/AOM1BuN4yCszFv0BEElqc7bnTktfWpGDSjtsRLgl08E3mO9n
5ZlaoNZBu9+YSa4k5RWiDVoWc33dSf89x/2OmOEcmzJAFR2KjMdJF1MEOrQTkTseSBlNCIc0gSmp
KY0wUoj2Fw1k/IuFYb2wCn7i2yo9DeVssXwakDI9atoXnejwkliimm4RCMisyS6i3V5QmdE/lNMv
sOmrBBri75/oadjOXSvnEJn4JCxx/cn4xD8GDNHMVK4OGBMyUY9ruihS8Bt1SQtN4Ml8edVMIoEn
QDf+Sa3OVejA0df6Y1TGuhwOUCpP0O7gQlNFVVJiS9iqmtDVLX5vgYVSFb1beOA5qiFt7teK9vRN
QCNUu+iI/wdrZMLeb3z2VHaoFlLAcmoASt4D2Nl0wtn2OcYSTSYMVuNpU1zxD+g89oxYVmakpVbd
J2SFZtQB7y36N7jqVUy7WghNIdKLeiaKdFoF7sseZjy4n6NYwxGQGminbKDLPhRyj6dePIwHw9bk
VOXr/HGROiKrZZzmNHv3CRpIHo3ookwdldg1vuQE+FQDkERN55cJP9bgpkIzcZO2CwB/RBIyhNGW
qbTqtiuG9ql+PuyPzkigPTJO7I6/uRYAUL5NEgnP9vDzBIc/Okr/c81aIaI9knka8yOF78k9veyP
bKkURo2T+84SyfqbEgdqAFoNj6q6sGWPH1xOjSAe8LeE4ZJG5WaOCER/t05ymUQDj/JgY/lJF77i
uEB2Mx+0InTfTL3Z9fAkSwa+kLRVu2zCUA1OdVTnE62+VCpkAyaq0GAWXxU5OkmX7vwxSXmx0/Uk
me3KHGFoxj23gromTRyog7GT5Ej3W2U1YpMlyXWWknHDYNlXp3tvbisBwEtY5hnTaSqReIcnMWcg
XiKSsxjnyb1OLAgUtIhm1OWsWaSS7FhU4MzdK3zLWkjOxOG7x9ae0f57lWhB+l2Df6/PREsLA2jX
yUWelWTcMjSVxgqURBsenzLsy2CzOgNHwurRoDK8EwDsbukQ3c5o3Nbo/MYRblp75SCMFuTI36WJ
TR5q1y4XwT9cXZoMCmugYKVNupnGHnsQM/bsl/P0LyxClTqduClyeGlnNQcxPMMPgzi8Q+fztNr5
TXAfmJSUmtxUvbKaLFzLv71kz2kuUqADQC5OWxeLzAnXLgFpNTnMI53C/zPicwgw7yipzhqX7nwj
HcWOQvzFdDeHHMuLtbVwfqlYMIJqdWYn0R91tcohGP9mwt5h1NYa3fYEa+hSVKYDLLlnxkwSc2jC
I4LqxkRYiA8VvUnrZYjbrGTXfV+i3hQQBBYR5DyLjHOO4GE0pyQQZIXjzRc6ptnog2KtDCFckFXS
3UcTX9aOLzdsSTNVQ9IEZ5bEYjJSO/C4wnY5nHEanH+bk1sItcWjb55PkcQ2eqBqczGuuSAQXk5c
5y2PdDgZAxOtnEV/ghvKEZU/S7fb+BomzxmAVT5z9F8JwLqMlEE1pMSzaaysPXdUxvEDJV4ZnLcT
NPBw4lp2+uPdmWZ816LstS/D/I+XAqIRI6wZDPl532Ee0CsJYp4KO8YuahU/XjulnJ4zFjwFipxl
ZyPV4PsK1WZfZl4raIDFe/QGMbIW5HbmBEjWG95mVTaehiyU+OH0pOu0cKWMPa8uUjZwpov96qZ2
Xb1pDNlkm5bdUlTFkHwmBLuOEFQnXAKLQop645gn5SRiFNoEOGQR+9lcsIQGIIks14j0pNiCAzuh
QnpbjvhfQcRkMkr4PWhWU8UX/gm8UjULjbVhznDdN4pA242Wzmk/uHGalg8oPlHamwq4+f6o4OeS
WX4wABkqTyZDD4Uluw01fE5mjl2UnoTTHI3uXBBz+iaQqKleSgpsEp2OgGnhWevEcXAd9txeamvk
XqvMlQRqHLJFZqiekcpN5a3xoWo02D/Wv0eVx0nkEo5MJvO+P7FtMDqQjLu16cSm7EOuGjrzae8B
/D/KeK/0X+DdVxjP4JDsc49Kr7gkc0Xg7JQc5KaJUVB3jc14W4+48Ud57gTVh41nWtl7d4empBdO
F2pm7Ea5N5qwB0rGEFvVxjPbgE7LdIEBzSwU3FelN851HSEARTKS9lJORqNlk5CUxdXLnNUiJoXr
sYBd8WFEfrhdx4j8/3mCT/V5pF9BQm0D4NOwRQ8ltmUil3aPR+s7Rsh/zZgOQh7VYPtAtWtWTiL8
H3/Jqy50iI4iHCWE79kNzghkxkdXzr0HKmwTQUy1WAU6Lu0anxh+U0OwwTdOSyk0//bczdHb58wA
Zq2SGhf9smzM+XuLqN7Oa//7XlJzxvcyvRWLJ/1wI1hc37uxJcOd88cckWnpihJl2jVHP6qtgZmw
I730t5l4GaJ4jmh5ZnY+JsDpxOqp9iSBO2IF1nxfDAcpD4tfBq16OUxqiJXhgR7e6ZIV7isjaE8i
CPZDTRfBFQUvfEJsSU7d+P6MR2GfoefdaS9qaAu6VXoG2yo+8Zta7jDzSKGApsGS8Yau3CQ//BCH
DmNSk9bLI74BmBofF3t/09W5U2/bOaQ6xLTgNGzFq4bdNbEclu5xVhyLfMnyp4l1an7OOoD/T3BU
ZL29yhmHCckv+l5vIBvH7jI1dOsCjCV4fR+hnmy71Vgbx9cQTTNAPjUwG0A5Px9GDLo0AUK5byuh
VQq+FDtbjQ1QP/jcQob5FF2HZ0nJDSxuXyDkeM3QaQeJ8wQJtaj22UO6hQh4xQtOhbQOha14vjb4
FlZzZlQD0KRiay3Cz0k0dgTeV87pYo97njHo/3tud1Cw1MqSHNhjQJqnUeoaStoNlH9sPt94iDxU
N3JBc4IpnfJrIjRdG7otAGnKSStkxkVj1gtFHheHY+66deg9aBwE06c4+7cY27lA1N7TZ2xGssx4
Gjx4Z2WNiAjrK7iNOFdPMXYdGMEDohp/KQWSRfo18yldAUqfeoRZpZXtOeUPDGg0BsA18FFU7Lb7
d4eLgNr0B7XEadsR/KaMcY7quU/GO4kaonkh6cL4TzlG41LpMdZdHvSHH6paH8sCloDvlLchJD39
eAodCTDNDKBq97YPZe84+8wRp45RB27rM9A+d4EYIrHU5FkPS1nU+BR/H8PBgLb7tZTv66hHyWqQ
F81oCaclG4glKX1ClHkhGIZPC6qDam6kGg2Bnep5k7Rw3dHK3nSSWxmASZKbIZ8qFSwn+ZFvG1bD
qOG5bqzyjV7rYWhqtRME1AzCLRJs+KQliFR8/588JykZiEU7G0J1h5yx1tcxzWF4/2KZ0+eb1ged
A4ehGL92c732XQ94hjGNEwRNUOAGKV6uhzBUpu1lzQIcxx4FWkwujZckTguBXM3SOJ4HLSusq2dx
+4dsrT0va7iMropEGvXYijlyScfPV0F4kBpK7HcYeTGbWRyv9sRYtja27CoVtv2elOB7b8fVdMJm
HVeJw8tIiuYJ6aUrJyEl5yrTDSiw6/71lR7X7kYXGFeeKDTZe+zXiAVAApDekRNWUl9/PeOf5P1T
1agTsiLbXczECJWKwXQZ7JOyPEBMPYen2oSojSzZgJi+31uKmZ49Cg6EEkWTjaiBu87ywGNQfyim
M9Gkut96BfFZbhdZUMjniV5Rs+xcwn+n3fEQ3x7j+OddnhjQjz8HYiZhj8a5N7O6KuXsSpO9tSBt
hKFpTa1ObkbfvnxF6IVyd6YjNodtyJN+mIk341DMcP5lLWcVOGH9n3dSmq6bGBzmECMz8PcHJXjS
N25oMucXt8EvLWkOWYAT0rS02DfTUBsE/9cAbXZZyAJoP8l/JMUgmqnfXQO0hWiXW4bPxw3AAyE7
V4u9JjKgw+aLUFZQmyKqENJfn/zKistsMUKajq8XsNmiRAtZ71kQH2JQNRkwP+859bsMQgWmCb5j
cY/RJE4HLWBFrq9Mq67l+vI2yvKQL5shPumJ7DCelKnJJN91Xt4SgfDmLcAWnCwM37W/yJxK/ftQ
/QHAveMKGQPYpvEDM08vPzsYK80X1GowX6dArEa3kGPrxUGu77X4VKEw0hltbTnGc6Xm7QpDhr/x
lNfXRsuOs+WstT6g7ImIb9cN11QhV9ZyhEpJLVZIwjKWQUxSTd8NkrO3KKO4t0EA2W9kwtfWDx5I
q4sUxxolubp2jzvz9HLa7L9DyIFMrEH8o1L23f+hu48/hP1wtdBMOysucuPJDZNjwbACf4PKlK5S
3KPyGT5c5wtNlpW/cKopHs7vY9zy0HrO4a+ei6MgdfwXqZC6fWkYLEeY5c3HglbaH3ukkH7xqygZ
s6FTv2Jww8TFjMOJ6bojduW/OgaV0jJTLofoNJa6QOCzyTVCpHNkH7A4vqrfnuDQTudd5HELEgjt
39CGO5FuQosavpmBSbfyxFeoHZwACAPP0FVfidCQF2ei1p4Xt7acw4vjUBfk45en4bDA8ZTB6IoB
08QVP9QC/H7oBfd1HUkzT1G2dRCf9azMRsum930CTp33ukSFzaa57735BwFM9Iun+5XmsI/WNeZU
NL+dm1vAsy2GFbTuYiFxjtJyiSHq8WCodo4BXH1pwm/BizNwBqA1tv0eI/USyvODJ2s2Z8kFqZUq
h+ZV2lUmXlMLx6l64AHjB64S2Y9QkxdGGGFA5wcR3UjZ4Q2mgg1co6H4bJj+gAXROmyUl7N2MCWn
RBaCL52+WEdUVP4tPD+aR9c9l1jt7d3fwvNVVfh8P8GAMGGKGtNN0lSBlsfkEffT6JlBHK5OhUch
4cOBmlwYEEwmgNpGvx7Q36SIWq8ibG/MXZt73kmJo3+N8gpX8lJCxcbg9dWmhWmqdbaBmvUY7Umb
uJ2lf2EQZxL733tC4Ss2CBxtYD2IN+uFnGO5+SoMDzSCwcx69XKbxIM5hfTZkAxtrUp17z9cosfW
qN6BufukDGf8F3i+lHtAg2SiFjYGem2fxClhi2Wmw2VKN1Gjaytaw5Ot39cMjd+CRTRgAfFy79I5
8NSvCKrNZlv8/BbdpvhBIIVmQmpwAIUemaNpdiayqsxd/iVms1kguiRszb0ZHUGp/yFTd88r4IGr
WB4cC3x+THzr4+3mtXM3REBm3B6dZb/iAkfV0iEKxjQXdpLr2eVDr80UAEZOLxKWLwZKCkLZ4Tft
c9tbmJYMCoExiLUEDYI2WKuGzHonb5EUCWPwqrFzLAU5e3QKUr0txoyzecwVT6WX26pTWwh9NSNr
zC5pGxjWHrGoIwsY0y24UIi76dCNHmY6eSZ0MDlZtn8PbF1+hmA9KUGoIP+RmgQ7hUji6UzvBb+J
uLDQGRY61AcTSp+K6OngG0EjCYsoRs6x/9zB6vSDm5PXI8awD8zzjFcB7KL1KHjDyEiohC3RVUsO
nK2mSKhm7YUqOqPAfbG2kwcuifq8+XdKWtyCn8PA0xfI6VoLtdv4rztf1p4DQBEez4u+Wd8+m0uS
DVmOWITpHjsGsGo8CjMlqTP2dpP6q2ymXBhcaYsZLuefewizPQ4x+6RfFNpeMjvtfdeFwM0fh9Ky
FJ+3msHY+PeRkXmOc/wy5O/eC8zmfH7WA9BfAs9aP3qt8zvhwVmVTzZxWJ4mSHr8QdSptXpzobou
Su43KK11YiNW4CGKpmun8jhu5z4RZax5JVB1C5Hccz+TqhzNC1ClY7rCoSFhjQfoyKdh1uCG8muh
XtNs6biW3t/2om2dZ6DfNPwUViVRsNGv4dCaHHa/PgmqHcTMh3hM5leIuPIbygG6fwxF8GaY759W
q2xj4XeiS6RT4EdhrL3wsJtqVDLhlanm+DzUM2Ol33qHRb3r8mp3aV33kuJqDKFk6Ftfjdz8HxS4
jvpH08F3Jz/IJuz/qVEY+Yh0FbQT5qFsgXOHvbKpqyb4qfCLiRmuUEne//+K1JkuIGQcJSEfJ/Lc
+YsVvOOPiEaljP+1QphlLHuIa9fGw1S0YurLTH9gzlIl2xyIG2ghTIHEcYrA3Dl4TtzhwsYizfiW
cPoo+zlOcC3HlMbwAi8XiByLnOYZsUHfJnaKNAqGspBUArAeuj1vP6ajS3HJwN/thps3ah6ftJQ5
1ppOYylo/vcJdloXM0MEEtlzZaDxaaLdANxALY/V9jUxh8MG8jNWW0YwvDubyWq0Kkzu20H8VQy8
mTJGChRl0fe2iTQUGgr4YvsGqV827bkmGI5lsGZDD2RC5T7T4db/4c5+1d7yZkHmnyvh6YbyESne
7NKDH8CvPovajn8o9VV2N+L0c33G63nEIsvaE8EGOUzduC6qRY7lEpA3OxUVV9l8eefLoWLnj+4d
cuau1cm6CrGWm2YMt4rnzXoUg4RrOBcrd69+zRG3sVEo4oJa3DoZxoros0Wwypo6SPaGAeG8oJZt
mLI2Dq8P6AnJALpQ+FKf5UTu7ZfVmanw+9j2rlVEa9Q2MHVQg1s0EHg8X9VqlHjykEqgAX2jW76I
vGJsA7Y9JE+1ATp77Ganepfz0MJIfjt8tyYw9IgRlXfvLayITk9XZDHnTs7Fzn4H60heSqY25GLL
0juD9ISbdEWEIsOMwHwM4MxWGk1+q4HX69moVyB7LS0wa0tOZN2JB9F6695bO/9hn8Kh4sBxEia9
3NUrqDm/ZBiGtNy1ea4P8/OF3GLZLERkF1wu7VxBuy3wlT0w8rgIaV7lwuUC/Q2qAcex/xWAZGlP
zqKUnI+i2IWSDoNKuWntveCZkUPLtHoOBLoKWyS3F7KIG0YubUp436/3fAHR+IPZP2VHC4e95VcF
LgGyaiHI4fVxXnknAp8yvBNoDMG79g7y/7+Kf6VGdNNfb+n59P9RyJBEYU7BPy8tjpJAGpP5uTPr
Ls57tUq6/CeKE+mc5h9/KoUZcDlHJQlVGZVQ9MpcfIibrU4uN/jojD0zwcJhlXlxAHRC00oP0r7q
esd8Dhp15pEj6ulhusxYNommHlchiga5LghaXL7z1bN7GRSKGKgsviU7bMoPvZB7my2ef/mgbPqt
tzWfP13IKUnYfRYLpK2bBXuw6emLa+s74FkobKtGiJ2HcVc3KjYFy2VS+W2UxXB+mAccsqfvsYuB
IwXCmGryV4YNWHbb+zmy8Vn+KR6z2qDfFZv4nPpW6wPxMpR4iQH9XeDDexbXhIbt1y1KXW+bNQZy
9k5KSXOJ8W8SvdvpdDPhBLgYjoxRHX0ImFjxl4RWVR0loc4MdC3398QiwS6iEo4zPJ74OJfgd2ch
dPN596mqLgZ/uENa+EgwPducoy/7bnpU03PoFyZrdGwX2PWNf1N1B41+tp2y3IFW+edciVxnNx1v
z1z186vY4fVoPbeZhqztthzHMVsiQ0O3BvaNADegHelIto0KyCBoMkyd/3dNZKD+69tx9FN6+ymP
Ys+81mbBVE8o8kAxOT1nvusMau1dmC+tpf8ruJ7Lh2gK6PwkPVCPEcukttYg5frKR/EGSad9r3E+
5MQNqOanJagMlwl4EgXcElCnYv50bTGl5uL/YGtho1u3Xtduuoy0cAr/2yIZ5ZuRM7JQRU77DvO7
u+SuCD2LkCUbJJkhiwYdqL+cujRoR0TgExdhnoWocYZb0MCQZ01qVzlzSAqQ7pZICHIqZzeNW7sa
3NDiFzRGcXvbJfrXxCItuY515JaFnaAERLFTriUv+rthF+7TGcw71PEQvEObpefuBF8/8IYQqru7
06UYap0hLoA5XkcIrFxc78nokyNMr6n9YHaPzVZ5xUtCcIB/cc9te8Y0Xn0Q1tvxYL4lUlSlHWN1
GKxG5jsDyoMueb1Mfc9SUmj3PzURtdoDBNyTJ4aklhUBUALSxHayP1UZC6YZH5gXHJy6DIAIaVCp
9tsx5kAmqVpf9BG1NN6U6tPSJxPCaKS9i2gNRKlyYEN53iSZMeLJqa5Z2azWPJNF0vLVgAiXNDm+
WTDdEgA2XaaRrzB8o5eDYPBCn6QsLPCYqwvrWw9TtSbYvsj/Oi5uo6ASfoJWEXRxvTg5Ai7JzaC4
PKADQvwhiPrZW2k3FhgPBp2CtlMaPf1M9CASBPsJCuLvCpCP4x1ilhWMDZd7wwQPVb693ON9eS6c
xiJnN1Vl1u2iJr1g0trCb66Joo0CN/KeoK1tq3l5cM4YDlPFUkLqe7MNQe17tiGaMrH0dYkDBCGy
UDCzb7xGI+GrKmrE7aQKfCT5/O+tmWoIZcojsVH02MbA32Ia7AG5I4wYOT9nuBcDm0ktGTfc3nk9
+eyzr8UZypo5fo8qmh93wYM8qO61i1cgTW/7lUNXLdzR2BbF/FqtaPH3QNaDvYT9jOP2Ohyc6zgK
d1USXyvOfoVlk4TS3yo1YzjiOf96AmsliuKfE6sUIQW7e+5alfJbjHREWY6Te7fUC//Pz+k/pS6n
/BmapV0IS6QQzun5fCQaS1tA7rj4Kzm0AHgN2PsEy35JZC9Ku7bncueKHhG2QptfnnrV017TMHvS
qBlC3P2fesZEeOQpO5XF0rO7xRgQtcs6GFKiSOMX0K6GSYlgdtUQXqGAXKVko77tAYkGT29O55qS
6vcQ9sImauY8LEDe+YbyuqDI5R6kRUe6DN2VjWuWW8GTHVVp350nYs/T4qQXY6usIWFaKArttqX/
zAWzo5rvTBKfH378abeUQPytkQibmpeex3nl7uaOpiGbiD7ZTIoORA/KVWJR5RpAoIhIdYJg5O84
xrFDfj2V3pvsbMhpBPb2yPFv7/Y8iuRRSC3eXakUkpE5610cnPubCwzjGcdeXhqmMuqc46IZgy3b
nJfCByNAQiWtxCvWjOfq8BLj3qa4x1i4LKIBDmxuhjhmeQGy7ARnBPWz+Imh5msFTQNmjBOQef8F
W2C6suDk/e2o5i0RZZ4p1tfZtpIH+gB2DHAEUaBFu6fm6cF3jLV8W3NVDeGMUmeaRGLRdVBkl3B9
5KOi7FxFkNrHoLtWuOA0NqNmukEA5BeOjBhKt9MPXIJVx3Mf3R9qWv9dhRH2a+LNDVOkGtfJnzPj
QQmiUkDQGydT+Xbuug0O4FaShqXkb2z8CPh1YwO2RpkB8Jf1HaflQqtEMCQRerhv3b5eoCu5rXUp
HSJY8mBXQ0HsqvoxwuDcILU5o/UD8DaTTfqCkK18DB+uMdLX3ve6KEC1lPljQ9dX3XwaqBVASRrU
PCZM191TQNlUbx1AXHYpBS1ZdtPjqmEKMTHm8PleQlvTzdAPXvv5QE+PWtsHm2nlxuuzEN/+nsvM
CKZrsOujjjI/FruxJxN/iaUYAFDPV1TBDwltUg5oOnnRaNg/z2fgnbfPWwpE6GYLBnccY/LCZ4e7
zlN2JiwLZvKirPf78RhM/Yx2D4wLy6URz0IRtkxVpZ3cK8+KoEljLprY06xMeP8fzCNpGCGk/b0N
6RFcfxPkifVsSCbMc/e9SeGoY/7e2hfByplMGYQSV9Nc6FTC8vWvcQK//hCrNcAJFKURTyuvbDHg
PHB3SeqsGsOMbqycZMIW9njaAk2Jo3N4iBdsGwmwgiamAeN8QzCmUfjFB3KWg1D08//e8VfYtWOs
dh3q0D/ivuaeQ8BCiJjMBfAYEy6szSXOzIODzgIaCB4Tk7w20Us6l/nnRrpTnHPgSMknMEh+A8go
dMG9l+bU/VmRV7Pw8JGaUE13aQLh3PxOThjUQUmMovAj+6RHthRF482Ro+F+e+wDEPxVKqoh5cHW
jzmEYC3ZbXVFOk5Pycven9ygoxgfRQ1gJp7iokp/RKlfg0eIDF4YgAJHZszIPl2HcwRWyK+DpYke
ZJ/oUCFZldgUJL/eE75ck/TNSFbkjLL9xqJ6HWqtaS8O3LXmH8+rlnh1fZ1x+kxUQjU2oHYefaJf
R4YEjoba+9/ndY8yjWBpQNNtKGeW/5GyGTJuWtPXv9tqeHr8AmGUoRIJeJXoBDrfPg5zsNuHMP9x
5VoEt4jwbFxAna9OhGNQ8Nk3cqbdp3oVNl6mkVyMPxAzdr6uD6btxJNGUWWCJEi35J0GfKeeEViD
ff1+4o75X5XnzyYJkzGBdThVz7ZFfegSH1YmlADFkKCxH6AYGxXWmCP8v1Ghzz+2zB7f1zVqdpr0
0DLSpB7EJQSCUmCthOwC2wvBR2P5QzKrCQnjwV5l5Rh3FEk1QaI9phQR/7jW/iO8DT+iHAHQIryX
akHVIFmyiAhNTYuah5Il74VBI4/WbzfiDbj6oALouteajn7F6ffSFg78HUGHHnTkm6c2/3h8a7GK
BUce96/y9+oBDycHtJKy/nzeIZCrxEORpAbNcpurIU+4eBb/ASTgR9dLJ3mOZls+E92jhj3ua7JQ
QZFTXk+8X03wFl7jEWcihKnX/am0JvUM6z93moTI3MEOQW1PAzVh0CbDPR31ocRslSNWAJbgbkcL
olFNl5Bsw9bBZw0Eb95T3oJ1+e1ANBtVcUBphGro4GYbUHOjlAM8aSxP1hgvjhvm3HaPfo4gRti3
O6TMZ5rcRaLmF47b2N1ASqSgTwWIhyPT0TxAAGna7OogCy6cYV1jG3IM1GEh3KOA20BUHa6lQzdm
fA9BB/N06owPfZN98Gy5bXb/xBcng5DtHNISlYcrKtbvuKluvUhtYJQdse9lm4Lkzt/KYDlil/Ux
k3iSp5/IcNxwL/XKwsUL8xuXS6WruYridvnAT9MqhqaYTaX1XkitfkkPfCydPVOaPNadwiAaLBl3
R47C78ik7/ZvvQCJ84oKVNqXIck7RkK6bPE+g/95kfreK3GHYF05/A83m+zpK41OUjayKzV99Hkb
au9ZMjCWjSznGhEu5cSvnKeH3jvUhZeoLDiWIsozCTdUHDJAu24OrlUL0FDQ5rvNfSnlbT7q8Qxj
dzbg2o0f/oa+++6GolaUlBCuMCW/+c5RX0y5X4u4JUCAYKJj5UF6IRqE72VGirResqrP/lsvrDpq
bNtfEUwpi+mWTitvPvVIDFKPhyzM4YmtkE5aQjs9ssV+QCG+X3h5cd1pOnypDTQM5kScmkGiiUyq
XeNTKdAhLX8/4ASaTGD1D8s78PUfxzBRYcu6E6Kd3BjvsH+JtZ9qvpjAEZNip0Uj+pwQ04GO90mK
ERe8/IFnKax09MxwIeq3tV4UBl7TClU4+Mvh6xQKTIF3ApbXm2BxmeHQXRtIyeH6R7FqV1zAvnh5
Tzz8XFhitQt2aZYgLonMqrG6p2OaN7g6rTgrmnHtINKXE8KJK88M9an7bktvnIkcvd4JQTS36e43
fthIqy1eX0mXRB1TjF3cppyh6BqKWJlP9WUyq1xqkzptNrYs5nQZdVZhS/idN85nZa11pLXZIml8
15F9MrtJoO6L0z7g/NY9AIXUP89S0nDeSSbPydqNEHDwNBNuTtPFVgnMUDJVTkwEQhrvQUgPeZFD
OC5NkkUrfkkm32qHDT3cPBDhjwmpd3Rh9s5/i/PemFKSFqt0teLGLvKasfowuFaaZPJLQMway/Gm
0pLnkByCy4Y13G4EZbrSExd7jSj504beVfHzxmuR1fqf6wCTSk5BA2aP+R1yUQwHLW3gBRJioEkS
ldGYPwtt8zkNLjp/fNhucCcJuwEwAHnECbvvT7aV9ntSY7+nYE+mBOqX+ikmwx8U4CFgn2vJkhXg
4X49baUosXqpeVWltwmcq1m2J54lP2/REiZ2Rwe440LFR0gjnlbBjlZ9sjw486zO51Xz1HCt4t/A
KRofxf0qZAgnEhJNElRzti0xrB+aNt3jnHLa9UQyUlybG9M02zvWZVi+xXipbf7VN50pcp3HVHbT
hAZzo3iimvNEoCYNx7DMaMVS/IYHj/7oilsBJFgoeD6fmV5HwJgoY/y5/CU7+4xn1Plg+E/e6tQt
4JmFIi+cisruIekxrfvgONA+pp+6P8z9lyPh2Fg9M/gCVn5DhWcgBFRLjAyxwTDnti0Yvtt9HTBo
Em1iiZRygtzPvmlj0HXV1rA8HmR5rmQRA8a2njr66LQGxttDTFJbXoYKylFwplKSl2P8Vk5qw6Vk
GkNXX+2RIQY7MYknuTssy7RccXhs1fA8BKcmzK2RSC9rW9DAY2PoB0Bnx64mH12hNHim1VCelPJB
VPLsFcbjr+dZQQ1YbQbGRH97F7sY1s+wWpmyCCFN+7mv8OWj7iKm+uevvy+1S36WbBk+o9KvizYR
lMxidDbdenP1PnyRd9cFCqaW0aeltzDnLWHMssivv0X1aa5GCU0vz71H7KD/qP6bOlQeNQeoaUZ8
IU+8gGep1BlL/tUZsqs21LTvB5zc9eVx3W1VIkC8dliJAgc85B9ZCWkB+h3wLRXVI/IAX5y9T0zI
EhuMAsKwDctaMbIMUeaS80svHQOX99AGpwTv5FGC5FqrL5giLFhh5WGZWTQu+j1T3AQKZT9SBTMj
iaMjmGez1MeZ0VLaX9Q4eUzzoMw5JJoDHdnB6y02h9iI+T+Mq53z53QgJweK/+p+wNzm3YrKEaSJ
fhbAShlG61A0dR9wpgy3lNr6f/luOGUIip5UbhrHTzcZzpSkgMbqsptNQz29zI+Dw3qlxdso/YEj
CCyXQMBKEjdEpLhchwgyXqpMsCIOKgP8wStWapsYnQnfBWkrwJ4p/zFt/JGHQH3eoyFEByjA+A7A
wVol3PX+oqennDtK5MiiUOVSyu+SnPfCK243x/5M+7tHDc7UvQBu0ltnUqiJ2VUdisAwXx794RDK
YjIr7xAi5UjBFqbziHcdORpeKFLlPtRwWmsP+eW5O1l59+s+hQRl2Ud8ozmkHEA6BfKW/bpP5Z4/
MtzKW36fYcEMJKRxAboiErKDcd+jpjtba1gvLrnDv8ojsjUVUMm2jIMfQlfZdkQOd9KIk27Ouan1
A+Fg29dYRv3KcueCm2x+u5phn6kNRvxppXsO2sbzeMzTFggjRC7Uf6dX7FUxKJThpJUdbsh/94F9
rh1mCPRlpZBLjAQOE3nABhgk1dXXTvCAxlgdeaH+qhWXHmF4L5xht0VFOckIFIVclacl/5teyXYs
avt5do7LVIc+64Iqrv36duYzdl5yLknzUYd5SrOaGs9hJ4D06T+6uJNqNOVhwxoojeSGwdxyVY6P
E0VA0cmjUCbxoWHnTXE8AZWtPiWimsSRzQNa5VwTdH38DWX0JVpSSEXQIjeU7fRTUDuex0CC/aUf
ZPDiPcMmEpHFX8OBtUzmrbNQV7+M7B6DBkENpR5dctBl31vJ4vVakTqn5bOR+Nf80HSpK8kqrevQ
ByrCA1uVdeFSrm3+95k4buv8AJznZVnQn4p5s/WxURQs9HrShSl8AelEBc8/EC3zo97qcJ2CCB5c
t/JvYoVVxkVRxXo4yhsx6x09AWNw+rn61GiFobR2lnemqKMXnqt+lwnUn15y4+c0ThY5Y2s+8Tb8
CPM9S6zFHeb2hJtASEvu0TuuD4c5uUgbKwXaj+4jMcJJxlmmajdjK2P7lIUOEAMcRbT1uJgUZkZb
eF/Pw6jTn3nBFuMBNudNUApE7Y3YRvZt9l+azfTeAlrm5HKXbTgN2+tA8J/SyhghaUjLRP3416fm
c3CxYdCXXf1kDGUnqSh6T6/60+XeUs1sQW63GMTyCt4SItL+KzPZlZt0IIYn0YuiVJks4Sz7lqlF
39wbHRohTL1z6MHHcZkeJvJDTSHzOUCyc7DJrQ1oPf/KwJOYqijcRRiYI/uZhs4Rk6qYYbtrCfr1
imL3YhTw1NSahSKD3xZ6EO26oGDr+KLXF05IjEX/peCmu0pyWE1nN/RgF5OmVeYSJ+R4JW5zGK5t
Y5JgZ99UfaZYOycH2dlsfjoU5BkakeKhDBVOttnvcNcTp+9Tq3HvZpswOIqGBqBL6LcGHBLsS9st
g16FUgyzWUuM8R6boYe6k37gyUVZzmZchi7RSf4Bcgr9Q1D2hUV3Fqp4wX1tpIhPZIhRpFCi572N
PwT03gCUdVC0Nb+X8XfBmPddPsqrnYK7SEleEcNO7FouftFz2EmcdSR4xTjZNLXhzfaDqMZxnGZx
/OSgwiJpNjXbutsvKITnxHa6seZVY5KeEtPoc+GAiDzLLnD1xBoAE37wnMzvug3+4hZGfLLjhJR2
yEUgQzxptP09HEmWO4YPdR/1Ie2H6J+fI5bBM2dtZTIOeNBVgyeD7u0Ujr0N3hJ8JpfwR8Lajeel
ahbGtmhr3/3fUae/0NmxGyAji2ECr4pAQRSyBhQweyMELqhEEHL2cfFE5FCJH3XbZ/zfiK/bi/80
9DezJz+y07el75jAYrYOQ6HARd5uNs2P1/YQAxjAkp9p/LkG21l7TutaB2n0NrRaMipz+g9KYfka
7Ou3P4ozj4Bhx3JKrN0hNsfR2cPPSmnEU7fmhjUZx7VKUYttdXzU6N/JUIN4Wua/NmCdDWecyBeW
Wxz3PKuJCbC0GY9eab10VuEPJMV/VoV4mmFRjOJYIlwadwrm8fXt6REM+rJOYKWzhKy5tRQ3eF3p
dzBd2T675AgwbXvrZHymGJ8Pwf3yrYzFkrtPi+mNwnLx0B8u8IYe48iJosg/AEZXVGY5phu7p0hY
M8d/f60llMYmeVabqVrVBe9zPa6HTnhAhfCrGCy1XfwO4UQ2iuGuVWXQeeGN+6RKsE/VQQcM5/mb
mMmunMefnN9n2RgP6x/e6B0o1Cmv2VAlMz+4Ci8RtGJs5CVYUfYf8Fuc74835ZoFYoFNwndI604w
nvAI0zFmoFGrH5IajZTeQEwasm97Yi3beoLVGYtFfGh4BBeROkmStwhyJdkWR7fXUhQheAcgtklS
Mu+3jvkq9UTwCW0HD4zo6g/tYDWX59MIeOXPnno2Y7+2yLknz3NszqBCqGdvevTrYlWlEWjk7UEC
ax3JvDGNETpHusjznITXP+KWCLi8/bx82Lu9PnGvSU2HDdJGm5pviHY2ZUu8ffYoiUQVXf2lijiO
Q7gOAXkZ4qlZwGge7WBreHDczf5XzCn+NzkXtEpKt5p8Jznx1dIsw+SyE3xCUYx9tQUpl4dYqsjX
OccA3pWlCgw48UKOD14gqxEg0DgNstco7A6L8M3oZOk4MLso1Gi6LRRquZ5Friu/qw7cTnEm9vUT
fgK2QW4Ck1twCe/Y8zJd6QKdikczCKgh6hg4T2lsIylI0XQnWvuaHIF6fCJj1Yq6tcRN2lX4r4T6
tx2CqEjRfWbFVGRMAUpIZpH0KnYWd5mxHYC4PTRV4AiKQ0jNpTTvsIAAWkHXpfvmR2MKPi82XQdR
SnH8FRUSlDziMaQcue+r1swMr3+b+x2sEpKLlWJVp6KoaWDv4q/DAdE+IShLhyczHX34L1VrSI6Z
bVGrr6JRHKV1lk9HoxCHp1IJf/ujYLYpEMR3NAhCyCYlmPRuJY+8kTgAjW78WsHOVirVFjtYLiqA
KaUE+kTUuS8odgxycy2H50YDqA+ImKbWfRpYUvX4Xh9K6SCP4EbTjHMV5pZabUxsmnPsN9yf6YiT
NVOXHgWkJoSVAyDy0ipRjkqXv/WjlEtftSn4lACr0mLUewnfXabpqHAA6JyYN8r+ymNWcYplQvOJ
UxyxsGW/48MYJ2thGymSqXZs/J5HgaLqA/ryRlzmKcdDhDeHW9X09rDfxMZb8W0u634m9uh9Aj1H
yO4oGITrDN9r6Id1a7HmEjQebaxa4rHQlaX/SxNUu1qCfpJzsLluHtsPn6KfKBxeIt0iomiiYWxl
ETpGRnLe0ZYutlctJwR1cL/R2ND4m10CdGenOt1baYjfPXdqHdxvernydXkSSFDgZIKnhVAXmd9t
Ia1MazfPZlYriKv98uExjk5XrCOo4XyPnjQZdC3zPLLB+V3pWYe8+n33vqMTi+QT/dzOQAiggHVg
e1hyllCNLkQo0MmEc43u99j0Uc1J16bqHDXfLI/18W5PJNbxguQuQSTzgHz2fekyhtQCyh2Er2Ly
k9CsB6sxqXFK7IXrs3vg+vtvqvzDncKje6zd65hWn+4PtXDMxh0UyGZ5OGSTcOhy33d43G79+6Mb
8jxH1BEb1EKL7H61HjYKace/g6xrXUdKmszjaO+FY5oVVKL/7dv8iR6vqXUmw2/VA6Et/vfDvtnA
POEUJ2ON1Bo4nYybS3Oi2YWY0HvodIqMaGMmhk5jyFWOYgftRSPyq2Wsgd/sf6TJG5rkH3yJMgsN
FKcln0PN1u/x+0p1d0EAIxLvGz4mZ3jRIVsTBj2cURFRMlrjmfQdsOFNFcKHvk7gVJOoqZyFpBWP
kmt2UMlry3Dejs2Lu20jMg6fz6CM2s7mxAoieYGMPjlZIXxfCI4kVnU/1ZqGHN1FCVPjJXHIJgrd
28j5t0BPof4odhK2kV+CtzBM9+2DV2Il6SFUqLwSgXvbUPrsLRdG3nUCisTXbKI6TRUia4635m4g
KZigPXF+Na6RkNtIJsxSoxLY0VP2wZ+WEP3XVXfXNCSn0m+K9FERM115flKYVDEhDVwc5nZb7xc3
KDc1hcNKTbIerBGFW+xfNJe55KeT5CRjDfdGHSqmn3mYW9dLaqIEV18gKtm9AGpHWabLtcnCSVIL
BleCbErkAkhoAGtRqBAVIqNTpGdZoyCtwY7p9n+5Bhc1ewYN5oE7mLNB0HLXOZiZtFfWbij5hLzN
2Mpx5F9AaSwStaULj2G4aBUUc/YjuexfWMwUsB2vrENXuJuKZdk4BzNUzpK2iVrOf8cKp1lkNlYI
2w+rAttagpiA7nva8fqoRcsdO0tHo69iolVO2oAQFCixJ1GP0MS/23F/XsxhHl7BvG3P6Ouf1eU/
iwGZNKSiUpWKcfYXzMmebXXkpf7UNSILKIw6JzpxtmDAyRj2INDqnm2P9sTUhot8BY2jrZ/P4gax
4ZT66TBsUtmR2idtzqlnbGum1HjSxN0e7huvEeBJD9QxbG7u6/TnIKOo1XxwzcO7cCF+DG7wNML7
1FVQayK1cUvTF/aRRQkrpV5WNINh/zJko+pcAwPCiampL9kl04KgrKtX1DCNvehOmZMp9yrZ+StB
YoCxwYTeEJQv2avPVoZH5WrXqX5Loj54Ya6FFlJ4qUKMnGFyd/dwpLlGLlmyWFvkoQdeJ/dRk/jL
IXfVJzFHxgrfvAsnEXr7aEPO13syAo10R8ZHSZN/7/lNpK/3pRm2DAw9kM1dEFg216KUVBIviK4L
S+BT1n/nlOoAdXhzFYnr9V2K9BsoG4woo7fniZQxxuk2k6sDYXXBiC+MIChx13U/shL0BccOuHUM
pkHFCVAyH9Fb0058QjrVQhvNnTUUkQoCrj3X9WDywIre/DKn4AMX2TX523mKFCXQpgS3fuaKogBU
0wBB9pGQ8IJUsGXpoKQl97E5XmNQcHoQ5Y8ICRQqy2B5vyPX0XtDx3fnx8EjW8I7UAGlZri2hKuT
yH2UfD9yGywL/pzTacETMWcmt0obSqNWS1bsfkbno96GDi72rI6SOPxA4rgYP6OjjcF3kFmargej
/X/EcgEFiPsAgzGKeOQHqgXjHY8NMo1WyhCkqqlb5ss+8p1unRobl0l2BSUjsRucFhkyzpnO7wbo
t6yi8T2tAqT5xoJR53BZTzNEOWj5VP1uzUthONgSAW9aVCCqqPfFh9brGa+iYXnudY4IVZD1rDwm
jNV00d8lffWs+43Oi6CWuTLej72bHETk34uUBZHFxnMiWDxGEkADmBKVGUxwtcrr+bDQxUFrYbXg
szPh2QCeUWoS0rG5OzDQkZp8U2IrNCQNEJpILfCiIqfKuz7GjeUDC31hd4FLeTDWMxEF6iC6+fle
ImtXzkgAwdjt6Tn9OBqBcGUCVEzmuMHNVYPGLaialDo6486Ry+ySFqjAhFAbVzGF++41su8PTmP0
xywtxIualUp7HwTw/vJijz1r9FGUHC4Bv2CKiPwHPwJvqebhs0IzJom7I7UV1koaPIXyqCUOlo23
s/uohNEAOLEZjJalgyopDPIvgvUNppsFs5a/xf/HMOo4nDfyctxZswRTuscnfA2Em0nqbPvNwW5y
6mB5r24J3Zg+iMhB0WOr5AntHLxZDwIiUHEHJyetvxY7prOWlmi4PI42jRPrK5k8pNwwnQ4aIi9N
3xXdR/TIb0nqkDlE5xaGyr0EZg58W70iBDetx1XoMPp9XwH0QhJvXMdZg5rKHIVf7t95UWt72z+S
bxNotdXOtZhS4egr6dk1DSsaA7gl9/6AM+zYVBzpwHRVd4+tvPcLtlVRysdMyyvrMH46oOx6cCrx
MOSqFQdZCTIqtJ/mseDurtZrYu3l4orPBaS5Vv9571OjaAfmUB0jWJaZKwTyG3qwJQh+sxPp0Az0
zlMGflWMYxN92CcyhkfyOWn29GWq3jy8gWxSvs52MGBW4+U88WcGX93jQx253bI4rWWyF6mvXAEy
ikqs6c69hDdn+lIHaEOo++jOoCWaIBxi09Z8BQRzXIXWA1er6HsZsWlyiFu3UfO+XfFYajx1mNTa
VXpEf2S/hJ0Y6+8/d2C1aEkWc2HKvfGneFvgIZg6GymiBC2lS572ZSN8M8KzgzttLsIPKFpNnRJm
O2hZ2BRXe76WEIRH40YyOAmtfGJS0QCQG6qmV6GtV57dZriaDfJ0u0p9MWlFW9t7qbAVhFsi6Wf8
JjPrbn8ArCBHIYkNAmPsJEEVkznCUtXmL0eZ16akZu3/AjLu9QN6isX6hUDcsypIUvUwC9Fvj8eI
sBxoofLmFkEofoVOLqWOacF1D0K4RZlZSTYmHNArZdAu9laUWAG5BsZvKs9u7dyYou558pGVb0y2
4QXjsxyllDVHHoB29ymtpLclKlGIChxVad5xWpzsseG/wiChWFEZEtfQSG6ls80OmH+J2wHAKJhP
zvRnQ2evtOHopHEllyMSq8UX5llP04mdK9Q//oNlafmeRrncp4W7g4eRLM9fIoSfrwUmE76Bw9e7
Cd3fiUCEECaJR6fXGCLhOUnSbTIZuJ5i2t5UX81iv1nn+LfaLrRvoZ6UcLKt972goGyMNbrq2h3E
aaeSfXTBbIpI0V5XL+bNg+/Od4979sngmFzcLzLfkBZcU38ekZgpJF85eg6qHfTuFo7IPdADDdfr
nbd0oQJIuFqF2v91x2Bn1LbSoOVcSuJVX1C0SAKA3J51i4P/A4BFv21LF7Regf188MKy3FAYzX9T
bnaOZOeX0sYH3tKCgH18vDou0ySqiQ62HWACttH6mna6U4Ym069slLzguNpRdwSw+LCEPzCjEeNS
gkgNeNi2gpdh4xyxKjpppJXAfnuX2/nqZw+L5c+TOXH5i/8vH+UO79nD5MK9uAj/QyANJRD269kw
vQAaB43G4TlWqXKWfkmcmqNm/MNbdRYzi+vZIULmrZtdx9MUhLs3x4iZHzi1VqxI9cEdJ66HUFOV
R3qLuRB/k1+Ab3egMrwS07PVqcec+esEkihNEgLdBL62rsXROjAo1nv/zKJumQMzMvLb1KpMiCAi
iLd1/vmf8+ounaFK6hzIfjVXRjNnqd+YaT22TnoE1veJWOhA3smKfVPrfyzvBxIeyvk/fQqsm5uu
z/8q4/7CKPUXt/vn6BTAZ9o9DZT7MINliyITypZA93250qB4ALI6MLo8Sro05tVYBb5B3/9harZu
xXY+6Jr6gDlEEfTt/y31qsfzubtua4lzaiNOm6ffp3B4varc5U6YKdAsBMAs1lIm7OJ2fBSCBd6H
hNVyv/qC5iFOJg3RIXw+wAx5WALAaFZKaUS5G2V+D4l4JCmG/apU/NNLhIxpLNlZ6KPJlOsbGHc+
tBGeKlyMTepVHr2NOpsEJ1IRekgNG1Kdpo5qkPOIwg2wFSfuyJF7NKZH1N5U+sFjsQxwRTQLNn7f
+7rmZaCh+h4wr3V1Sb22m/mGVEx4iPiKq9sTTgzqBZ1EBX/EYwPmh/4Piq7/AuUF0lWXf2+E8i67
qLNotQHTnfzlHKBMaE2IUh1EXO6FetJoPsKQmvFWHLwxHDGj2LnL5Zgjt1vyYr2M6nRom0EGfyps
Nkmt5tf33SuqShFvSBgJTTWaawW2kbegKqsNZx0V/7vcneOtTWOL+mRAhKhAoZqfBul2g8HJ43Fv
S1lDXPWEBqCG8lE5st4vTh5ivpZdGFPCAzQmLmwpaPW+cLqErwCR1Gp7qViJwkxJlsDxh11pnzNO
F5jKOR5lV1+vhe9QhaXjZY/ttHGsjDc0gBAfMDP92aJVPHMgoK6/j+Dfd6vRnL6/Pp6PPDGhBeeI
+Fu4xqKrxVLBWV39V2ufMxVQczby3UyFIqc/Bgqjg0b0eOZmVB/diORpJ5ihdP7AYjir+qg4Y1RY
mtsYLlC/W9cPogzs3tccoNd5UtDtX7tvhcGJfnAv9xpE+5RNJuAsG61ZcgDGMhJgl8GDjTHWdJQ9
fe8R3NEOuegzhhH/gNADMpL8MVgks0NWZn7YhD8hUvky179l3yvS/ZaX7OIFd7tALG6ogHvnF5aq
+3fqp4+siGYTNK3FcjeDfFx8QdMmvuCLhXRhONgVByeh1Fv02P+HF2Mt9Y8hAOdAWU+JDmD04Uhq
bLJ7Z0w+zCp4WyYxj/HrmHKJx6Gfgit7JSt3IsUTxRir+rHMjAlVdUgPp/Ge/fc0dSak/c+Mlvw0
u9xcuF+IVNI9yDbbe/Anvw94soUKKQSWkIwqNayMJive9oobrhMPI9MtFj0JW8gXvdZR9qG5ZybY
HrrTvFfUONhoNhkEykaRrLb08jMnOxyPsutQuCZ7QqI+xshvedqn1D81KQriTCiXbzHcTgGu8bMk
t1u3rgLiA71IdGkyBFa2avUKjfTlIaRaYJpe2uKZqOe4MlnmuNil2kMXF+qPNFhjw4uAorCfoLBQ
Cgw5z/wQzFyiB0LVf4YiGuEgJ67/B+sZQjKn4fWnKjMtNNELoAp1GMo4cyvYPgLqziOi9MosfzpR
zWScL6n76v0SuUkz//n8uikDGiN7TpEK1YkuI/mQCS+wyaZ+MvG4WDy21eoBHoXWsJkMDZWYqqXj
L2QAkVIgJOJw40lT4vQkCC8ralEdCT3a8Iy9h6tGxZNRy45M79q1BPuzTRx20uZ6xPgJScOGmabc
/odsPyyGxVgr9K3JHqL+4OgNNTm3YcdXeJVpUGw8vSBcNdqyTr4thL1ydWnLZkOWEEQdFA9eL6a5
cvo0miqzsXs1eqB4qAdfkd26er6Y0xQGYKQC+qh7U/7L9Qf6vg/cqU2w8FQ2XfQaJ7Eofnn3WyYp
ntUwMbnCEs9Eup+iqIq1Diu3kascRU4Rs0dkfLGrkuhsdKBNIxTaIv+8gO0t8t8ODvwNcjbDS/C+
RBQt4feMKjpnXeiWf4NMXh0QagFertHFWhQSSSWC588Xeofn1BFZdTyYTwp7IHBsUANi1FpyEonc
LsBmKc1qFQzJNfKYpALww4gDbjpk9JgQOZ4FwKOIcoJxzhC+1KVl4+TUW8ydgNLq0O4QZ+7Mx5e4
HmuKQqLvBSxpE06aAOb+CwgVJrjZ3loVLZ+VQuF9f/zcfHaw7MGajgcw+CYeBQndDTP6P2gtUjc2
6xe0bQrnVrUZBvOG3G/0D9Q65XSzduORqIx2Tp8nnz1CGOrVx9qZdM8zurArGbJgpcraz2ibIaAe
h3pYiVjATDi4/NbJoI9IzBn2kJodDgz8J8i4Qq287BaeJ4lxbZmFlfDr3pvIc9wZTw8tOAomJATN
zxfFJ1dSwSOfgDL5nVQfcw5otGuGrn38a2oLXyUp/7SsMKL12QjGvwlOuFg/sT+b7CBoDQJth/xE
IjdRH1fvlu8TYKuRNGXV8bao6wdg0RfIyORq5u753lBg2reG80OsQX2nPPOmcrqROHG7GsKdVkgv
Mwspw4RSr1RA1tqy0nxRvKHUBoJ80b9aASYww0iZuCLPkOLUh7ktRBGFmr9UoJXk9KHy5e7evmkm
gJX3CHEYY8bZLyRghlN+wk2KhOBz6bJ03i0YOHxv9l52dtLJ5Pu/E5Twm8Rg1iwKsBs3cDPHPPG8
6dD/uqTo8fUNLk/44C7a2ofkUnsau3mVTb03h81igyZb0zFD6jim2l0xdUkUWFgdHH872+WXW9ok
QtaUqY57zUIhaM5bvyC94OudzK1pagUh4MB7AcRRqoEhegY/qZI4CPKI2uLsy/Lre0/IFcuIb2bl
VaJxXXaqT4K9rDsRy5OnnFd50nErmO+yx3xozUS+gIZwCAkw+z+O9T0vCA+QrvqIIFa4WvkfL52N
24e0BnNs3d2dZ6WHrSNPrYFj1mxphqIBGS4UysflWW1DdDo/yWcUFlWwEyRTIHyeDrUJmj+jIdhE
dkFKXQ841xRMLUQZzmdTE4lw3q649CzrE7DYOD+INMDQuzwdAhomHbd9+USZwEEhOAGp+yR1uqud
DsfCra2rnkdJACuiLNmA2LWnBeZ5XknGXE3utDdtEwc12QkZBQyvZ5dkLPZu/7VD/XQ7FeRRJqpS
5/bI9hEHe9usv7aJhQBgQB3pXrBDqerK6T+5NA1mNq0lvlE3oozazgJm6JtoXvEHp2qib2U9w5W/
HvmHstOfRFbGt6hpqrIJhYKoILViCi+eMml82wGxjyE2fPHPQjDszAEthFU+wNH0Kjkp7HF/qSer
EWpTgWR0zb9ojAH1hBTi3wEwftWpD417gVRHY76ow9/YpOvQfu030ZIa+TTsVIeIv3DmKCPheNaX
8E6hcWNvE6CXGICKwmYX6S5DSznKaWsMZiwueKWskLCDYDh2iPL8i+hYHPc1P8AuKTz5kqygBEB0
orTbAW0paph8SCw5MQHXcXuZ+egjiWf6wQaLXdSBW6ByLtCWytZ5rje5yLYdvCKjthADli6nOsoX
YyoQ2N1gtP4S0SdnfyNYZKDuQcUAGpFvxR51hbE5Rk4/Lj+q+mGmO29f4O2jUW8j7iGeEjDjMod4
LkIeE+dscTlCIUxX4WjS36XlYDWLrBQmYo7lA+mkt1fFk07qNtHClGjn/Du8zUjEyU1IKz6SA1nQ
i3blcS8Cidp0dxXa710xA3mCfe/XKdUz+5NOqPBwmcnYY8O9byaUC31w+dZhHpntlaxUT/y++S/b
JZoqKCoHPtK1fvBw50peELSGd511Fg72eC9+lTwRG/n+nOkIz6WWqXoy/oWK2jcgsAFLQXbWm8LR
cvyGFGLhnt/Y+wx0jsxZpL3msBgNCRSgx1Q0G8qH2VItWEGZyHFhGjFzBW59uvnoG0LKSS0xyBlu
p6iq/7ZzC/jZNwlhMIJHwMqgsmX6ZRY3PtLGAKFU0dLcA7tG21VrIeyVB5zz/tItIk7tvOiL15Cb
onWq31MZuQVaXzP5lxq3Bd5l7uiRoaUyjb2pb4ddzs+qgxfAgQJ2xXcBW6tnTsye/VZNYoLnOG5r
gaa5YJ9pt8PfumzYEWVatTJnPmTZoG5lgw2kbnSMVTksGMal6FscA+4ho4elS00iwpHRNErDPl0d
kmUQIv1LbVqPDD7ZRWNt6QMeDRllJ3gCj/h24/jV+8/wQlA13Us32BN5kSsn0UoiCDGXJqk1VJ+1
z1AHuxCuk1BLQOftwlGB1Ihlz75UwIQKb0Xvf25JhfjH+SX1puZ5vpmXmAUiJRXyF28Hy56U0SyW
cT9FI9rFO8ioIfxud6leSezUDyh2KNooEtcs7/4oM9gUAPpTdrxMksNnZ+RQ75YI3WTYsQeJaDNQ
0Tgsd50kzAGjclqxBLsPDR+ydam26IUKZy2Ifc8AfD3xs1lqac/CIG1ST+1mi8MYhr+CBjXnQc2P
yDL7WJ6KAmT4beCfLBbcu+lYUdkT8azxqa6BCj0Te+y55Y53Q96yQlUEe9XPR/h5GnCp+Br4IAe5
SK6yvMktBQqrqbRObBowT6ZUpvcxHFN9jzdQzQ0k0MnuJWC8NlW93DwUTH58D6BL7DuK6CvDEUCA
tnPCWbMSVPbWmsFeVSYdU1UfLNzblgDp9E65LKusm+aN48qeVGX9tFjfD4IRKfG6xVFpwv9szdeL
T3nSiAy2ssDVnQ58jZbVAu9Vy036caoL0BEtud3l0qhieXbDBthFneZc5cROc2AD0R8xHh/EMqof
t13rpSfivyC+o+Y704PbQI/mkFWyH2TvHJYzL30uC0CeA3so6TqlJswgPhGWRT861KhWf3HpfpO5
ZKuhgPAqUTKsLnKfUf5q8kPHKmMl8WoIZjIkhIC+A/i1R2VP8UDcXIlnLEdzDSjJ+tVK2YGw7Ym6
HaqWydc/kWfX4/JZXrXj4eWy1Wipz9r8U+IY+TMKfLFYJ7GuSHJN19daLblUN2KmbZaiQDLSpb9z
LEw6afIz7ASPPR2WeO4BoDtAazmRAaCHvQEutnyKYdxrLmpr211TD8AyWI69gnk1fNYKe4zm81gz
RQg5TWRO7yTAFJSouLY9UF7FZUedU/YCaQHdTq4eAPMTW3fyEqSMUPgTpb2pcjNj7yDQGnU7trvH
mTZeUJgWgw8kNyMBjgqM7RE5xtsMLUz7mfnKnVzBZItkuh272Aa4dKPXjYSO2c6lBeCyjEdidxgI
pPidV6AlyY6TQHHOCIEOomEjKyEX0MmlFg0NJNdmyTF2oCgi2O08NwYA1FeJYqbj2Q/bew+GQF4k
lYFIGqExL2S56LZ5KQEGcuRsOcABUnb7vadIq4Xzatk+nJGO2Twm6Hu0XT/KY5OZCmEpcVCWwR3W
Zf16T/Fomi3GWfin6Py7yCxc8aoHNaicoeGjA9ZQzQl2cRFIc4n5t11sil3MXtizuKuM0nLeikLl
yLI+0Sa7YsuYhHfNixa4nKBCc/I0Ra6pAxaiVijpLjuZ8PAiwjouA6i3Jv/bPliSLGUbWQzxxCCW
+OiGccB4RldFHqdjTwN0Bu/pR4s6RhfB1Wbj/Wm8IO/C88g7jl4M2IfJ0Xpe9Uv3zdu/fQccex30
l8K6gFTAzsMIRfdQOokkIcFM8wfJOExTO3NOEc+KOa8bxgTkrM0EF1KvwUwjpRcwrdvG3iLP0sVW
s9U0Bv/fMUxx8BLzZ8l3eEZofPf6p5GYcj5u56wXLG21e+CuVaclzfgwATsMbzgW+cOvtcY/dCGY
3zg9ZBvwlhPjk87AvlbiOnKHr6O1QyEwKrVIGGep79LDK6njzbGeL5cGtiOBu/pXVkj4VajmgJZy
svEDoWh4LRZ7aJnmnt20XKBgBBEqA5/5FGKIl7b+/puLpQeNqSc3qft04r7v7XGTgCtZix0GHon3
S6Ryj6ZJM6I+8j1OZsfEpI7iM+Rib0yuH7IJOl29NCJxvw21zanhzBaAmCp+LEP9guxf+5IKQao1
lDerXA7m4KJQpGqx+dtD/ydjjG2NKhsKnrDJ+qHHbrnrx2Aixe0iEcYtu4bVJsL3+IcRXBPDZgP4
VJoOCJXTdqZ1sNCUpYHCttkAkha3FBcZkKkmcw8wuwPw1o8hr3Zm6EgmQAvoheD1x/5lGUeqsX3n
XpdBvCVl6KMwULQ9sOuH2mYhntZBsLKQxZg3nItWmqkk9i84ObnxSOk65FJoWgEMKEOI3ADrS1RO
nrmF6OHYM8tDucYWW9ZMgkz8iAeWstRW+wyKBIVyV6mN5qKiQgoR8hxcfHUZtng9D5SoAAPxroxB
MOG20w/fN81mK+F4GeUhFQ3M6oYYQNTfeNQaHk27X7hoSV/VJf4wkPzU/j1sbrAsF5v0clgr/fGv
H1BgeR7S/BIbMstG12MSAS+9nN6TStjj1HodYwrbyqWOEF2FQM+MznLfu/rv6gTP7/wDh9/IkNT7
Mlj5eWAAFHtUEuWUxCrsVtagtb31Tt9Os19GGE8xOXsS+yKrBz7wuDZcEj5R+ifYmBMDTAuCW7Zr
cpU8fZX+XXn0n+hV6ePFRXmEPMTSPHPC+G1iGJH4djLblWQDXxj9CYhHX7Q/6IMnpInYvEv6zmOs
7Kb7Df2pm723jWQj0zvTAcnWgbImkRQKpQg06aQsxNbpKIruoO4jfVIFIB7c9hreyFL+hKSLXU/2
32xLjEy74Qg0kEyE7emWnc9wenzj+DMx19MwmBhTsMqManSxjAq1LxvBJPahPaHGDnG3wxFmDn6a
U90jMt8ngF+nbNyej9YrLwDR6Vfod9VSy+gmmVnybHOUeN1A0qLgx+4JTOO984dRppZwUNHYLN0I
XSdAF9eEbrmyPd2UfbSl7VmG3bOLK8uWKHupH7xTqGz7CtONwISuD9rEQuRzfvWj5rHLK/VyRxEg
JJooDnUj+3goNUe9Cpw+0/C4j9AJpIFC59dBPoDAuBirOz7yzxyew6IMR0jzYsjZlMvCP/2WDY06
jFRCCXxvO13m4KPjZY0eRvSK+gvd4DRdVg+8RmH5qRQglNbAFaSzVIARcFEOaSWUotQsycdhpBBn
YVcRE1hnePPIywgrbA4iyGBx/K0/u+5yjfm7DSChcax2BgqtKIr+aUYtpuoHf7uCKF6nUAd3jkMb
30O39wxuhT941t1eO7JNVfTPlpgD3Tf3Yp3FCFxC6o+8C6wbtqjyFtA1P8DAr4yOMIhd2Jt2phk3
Sw0wcJhizhc1g3RuDCrn2jjqx91VWeV43PG6Ro0t53wDY46eVlV0kDIM3m0WzaP2NdU6yMNV4uth
6GnwteRJi5rCc3y3yrCFJcT3BK765YDy+k44052KSmCVLz+LjxbJtCHUKyOq8RTWxtbNeSlFxEfU
tFVv//Cxg4H8h/jQgUHgW2Xv2EyMQpPxm6tAYsQW/EuUkYmy0kxrhO0Y7YJ8EScKYsPkiVSeMrdp
ilGbCK9IffCwaRULtv53huSMu9itlPjH0s4DUM3hF0Cfuesi3IB05g/DvbAITu6Jqzx6Oy2P0F91
moPTuQkgJlQPq2U0yfngyOMXkqWuE2TpG3mx+8TpshvF3YwQ/eGVKTtHztKWYUng6AipG/Rn934e
FDTtnMBkwXqsUY7EH8eNFyufnDz1ds9YfLu9vkRF/YmRaHokFUfbMjBn8lMLYAIsrzPJecrxPoyG
oMNC701DsYBLmYNk9b8Pg6OwtYEC+pS6WIPoFtehrIEaDGdrYzTc4lM0XW+iCdjfjXOV0HxF2Sul
/B+NeTcHPA6VBz6FfukxPFkpG9ixI75Pfa4w4/MvBhdHhF28rpz7ML4559cvPv4UT9BJiQ/tLw94
AUwwv9+wwJ7aspbaRf4iGz/NpRgdMeqOt1Q8lf3c5y8nSCB+CsgWxZdoftvmzFva2s6YGZDzg8yt
vsnECJgbKSuL9E5nwyPXfEu29/s0SzI4yBz+NMRP4QtYOyJgC9tpU6txLPl7W+xTBxxrW8sP8R0U
pCGzeJ0uR5xPsKV3ba88yVS4rMV0f9ar0BpSNWfDc750TkilwDcW47O0N3xMvD1CuKfh75o22XM0
RNahiI4PGmY5lZd0FQLrV/23uB60W/HcATJWKri9eErEHDhiOcpzr2dibbm6rh7qf1OSdTwkO2tq
uC+V4XpDmV8gbKCf4AhWtY7Qx3p8JkVHQOhR3KbEeyp6LS2oRTYZEBEsqcToLLX1M4+B+nMxIHRC
LeOoLMXz5sxGGhrDX9YjMSzfiFeb/bfYfpCTG+ET/o8EovcCueDEy6vv+SBXA28gvIAFU66gxVgq
AFn+xZ/vbWrmUWWB0LcEjQ7ODqhw91te1Pr2pet3JE7Uo2kyioR7Q8ZvDkvL1pXDLpa+U/Ml0jdn
/akkeA5RGzzb7YF4+gY5UNSq6SSC6WgYgM62MFKAV+2NU963sPtO/DzxwSoN4q4QkSxwTsnNOT+B
xhhCvbWzZ9bXqW0QHqCkbrP6eI4BeINxlz8rGLuW01tknfeEwDd/Yn+rr3yoUAWvb+ZUUNQ6gv4m
wqkNVIDb1tYJtIOj3RqU6T7WBcV4sMJtwaLJ2fCw9lTICiA9XC3mgRkYtKLlKK0Ei0fQCQuCz42G
SUNQkBTyRfszG6Rdv7fMonZwosSnuwhK+9716ID+Y/knC8AIfSZww+4pJfbd0mX6EfTmwFbyQ99r
Qxja6PZJ5l1Ms0RhP9wJf3xTpj33r9o8thkAFK9fDWWo3t382c1kuSqLd7wkk4pbtUpbbYD/3b3B
c64gpdgNlVX50MvpC9OOD0pSV8vxQSAchTH71PV6lkM8q1gxZ5fPlqWuc9IlD7xK9PPfT6+JukfK
vWWstvwc0q+tyKx16/Pa3IXJdYF3ozzlaVk88Gbbc24u1bkQdQQqrTvYqqu4FZVKOkankMBQvpUf
2HQ+XuVT6A618v9oF1eqLY8D+nJ9AABaQ8cKKRfooPY/dCSkbf6XAOVv/H2DcRYgsrNKfvsfvTaf
rCOGrg1qQhAaoItAaHIGAEQWUKu+O2sbZ/9C1jbNuiYovnZ78eKgBS8JJ7fU+R7hBFyJi4+8W0q1
yYSpyGcvJnRAtRGlNqUPXk5eNIUdeRQlGM6LJNt3qcHzzb32LUb6/sGPdvZ8u9/Va7l3lbc+IP1s
F0NfZcy4T9gu5/rCXfYNemdP6gjGEKf8Bs0Pqv+1pw7K5n8S7D6gxCe6j8O79Ai46iInStqHATJO
lPm8JlXlMwgBgWZp9vBESVM615fSK/Z/aSMpiOxmClH2TZMCBTHmNJJiObiQyBWRiZ5Pj6LLhEAp
g/7nMyfexcFCfqDrZf/gQ8rWnJxqpp5Kx+E84EURs4veSETkpgN4Tg4sUMiCNy+B+RUgMR4BR3N7
4YFXvhQtwfk9SUMPCjr8mDyX+eK+OUI0AHFt54Ha/IOTLX1bHVgMnHfBQ8yThHYTWqlLY5SlCpWB
4KfnRRpYhpnBEuLPbdBQ5DCNP/fovuIqvE4yV/aQJ5izxnpFkOy23P4rhMdguyM/O/PoEQ5rQDsw
b98/nOT2r9XPRwwXmu9hKeiSKxsQlr+E01YOt1Uhq93zV8cfTIHF48YhkJyven3JyXM7QfES2qfb
6zkiBMocjnWG+kussk6VPDS364I364UGJKPyAn51LNSOBBO3j4bGEWM261gFFE4IcyM8HTR1K/3p
Q38bUbmPqZ/5M4XqEdspEDQbFo6JZrgqxoi+0T0VavNe2m0raQUMTNcK4j0+Z3ww5Cr/MOZpVaUr
PzovCoGbggXz8iW+vhyOCwHZBusXvZK8OXhyjV1VuZf+qBTMDMxL6uam8InMZYc4zUEmdbKwUM2Q
VeC5MnLZORMlqs42Qa49C5+tsaXATpLUUUI9IAntR8wqE3XCLcFERepEJ2uPsi/meoSyvd3KPYLn
j7Sceppimn/vOdaWcb/F/Kt+rI0GQZqUd1kFhwr48KawFkQ5vKp4URn7xZy96x4hbyTvo0SoxZyp
K4YvcQwadivUWa4DJ/awpm0bW3RCFZuoqx2ktMG+KbX+nFWt9d1cps2JYHrCZPLQPuqHya4XWySo
rWFZilQRgFzx3orxUfGsjIjt7kVTPEqIcRGW+wgttkyeNqEUbK1u32KxIVu7dPvc+yFKUcWZEX/i
2/hgwaUSBizeuzToSvutJjM/AHqb+wfC8GsIWvAeiIRRw/MIq7Ci6h5v8iHco5/PGj8QSMVlPpsU
4JKfvus6pp+7C6o8x5b5Bo0xlNCrZaqdtNe0KqMdAEbAYBavvDhCZuR94UcXzq+Fr14rXOI0ZuHE
iazGIYp30VAJXZPtC9ZXGqf+GtZsCbCGDIFNt/buDe9H46OyKaP4Ae+cZcGhVuXmYYL67zdjy+NV
wNlDwTgQGhYL+o7Jw6uCrUMPbQ4dl10pWI2Tb2nAHkH0slhm3EmRAYUgQ3k3t3Cf4EWX4Kt61YoX
ubyB1kKbxPZEdhky8ZiulnRoe/Ug/S9zV90ricVbPTgoSi/B5RnM3tvuw7yspjnQbCXdwjMiWukz
3TUDBc01Y4g7K+j6y6lmmqOyXZdeeemRfMoF2W/G/RTwmNmXEBg1jSYOflgV/5jKkL2CMjQd0SKL
n7V5HQgpvl0tBCxOlqPMCdtayAB2ZkPt2AZP00xXa9lS6JL44tIsaCYiqT2Mwm8lnxWGSKbJHUH2
wi7VxSm+NMEJvP0W5byxkSrcma8r4glqBCZHIDsgX98eeXteLKAZLGfTDIVnYikYRggFfL3l++o3
qPui587KM+OCYEJ8N7OSsLL8M5P/vnnIjhbVKeCEytsfy9ega494pknJU432qQelZu0bt+6o4Cuy
TPEfooAsYiAf7jGVtj2QiAWZZMOLGWyVtqjZzIvYSQPsHI0XYtm83eiYxaMgoIk2pOAP/ElgocSA
3aXC2uynxauIGI2yYNvtnYuhHzZ148w5qhXFO3ACmJ+2zOkhsR5jpOasK/TYC2xmUwjw+0uH9sNB
sthYK8mcEqmCM9ftc4A/aGnrz8KKgHZbN+kjsxzP44v40j3r9RCr2j+U7MJ2MMVF7kGBPWooPZf6
wWnUEwZmGiw+qFbMEhA6xjPY4S8BhGRwkDVMOCxTP9A9HwyfKqvYdoA6gJ/GDi98DE4/QjXuCg17
qg/7n0pUjAdfV1xQijYV5WJJS8Lg0JsjrgPbIZ4SpOMuW9sJjMjE1A/H731HdTyoH1anQnWeqhWf
nBVoT9TccgyHsZj3y7dRJOgrGAxn9ehFz7CuBJ1X85BNRBqR63/jbaLyY79V7NudVBHxHAdk53UO
3RB5UyabHQTkSEzjFqYjQqpELsTWqOTwQcyStaDowHMA4XYIvDpZiBll3vYtNtzE/jtPEIDIvF2N
WptsBNovcKKtzyv61GnL18Yl4hTpaUQCSgxvrNWim0JRsvKR5hJMI3jFN9qz4XMhCQacUrcpVBtY
HIfBJ/djK7+4EIVqBT+TOPTVM6vr2PdJFawAB+nSc79IFMzxj1rx1Zssiyw2AGyVDX9lQw4vukUM
vJOovWGxlrvoqRAxSkihTx/neRHKJpG+6ARFSLM1P++Z+DM9kAnE07JTYeQDdHL26S36pqDXPhnr
OBJqmq03KbEeiTZgvPSijzreXytXPnZ9JbETB96DQMeTgjswZemYe+bUw91V3rJ8MTAc0JGStgu9
QJlUNul6d47ZzGzWKjtpsBVboobzClrCYg3T949HKdRhzS06s4GMJfzj9PxX5znF6QrrptUl1U3w
g+DdZRedlw/96+T/o+x8t40hsZxFme24se8Ywl6UJPdXyFaQcxwCnZpXZ7m5I+Vxzu5XxDul4vXF
HOozi+m4dbizDlF/ySkhEmZssWmlPlA3vqmD0SL1O1n/cv+HdH+p6V916IJBHV1ERQAdRnjAkgh+
KbwsVJvwZc5+Vi4lc359r6RDBB48mKo7Ms32qaq5BB1EXDQyX3npmMJCKXzFN/Zotg1c5JwzztPd
zNuicbM0r+9wT2+PXJj18K07upRw/xJc3YH7tDr5RZWv9KKZlTWO1qJKA4D7G8vG2JvVdmDDyiFB
P8aO5jj/1LneK5LNvJ5VBqCk9vXZn+H7gmq614mgXpHDMqAQM9f+v7Sgsw5mRYzQicRQrB5OA06g
khblAxxTND254J8fPsXgwTruz4OYyFWu/xwtFGBnx5LzZvtYgdI4xltqjWpmLkIFDRQX+ao74KM/
BCt0cxbvVqvZte5F4WK0F4+2Xj25xV8DgyVoJQf21kkk817S3aF7XerAFdokCbr2KYHTxRcMVk6A
49XfKJhUWQE3saUekg8Ndua6WkYrY+Xanxk+69NDZgmsa0NUCq7kqBfd/fW9KNkYBNQLkNYHLvws
hM/YvGFt/YyuCDROXBpeY2i9loaoTmi/YMBQD0ikAxziwQghQnVTS6X8mI5RB+pTE18y92j9r94p
pF0Q8NEEOo0BotyYtuibkMuaVmA2z9CGSs7Kfn0l/CHWB9s+97SmSs0Z+bmJNHHd0N5q78h+Z0Td
DD97A0CQjF6KVEGdw4dBbdi7e4/eVk6nEUNXJhaTRcpbdwc/85H7Jevk1PiZlKNj+8yRylnxTW0I
K379j7EF6neJnXiXFy9Vsj1MqcdvXLzJRw6/O8acRJRi/7rl99Iju9hq3IPUYaVhgPfuRi0FWSRR
gfjoc8sFfmcyXoVm4anrvSgaL3U8VL5YSu7bKKnHzt8NyNzDCHcQoTwchox2aulEpmzV/p5QKVm9
eiNBke4GdF4gaUz8QP1TlxXf5KisGI0EFellSjjXE5vnxdEvIc+kXXDw3D40HWeshin9DVU3BiJV
KZARZkuodyE1RDPVhbBLWWW1LpkkhUbTvCGzTEpkuiYOsLsdhc7kBCUVwkHUmDCborM2O715xMxG
G4Kk5F+/6uNM3jHwK13M1hi9M5nmNgMychZbQ4XBnFq3iSU9oW5AoJyA/tyPAuKj1zH0pmpZxThQ
IJlX5F5bU1jnb2cD2Rb2HcJJDezb50CMF+pWSlqNiPcNBmuxdTVQe+TSh+YULr8LISqtXe5Ljah8
CCz+8K4g5bicotIJLKDm+uaC0nQjtBCCWY9gtbPf2YlFd2AkMaHxzJq/q3jIXw9On2Mtpn9ju310
7v9qHjw2ZgxXGVFCQ2fLd3ytJkEgbHrI6jTN+kR6FHIJew7/CpYY65X/9xTwOBeJjuy6TpN3G52g
nbCwaQ00wGLXmh11XDGBpqDqGn1uAnZddnHwiNVzvTfkRF8mdU2A1BsDb4gg5TBFYAfYJdXPmrmW
HLMeCnw7ZmzrhU4/ISblLonoJoGinPzQk1Kv3LYwdOXb7pQDsPzTnaSgn/xovR3YNqEZVYihDsvz
2TvLc8ECfGukz7P7X1Q12GFrsjhm13+oZdvvpK8CF40k3g3VuaVRGUZpscTaSq1MKdGDFVvxHZyP
Vm2L/i7jcYJel+LEJqQA/keR45GCLp7oU8tAGN96IQooaJSDZA3k1TpPxyVIfyR6Isk8rxdFjNTq
K0eItv1NFjjKyZz/5+pFOimd55nxf8/jDZHAIUJ94gK0Iahn/ctyKbmAq4PqsdZkxfrR1jPCctkH
lPe3jZ8xGv5DpiXCYRhOfSsJzNmU5UShi5eDvmgFtbwoFq+G6cOmoK/+PLZ3gyOkUeZ36QqFDCq7
n/n6RdtxVBvx5pEOwIXfnpPnZpxGWJrWIIgQv7k/obr+UGb5QHw8iUk0r1SrRP5ec6WUGYKduw/T
2zu8ljQYfwsZsOykASEHZqcPYYGJLhQjVXj4y3Y3QJkmLdK+PcTC/wy1YXZsw/DjBdu2+iB35iEt
StZh+TpVJm+8h5VSm66lh8ZZC9sncnh+Lhr3ostn/CVzejp7/BcQZHqqfZ033zrLmr4QUq1FI6S3
t6t0x/xEzTLAiSiOxQTmzB1dNAWHl5ayApfC8RItRZPeO09q5FRqxoaygWC/KYkkZyYMo2IWfCXw
owYVJWQx3ArrchuSymom7mGZzuU3jV5eSNfYhSwGHuwAr0+YfalRF/ddR5Bl1bh/O+crVm+GnFmO
XoDfhB9DReB5YEXjl+c4qo1qXxuAGJo+fZ8S1aIuFh6wpuNbWalMwtK+eX5PFSL6G9FVAm8JskEG
ZbEF4IQgRtSLg58HAqz4pSpcgoRZOeIlUkdaQo+s6WyrQrL++DoGZO2H8RVvsJFhDiBLzQiiZX0U
YNGX1bO79VJaG/w59IggzipUlP2Hml3yKbe4JrigZJJV0tnQdlJhWyk4RxewW6HDezDPxvTQq9H8
zpCw1RuysP4/AWZTby/uVGKV4kl26y+I52S+WFy49er/dH4vbX7/Mb+yjqiCjZnkQ+1Xd4AtSSw9
Vlub+PNuzjIuXkJTv0hQqsBobuv7A8TgbmRVn4GkKMNG/Lm+HLRtLeiGpJzeuY+iRebRHFAag794
kg6eyb/UVbmHPsvgAnXn2svP/omfePQo9gonmmPBvhvKoef1sI0Co3ZHlTABTBqf4xWdKnvGN4kN
XUYHB+kWEd885j+7ChbK1wnomKwyVnGPouELPBt7pZ2nJ0x9urGAuuveBU/ALOPktTEC6P2oBKA9
BtHfnUJ9ZRtIRzHa9sx8Ij04Q47hoQQrTb+0Ps/kcuTDK4F2nPEsREPGNNhjrD43atViKaW2DcwU
RjkDBfDIqNgEdY0wEjWFIOJaOV/xrrGFhJyakhwLnSxQyluCbo9EKyRITiX+maM7AyB9fGIES3FQ
l5oOiVJ72U/zZK+u9Oh7NNYjfJj1EPNEaEohQYa8uOtVc8IPfBQgnTB4pAjLPk89lP74/H0i43zn
9Q1fVKeQ4NZzBVpnwd8JPQkXwwHCE2/AJFNg5XRN6NJwlRqt5kla9/w59XpPWbieFCQFgB2oHztl
TLpR6ECqsBFTzX6clr+jv/PfMN6Zllq7WQs10ESUFtZRc/+FHJyJa034Hg5OwGHDe+gPIi63WomJ
dAtcID0xE+1yd8DXw6RHcEU4vMP7hTvPDIuQjAwS/IjKzqM10eGxeBuAztvuIVxsKDsBGR6eojaq
DJmAu3JLOwEZIACF+e+gPMeAab7wt74KE/Ks7WjZJUNVFL9YW+LbrzeduaCM/GTaTbngY+lEfqSA
oM65jjPzHVymmmEqMrfhBYBfZY4t3a34y8qrzAZVI73IdaYw7JvD7HtD/AU7AXTT/+//Dv3B2u/E
W2AiRQE+dp2iocmPfRuNUznXFQu5OeuGyflB9WIubcfDRKgRMh8rlDmZ+8cRwI3vFy1ZDxfrEnva
/wti8o+LtGt9lU9Cm0zf2w5cNg9q02+GPLZ4n/nJOsBQvvIfSv9IkNbMKGmmhdtgt8OWAQFyINku
Jr31dF5rQ8eHDdJ6hjDo++X1mcPt/+K4DUB2iH0FkxinLCkh4Pwl2OgAw6sPpRHPPsTVuQhUKOXl
QqA3MSWrENUe2WdSqbKfY35yPHeGzSLfUgfEQeUe4UUfQ746AzTQwavAddkqHipanoS1E6uvtLoG
JPbXj6nbdJydfWJsg44Vhch8F9Rxy+BZjm3UMk+SQFIdA2Aquyr9jFtnqmhP8vg/jaQy3AU8CjKP
lhwqThOnxNvSqePZ+voMQrRvi0h/drpZsN87m0U7ABoH0tW5l878/Yk1b5wMYZGdh4ZU9GRd65d3
TywF/NxBWtY8O4+witVS6J3z1Mv7tI6jBRuP5CTidWzYeLAk/VxkaMMp98Ty7Eklw5Ob2IFHZAeX
Em43Oxf9v8lY08MbUDx2MCEaF71utFXqbZIqdqPz68Rs2hDEFFgOCFeUE0o+f8Dmnqf0Ho2IOdk6
WPsJ/TBbE1up2udzHAq3s3NJ/3dOy4z5r3WkZmh/1CM4A1LLiYSLJqHfLqS2iT5a5f2+GW74bZRC
+IYh0ik+Qq/OWB8HhCIzGVAv6tIkGktgsm2sMgdMWoVF/cZmsHuzfKjykanpVEzw5Egy443pX0y5
8315pf8FCvbt1quLuNDFSRV1WUnHU85WNottVuCfHbqNGqSTUJlhV5Qj5iH7hTnjlpQERXDtoIMB
FmnvKJyColzMjI+oreQWnMJfgNG2IIhlQys2pF7tWHrsw9nVM6F5bwLTrixwy+PHmGKaXj7SZ0SS
WpAjMcB7ktjkoCjHMQDTjl0860CNpBm9jcRWnf+Hf6HVkXl+ISJAcFXkZflkmfou4Blm7TXw8599
lWS8/fEtZYJUVPwk776bkvpKAbbxc6hwF6LMPVkvtJ0gg2PoN8rSGi9ep6/2/9KswY4abKd+z2Yd
wnZliC5MUlHmyv4KUi9MDellhMxwP0F0iXc1TWuJiHbrqShdsuJgDzyUybOWQOG8rLDczeNmZLja
Uoz9cAu4QtQaNAAdLk/Qglfnn8H5unfapEFpDoPsQVg7rmeCDB8AeXNZTFirTg6Zc6X/waQHxIfK
UyuO2Xa4PNy/zZ0NXBwNX2xOaiVnAg5OHu0Qs3nZx7DGJ5BIy4myu+uOmcWn6tsC3/s33haTp3Lr
+/OYgWBswxOUwqsXcHYIkaOizl/Hjb+IUgZ18p/54eabLPNDCiFUXY+XLsY9+A5ErhZVzBSwq8AK
zvpjHEBDRi2eU68r7+Tqvut+gcgHNGMRFkXBP5mPxTwzfZY95nO4Pkt2GWcsLds4ohgq3XEiLu+X
jrmcmIB7Yuc++jMCtHLPXeN1D1DUbE9F1Sfvl3Szi3Rlm1RWNuDOwzVWdHlHOhv2oc0ezuBvStsr
DstDiqF01NQPrQaODYm9WH5xJiz4H9YgWD7OCMP8l2tZr8CT5M3gjlexqi+PVwDE7ibkt9LQ0Zgf
LpMTnF+Xvw9UfTZcYynqBrI4KVZV5kP4Vi/J3cLutrQml8FZcD4D3qIjNBLQV/9N2OqeTzChPZ/Q
qchZXEoK2+u9i/M403j57eTFZce5jSpPTMMP2FSbjCEYWaPCFPxG4DtWwbpiVvegz6tF5GxgYjq4
/VAhUXPdQdab3L8zAh/M/cTqj7vbOs5sauxboimSVw2Lr9Mlk+K69U0iTDXQNYAyDZtccY7o1469
UhReYQumkF954cWdnMq+mTiAg5mm5a6lKOMZGZW9NOjsFSlQ0jkI7/xrX5Eq7cBAoytDGRn8IvY6
dxMLtfZTM/nHvFpqo1skl8/2u9391e72hbGegmBzwwCHRAasr4MqG26ILYMry66oek7+tUyicngW
Sqj+6m6sjITAPQ+rK75f+Ievw8QF1mzram6ITwc2dKq1x1518BeYqlpcx/Xx9ViXbl4clAukis1o
w/cNLS3WRPRWE/olN8Xdo7JRTSSy1B3F7TqjFVWGuwcSdlZmVPbuCJMsTkLsI38QoFsiCd+LIRhO
P23nJg91DX/RUlNcSsW9QE2dtIGvRR5hCZFnh0mdDxrZSWWVDfaDuW7HAejayxnJ8SaFNSJLU97c
+fiGqB5Jw4EPgwHjL9vE0Hfysdsm8+oCHvek7Zv8CTKtCnyFwb3ItbumTV2NTmqabyWywdL1tNqh
wlb1+ZHgh1OTdMHlSETqFt9ukYdZLKm8fk5X7phNof+/xNrwkjss6Qee74JhGdYtJMfGo3Riv5EA
KAE7a2omStdeBUvHI4BFPBR9DC5gu37mBhw30jrvLJEsmMQToAddJWty6pLH5+zeFyV5NVUqBolI
kGLY1wznjtdZ/4nL7E2i48SlIgkGdXv/6Ga+o3yv+pcflwpaCEyTGkRIFrEtN6QMqwMhiIIt6KXx
cVLv8Qprsi/lupj6DA4456U9spNhOnGV4S4C4EvNJX899OxkG7FFuAs82fofOPpml75bQ0LUA60x
TTCAVMwrCu88ukMS99blU51gOEDhg1wJiRVTBdv6BQ4ASbY4VjdKZb1FGLWvtSzAFAjYUmVJcUVA
oFRYcG5W62YgKzm75AFcYpc/xnQYMi2Jg3j3BKH21TjpVebSs+i9PUJqpD+EkDm3EpHWCuxmp2QQ
VEyc1amr33mjeqIPRt7C3tlRv2zt5YeulUUdQhtI70Bxlc6PSP1SE8kZr+GXGdm/rLwW4uMCvirm
UZG2H9LZuqp8VpySx4QHt3xVmXFgM5xVMyfHfdxufBwrmzG9RQBzEvvLKE1o3ozqmeCKgvXjOgtr
+RbwxL3mvc7kOmdwvE0hTqRPkGY6XsGvNVXkVhQ73GXa/MMmfG4NfcRYFBEIYowFnLoyCctJaTE7
oKjpDZMXqaUAXUzqH3Zfv5F6EnSDTMulkTqC2rakyOrjDEztvsvdE4IiWQGyMJOmp3jc3hcsFLYt
Ipvc2/yta5daBSrnpHSlwqYJ7tR+hCWp7VsuBQxi5KR4sCc4M3dwnUOyOo7ulSBysrdEo09YpQEJ
8pjCrrdsrGFhP2eXkTO++Thzu+aEDBb+0zT1fKS4R+3oFi/9OS9/tk2OgcnhKAyV5vNpG2YVKYXu
qhx6go9/W13kiH27KX28LZnEuHdkbjWivIRBt4TH3aKCXu/sSYYr7eOniRj4zBlSKMB6eiXEcBmw
/DDDWZMxK+o+nIWGDPxj91SfNICwUZMztZWnt4irv4FxlvxWu4h5dVdxG2xxrp0VYhjjiD+BFEdO
qKsah0E3BnClX5qEQrChrYVg7+6t+M4L4RD1FYLsfuTs/kXxPtMMndvv8P7BvCZjhcStPjlwh+7Z
H55wugQq7XeZT96wBZMsXgRDNUuh8K9Td7wpxHto1oElpZdNDBECfAGpXiOaqKW4IyIDHAytOJis
3/CZeno/cOrLx9LvKq1e0T+JSktH4GQVq/kx9wzrfxeIN4gOBRwsOlY5dMNwBUqq6LA7peDdJf36
0Gyc00SJBrDLF91asseUM5svLlzROY72H2bo7cgb8kuz4t3MG364vPwtwar1H8nV5Nvq+Y+fWACf
ltAoQ+t32TiafyTFUyBohNjcxhFRVtIp8JbHL8xOjWjTAaOot8VBpLQ0V6RqFSuAJANCzvuxSwwU
ED+HL8rGbLFvcblbBHzmxyfIMLU027etSIcFZ+XUGj8tVzGrcj7jLlvYVTzqoKddwjMEhGAwuLbI
VcKpbMtFz017clfohpx5H38blBT/AeIvwSVCYwFcmDaa3NDYjd04Jrisg/4ai33b64lt+STDhCvj
Q+pYt21p+rITbg/MIYi35CslVdJ1ZLtmE3stCeLSItmzB66eTOerKxuLMTAmJe1qbVAs0AMO855v
er/vAp1ikW6qZbSuatAreToBps9Gu//ERj4RF2hU2PIWAQHD5OB1h3wosee+EuByQPkYmdy6+X8E
ryU42x80WVshTCA2i3OGnUAbV+mt6LrQO0ZD7PeKZexBLOmf5DtkgoQD8S4nhZCjTPqGy2iTiCqS
NrqX8UBYQ86d8Ry4ih5KoEwTd3B15yyJn8ivrNVHVkxAmSM+6nc8uJJGrMi+dWa0Rvnw0PxebnoK
qNQeqLMU1zgRRgSiWOtbQB3DxPGVxvGr8B0BDeqPCW/p7252SYiGaz9M2mNywOMjkMwWJTOvTfdA
lKReROWHuZR+CsB8eQGYWbyalSPTu4Fq8oRPDcw6TKlN9EGRrRH3qVS5cfsxdyflEHos9Xde7rnn
zFhOqTCpLtpJP8yzPt/jULfwcfYaIak1MSU3ejv30Fw9J0U2JYyTuqEPXYu8pyoyvbkk/tvOTZFj
zplYyRIVhYurfLAAv3yuSGEMixX5f4OyaZfs2FGmO6RMK2g6HsdyCt136epdJjzSDknftnrId6vu
n0HK4g8tUrVFRWpFz8RwrDHCgs+4loKDwKuovwpXeWIV1OYpXPfMvyuGH+I2fXEVoBEjqb6Y2Ld3
gAPhYvUuLJSYBisyGK6IKyqrwZFgkeLtk1ddBSQgL0r44DhMkjBg4TmNX5zrXROMcfVUio+avSY/
UGqmPUb3h6NCO+VMMPgbyoGG8RMmKO7RcS2+LlbIl4jLhSWW/Rb1KtVo9twdslp/QBV+Xjic0hAi
ZdW++RSMByAVpzvuokD4WXF42qq/h1jvJcbktCIxqLhjBWE+TQX/bet1idwIIVQeuTeQCfTwXHOD
C8Jmw9kC7Oc3i3fRPmuR3M8GM53la4un0xjZvM5UJImeZqEfYJbwmg+8SmAuoJMjVSedsxu8ju9y
mwlkICHgS/fB2XCdlEXFn9paCPUpO0q7lQz/Ma3C2AXsmjhns8rhTNXPanH6/ptWkgF4+3hRPdn0
aEQf2r/n+f56zfgcJ/949/0xryfY4IJ4FST3vR0sprMZSVeBlj7/50yoE1mGdQk5xgM3bTtour7I
KRC6ErxnateBo1o0p6/O53r6+jXEI2YyUTZCJ34uM3v1b9WQ9BpoHonhq2/0KBVm9ByEfthaskhE
apLf+StGYUkvwTzgCn4U4j2cOTdq4x6xitg0YfVzvbsvFYbfAtmgwACSIiSXk9GgOqcLspa8HN1/
puvKr4joNpbhMfk98m2gpy6R8kH9zcXFfCJlyLWJZOKEFqx7YMKlfEoPHqLHbQ7cAZ1QS4iUHwRS
4gqjZ+bNRgky5bXWew9+DuYIl1qSIliNGZgedwCtDtPkQEfEV/3YTlbJjSgPyeP86tiaFGjvkoNN
51U+HYfIpgBWUEoLk4bRvGSc7uXWsXYXol/9aBpelROUz55xHxmlmw2tf1KqaMhdci6hzpFYr8Tn
kbUCK+ilPB0XiOFV6j4btgQmEcHtfk2oPqkmQ/WsP0ZrjTU3p4ZIqwA0oKEV4HfN/9JzTW9cnEig
seTFvqxjMtKjZr4C8kQ/eNheqn0NkxQ09LvxzNqYVS4vajyuXy7Oha6/dRvKvgSZr7yxHmmZDTWN
g11ludRu2m9xcSfa00kjUlJNoivtFeRm/pnbzYYw6ve6x4TSfvBD7M7M0UNtsEg6+1u3QOix6f19
unH3TwDP0cbTODRjsqhkGFMSsLBzThfEfGVsEEch7mpf56vYf4YQm3mlgyei2q0+ZzonzdJzinnZ
nDekR/6YUXTkwlAd7bOTdXzhUdVKPysA6QnboBEO8C1klLKpgIiRqj6FnZfj1BShv0eoWZzhldST
29uVpgixynTq3Aa4DygIMhrnR+89ZT+Hz4zuNukizmRunf/LERfXgrAamPag5Wt3RBq+77f/3dop
KRweyBfhHsBcbDs9kRtx1L7BbYvDlkNhcqzRSr6bRCzk0HNU3Rf9AN7oWFP8CrBiUOt+ZzOyQcIm
8bJllpOKi6ibEfbg4ETH+So8S5lw/XXab3jcSeZiaJldW5DF6cai+bda/75x9bNBS9VSo+2RrWnL
6vtIjTzqNkxAuc+hXLa+7LJ/DFkdGXPTrfw5W2eV1yQH78s7zJBWLuxnv44IsfOYubpZSRmNAuxU
c93zinnrjsTVqAgtGCvZCxQEl9/xDgKamk7EgR7qysu2zNls687EXJmfBF8P9g5d1wcCjXda2xMj
IjdDc9qfyXfMylqp/geBzyY/QET+WRQrOTqzEpNtW+TwoZCbNvWWIkqhFD4j9hCbDKKrdDvF7VL5
0wftz6eV4YFYYw1FCQfkfkROC39GyHs2oULOnkWmJdP7BCEJcP2kGZ88W7GnqF8fZHAPF096rhzU
D+u2aLVSUs4pq9FA/l/5/5CUxX8NMF68RtTHzyLVLvASE9M2lwIwFVA47m/RhJGtHeSg4sEHIavF
hLR43zOSd0MOPXZIm01QEpa6d4efcTIJF2vGqmw7Pw5Gdhra0VPl5lSVobQmAobBdz03HvSPux/7
YjAycA+rw+3SETcr+KZtoJS0574HPG1Qtbx0EcONeS9LQWNZicxbOkfHoRLTGsalWlLK5X9A8G/2
V3fIm4E9alL9Ms7iFLh1NkwcWl36rQduW1CdHYXyOV4nzPrwP0TaUlKQdGysqEPNwZ+VNyq14ufF
THrBwrggtBMkvrYUnx4sV2/l9R4TZ+oIJL6oz93CRigCo7yFQ2IpPv6fZ/hOVH+yiyUnDECtLdWf
AO0KAHOy9361YgkNZ3UAKgIe9wrA3aRZJhzORQPyHGr2Gccj9PStgAeh6JYju6NMAxJXB3yinl8C
6oCsQE4neAhiyQLPzhV5lxTz1+IgbEtx5JElBCGPFyQNGNr+OdVxoOPnX4dAynsZ2fDQ4NoLtXQj
xddsfvDWMDzEjqLqFwPNLPp77ZmE4dbBJKQvWRkZQWCJZxkJm9FndvxB0D/wW4naslwqjdIEcGgB
1KbTbZ9ch3cUZajTE7Lip2iFPgwODLtUzIAM+cKGAtFVP0O7IPFYA5HgAr59WX4ObcR03q5/iloq
4WStnWDAchj2Goj7/5x4nkLa6FW8qvzrRDEBxlp3yIVPnhwdAoTsbp1hGU4Hlbc7Jnz1rRxrzdfV
+zTy35zMuXGFEutFrOHoDZ7xDq3oJmXs0d1p8UxV4NlX2DNefDj82sDDe0ulRMfxuS8VrV/jNUj0
QE0AhEQ2/2MQHGoK+9TtjL6prbv5FGePISRzkPSuRQc86zWqyHH29IkviUewpdUDcCpTniLmlr9v
neFIP2NnVudUjBN+8Jjf0ArUPxsH06EAmKRnO1TyWrC846jSIU9WGFGJj4FkK+YVMt5v93eQY82D
/zwMmtegRaM+9yOsxF5E+aJx4R9oj03DeOVhoVAmi069sskhIC8NrkCbTQbDEOY55pr6BuRFNUMw
lq47FA0sHUNMXl61PxnWPyZh+LujuSvZDj4PXJnq3HwkxT52h9pUafvY/Jx8rrg5avMVPcrz0U78
UywIggCJjMlTHuh/Aa9SaIZ/ErSwgLuK131dqWVRVtwB1A+vLkMrZQAIIImzVMYMxI8jRFrbZQUG
Hr89g4Bva7NyTdiHNPF97GDJ43qbX9WIA9BNzblGKRd3zzVuqpvOtRaJniM5+o453vQQzsuBGaVc
EJaADqN1OKSNo+4SwV2btWaQW9036fODB08esUGXlFjGNswMbG+NC5zkQZvnijd2hmtG/nwMRH1g
xqHgycib1VFEK2sa2MDjHtH4iCyZB1qT+Q+Ozgj5ldli0XYs7qR9eIPHsr8vu7oZdFgcHaY+KK0t
VJz7RI6sPmj8jGnWHH752/pVyAMfHQvVCtkKoSlnD13joCJ4EPdZd96r8ASYOcuz2c14bbMeJ9q7
VidkfzLfxquwPcX+ddS+xeSCS1QksglgiQFSr9nlPzXH4gfYtsrUb5Hwxbnq7YJ1wk/nUC/7Dm4/
VE1UuzGm6eKCUh7UgI2UFERi69hHrlBC8UtXGWVRB0I0ItB2A3mI551TgzBrVl0VaDJD67BtDnBg
0uRh6hcyfHttfB95kutFiwHzQg56vX2hN2QbU5F020LzX2f+XgB7GqWOJq14v4/0QLYUUhBEcypr
byGQRQBX1IN4GvDsMPeQJBOR9C0p3atsqC0pYaSqjK266I3SMwOZPUWL+c16MM4S+W45PqPM15zV
0YbTez8oxaZr++aiTnmU+4V/YlyAL5WceiBSBGT+w1pZ1MWYqngGF3lESQfWSuXJV/ImN8Gkxunv
3P4MlKo1jznBXChOLEukRcnKDYd5dmZZ1fLBAgK/72hwiFjyyYQ7tNdAPmUWVjkdoxRh6iuRBHo9
5o8Oiea/vvooMvRhCq3gDkd4N2CfSERsqzzK4f/GOjwLiPQtqCG/BdrQe0RNrwDnBJuVQJJeGwFE
4A75or14Ut56QyYgng2ULkn9FuEeXVCVaJbkntaPZ15Oar4Br/+8sar17HrZ1Gwto7r3wZbvWR86
pxeDK4DDZr7BGyH8sU4ahGtsW7PUaGQpg1L8hV+z8oDGZH+GLKvP0+Nut3yL3Iv4PQ+EMTQ9YbpO
APzNiVIpmiGCM8eEZLy33G6dcN58fbkQx6Z7SO1GQLp6RbFOoTL8HbDJdjVR8DMyabHDMKKcxcrS
9raWVTHddMtBwkTVZlZul+I+9AFHqBVZ4EMIvo1EYTbcb5bPspkqb8RR9YG/AtAVYjw3F5XImN0h
ZQ8UTyW5WLzY537WtvxWy4T56Tz579golF0GA4bRSA3iemH0lG9LhW3iUg5kBX8qntJLpQQnxc0r
mpT/2FSF+t7laGWK9WiXAkzIXH8SkexDQJ5BpgrE2i/Rsyx/sQWkfkCpMIZGvDAiMuEOjlIGM/Ju
9UQ08lKGE57sbTvX/GGywuNFwZYMY0jQDSNh4CGNhXVUJ4co2K+VGsiO6W7mbHadwJu5Zc7AlGv2
/aZs2iaWXYjzoHj2S0MNiqebGBYlJ0fkfeO9I3K4FRa0GSNV+tAsHB2MDuvzrWDPGcJ7fYxU2dro
Pbqt9TSExnwvm2joOTg14exyU8PfrSV4pJ7uNQcHqiEaEpQDJ5NtnXeLC4m7z6Nc8G4djonm6xlr
xmumWVkUhatdyizYo/JfSxTtHvVitI1MpAChuFIkVA3648qbi9gvdqtncoonTNwpJ5XIoKnAQvb0
oWtB4GfIz14xigeFl5WxjYrELJ6AMSei0nDxO5Fr2s/xTdTndpzfabTB+oRv2tylvpH7n/2uiLTK
YxB0ma10niOGVFEeJlNGzcC14Eyx4P9jwAEs/XZDbP52rus4IQ4vfsZPzQnio0AC9g+ATgKcY2ug
ETCEZabpY4KxnjIDjE6Bd18RuWPemE3Sa0AM0L6IK6yvSxqQ7o6cbMylkuopthWdi7hhoG8u3ZrF
/OSjlPyyD733nAdc2mi8RKaHSpmIsNzJEOMc+Bn5Z6kzQbS8LHMBSWWrkElMWXnySHgbOEEIV2ji
pnWnXsAf8hgM+hcWuSNQs3TmfvdXG2Q7uHoDciTtGE2zwmKMTzawIizJh9r+tyG4TV4otHSk1GiY
e195YHW/x2DFo9fYfbcDWvxRR+4LY7c5uovwwn99gE6hZx/H32f0SDjjepYReJVAHmaNeJzSK10z
SdzIjYSH1QfTvmvuFeeF+VFY8Zsga0CwEHfU164XNPWJixOVp8CTY2pvQT2HVvfeS6FBGnuJotHP
ZBzDeZS87kZCdGtFOpXV5n54H8DDagMZATebJOukBPvJHVmamGz+Y+5vzV4qNZNiMxO6GVg7LAWk
exbp9Gr3xtC9szHjyW23npUcR13VUuHjd0Cx/hpSM0um048+TwgzdWFMK2ZIu6TiFywe1CMqHYjq
tZ+jc34vxu7UytwUvUR9/k0C58EbltJ1FRCazIyrT10UAiIVG1idmt23dKo8cmkkdQLUIxEet2q5
CzCP2CpUo4pnNCB/g83bueMkOLS0Gm17uVRRRwBeJrRJ4BXHQO4pU2K7wc5cIPUG6fdOGZ/oUSxh
FBtjigsogE4KQFtdCv4DkzKXdBd1fe7yJDF07bceUqrUgfuMs8KaHk07mDwtRefqYkrXx1o3R0MN
K/payKnbRxWnkH14z1fZG6lhvbXXUPJcpD7qKWkJfEXZrv4HepN+vXnex35Pam8Env5zrDqBBWkS
9gprDjbjQBb6qQtouVWxoU0Jd9eQsY5BqkeOAMN65NSsl/8IYx+AsHVLnoul4OwwPb0hVnNXNnCU
toJe6k+RxWVk1v278ENI7RzfQSxpHYZYO0X2nCYB8ZtOet8QaofYcwv6F4duYJ3LttsLBrEDhZKS
+PyXuxzwPcU4jD6c94ooXsaXfu4mS8BTSiekNW9J4Typ9C5Fm2OmVIVW6Ih/iDU3gJ6epzdW4jRd
/HBn/01qL+kRhrNAJBVmJvUwME+3zDpoGAZhSOqfIbVpEb4504dgg0IWsc0DwOgCUCj7Rbn7mvUm
OSJlR2RWhV2DVndiFN03XXbQukUUHes2kFQp96VqE+6tPv4fC5sLPojIaZCP0qze7HJAEuwrdBVY
lDnW04I3ZanRnI0/S1nmSuDeTA+ylsUifHzpkRP8cOKUXDgZ7TGjBBVkmC/6Grvu1fmbFzEmSUiT
2IzjS/Frli/I/VaIdJSscpYyu+g1p80O0D/RV+nwBEdGohA+PBtILtbMd0wB68SNMIBm1eaITg0V
2xkeAo8cgxulZDz+HMcHOFTxjtLYZ5IPxqYxN47+n0r/X3PMZ+rk93Wqf0nt8Jd+9D8ooRkqA4Ic
/XSenbO2MTffuz9g+zlt/g74GfYVpJGxeQJB+x9T+ZqhNdRfgebw9xFCd2MxN3fXxAz+lxJAkKLQ
SPA/YyqQGvgq91e6GLn95cicHc5d4FEXmfrkoG6T9RDHklJxQ881UL4Kvu7xW5wiGl/pkMf0va/4
mrCWgakRKIyfY/EHrp0FJrKRIYlb5nHq2X4Tf8bnqIBU9hAM5M1uzNxNnMg5tC4z1hnm42yIrz5t
DcSWlyYQDL6aY/T9onBthdTwEn1yZJhns6fo/YHlYqbOrlkXvsOyhbCLD/97QiJ90NoKisAPEXJW
Y6mJk5QojgEcZw2LEL0PIZqkka/oSHfKhzTgQI44ICbIDde6jnO3z0q8mRUk6x1cPkQZ2EnIDO7e
U4hrHCkLCoPa7qI3XXcWl9GGbK0Ng9z/p+EZULY5sQ18CoKFNgs2tMKgdJJwparoCMXUCwjRIyS2
vj78UsLVQ6MiC/IWdcdxqo0Md/YM+Rp7qOK90AR+AqC8nvI+k+v4/Ku44Pu523XbMm3y0jLPcLqy
/k4InCIoUQrCL4Srf0cGxETAZfUgffGyZuL0ga45hheaswy15veqarvRVxfPhl1MZcQy5BH/S8oC
0yn5zHd56nv9adqQliK17PYV4XrW6CqN2qRTtQqmSFivGS/Mtqv5Bw/mq5N37G5YOlFt6NQLMc/U
Ifn1U8Xo7asIwO80wyNV33MGjC7ISkYPJJ4P7gm7V/LQbKkqmFSxTvsQYzIIoE2zVVdsOGvjqmnT
WbeHdhFT86GcHHy5UEbZwSN7NhNi3itp7tNGSOqcjRPf0xeH+mnucAAnjEuWrW/bnE1V7fTURwFw
Wt+XvqTUs3FanEzymsH7er/Vx0czm+gig6tRLeqx67opd1QDwK1ZehRhEJvuMfqxj4lit60jkxj5
8LIPrM/cLYJTaehXaQKVLlWMqbj/m4ma7Ox0ld70vzoygvPloBiGDtpN7uDlqwADGKvp7wNx4EDP
KcmqHz7WYV1QrIXxOm0yV6jCgkva31XfER1X7lvEIpfmP2m6Ta1ze+un13to+c/eH0IAaYRFUyGw
1mWJzWC9J3gHt/2NWlBX3B/n4OEYHZYGNmv+WAS5fWM1wBPyRHfQDe3xrjUmhY6HGu+nfBeFrBqV
hBej+nrYUuKXP4dQUWumPQSF9ed3e5fMa92+L63GSGdhIfXNm0BbadTNi8w47tVjWr6zChz9KW1o
1iJ3hAzX76iD7bmIPNdL3ACPMpx9gjTHE0lx4RpnwrA/ExWKGKnrAiQVhxOpU/+nnQSCRt+mzAL0
+tDtROqxCApC0v5Ze7uoU8fa6jN+x4iLt1PjarQlkRblqwdX/DkPfL24eoti8Eih/xLnMLxtyZim
85eIzDc6bEijtyAzfNBQZoV6FEFnHUqnWjhpGnh9RQ/qhEdJgqOD4aiv31LkzffVWN76hCLYd9eu
lsUbdGr8Z8APaxlTP3+v9da4zv5o/DcCTennC78YMqkNUvq+WKMa0gs0XAcLrPnD9fG7dDYrEVFC
9w8bxvFAcuL5gls6mVz8athLShVuyiRdON2zld8RavyEPeFiXYzYe/SdI566EScpBp2UP36M5cj+
2OzbbUSut6ZrIlkgVQ0npSwocg1FO06O6ox2omx0FLAE0U7u0/xcnKXUtKTHxD7dvhpr5GSgNb2m
5v+4+uiNeNtSWi/ZFjjcqu+tgpJ5eotjhSLUCWMXBP2Z6eJ/j8Fs4zmeSwRDpoN35tVn52xCYWFG
0Ok7EbBBIXqoQ3muneypzp469o3UQ5SvG0Sxqa3ye4fBSxQ9Gd6mTwRyXpbNuBTeEfG19+bUptNV
w8A+T4gHlLxTbGah6MbmRFljnYSObbSW8lmZvRiMMvhdSAgz5zLgzdr0L46rCOopzszX8jGeQyWA
woq7uUM8f5AU0FganQ7sKIb3JHkCHffl+0F+kNcH/owapvK7teccoG78tz6sBOXyFUiQe6uFeDWl
Yj1Y6JYZ5Me2Lkbcw8JaRwHhM8idzSb9Vrqylxu4kRuwWa/vSgugM3Bb5H9oWnAFzDzNpIA+MYR7
Fr+Mvmz9N+hwHcadkICY9TadB7IPOf21DcpJ9LMwinTqPFFMrngWO4OSowVhi9NrOOBlKYl9bPuW
OHGF3UiMuXZeDS7EcOENkHdC5VbCeNK1YDDCyLZ5znM9lirmKJyZpKyULx1Vgsylpad0Y3PLFCzK
BBUG8pbNN65ehKsKiKVRGFIZNUmpfDAk6S8Ju/1K8GIXHzSRRJMR+yZHA6Jnkv/VPKnegiTVGtwd
KXFqU+fcbvbBYtuNH5WxVgVY/2yVIGrYAMjJQFRjE1kHLqppjVDEEQL6y3igeJcc/NwQocoJPOEK
giYPB6kensEFG8YD2zIPEaNxfJZK82uiR1PQeQ8s4TumKf66hvpoR02+qY9LUGcSPrPRb2chIu7t
wO9khEsxzFXp8CwGR8V4WKkcDPKEAivB5cyUlep0QjkQFLzperBwff/d7ug3MR+qT+sQxcYCI4VL
ukjDYTnpz4ZmqgGa6Uu5DyuAV3MXO9JLPRJqm3mWHPKgPYc+p0ObGFaUIGUZg4KPwGcD4dMEqYao
BjPWdZF3GJBjkJ8RNXm5qdnlG3Xwul8ljmz4F8FIqx8vCmM9jiNXFauI/qEq93hqfMs9osnoPnwV
S5lRMDhBqMPFhkZv0f8qGhXl9q4D2HwzCKXlnmvb4VdQD6eMikwKMNOLoba6tjp+J+HYBOwg0nfZ
83soJ21y8PsCw8yGEOwupyPvOlc7/UBCHXSGq0pZnozivJ8m1q1rGbVgnXYDgJ2m9stnZun8+bhY
XSR58uVHeU5Y28oNUwPl2o+4m4sgKdiIoBtdzU9iA2/kZCPRVHCEaIvqnWrd9fCv/IaQ2r0zkTAh
Pn/24CwcoXVdFvKVupyWg1nrPTl4Nug+ZqlpwHBKBKeJkLK6/MVLGaz837bVxC5cdFndoaMsbczr
SWnHEbnRw9zugGlLhEffD7Cp6Vxg3h/yMyOpnOtYF2LhhsVOt/n2Eb1fMA+UGV8fceP0DtAzBwi7
CKw3bPJmZ6t8lf0NBRNEu5GTcnQT4Rrd5Xw0laoR8LtxKAcoIg+9p1QfxhPUnk2A47+F6SBJz3p3
W3U/cT3HbGS4NO8WCaACkrK2AkkAkwz19pJZcllmTNFh3QoW0SwRUjQ6rHNjQN7qk6KUy/lBKvTK
6vQV2WCNst4OxlnViHrwKTj7NfHLyAVQI8ZfrHZ/F+jeHyoJVf8bLUnSh4RlihMGmJSucM+UZw0B
vH/cF0yidoCS7YcABHcTbJc2R0vJ+wDJ9njMBLIxFtYbT4oIagYwcfkxkkp0sWrjFC+duJR+FllJ
gKlOzG4lTEI/CzcjtawTJyt6G9faGuzNgy3w/QGgUU/AhVj7ikfi1e0OimzxDvtgffY0BX+LNCEX
LsM9t7UX0JR7hRZHkPLIfGXFExfEJQMV/uuQq84BN07KNrflBuzWVI/aN3+w/eyXNcbVEM17l5h5
nNRctF9cDV7o+TJE3VOkupLGClyal8ZIDtrEDMKa+56I06HVUIbjbXEqd3Sf+QelsOm951TanEFF
7vKytlSQHiA1C9zqZDuVyIAGG2Hbr02wEKUtYzYa1xiHiuqCihnB/CFj1DghCGpa5PzC4blWeQE0
50rHB5Qr73A1IX4MQVBNcLQJ7LP2zplwmLDxbZJyotta21hNi24c9haZhI+RsEcqOihTpVUCiEOc
824Hurx6XM9q0LVb9CP1KtUHXHJhLtNvMN2q9qj8t2LPwQ9kVQRfp95rGmz4lbnN3swEKcsq0d0i
PfnjmNOynUunlauG8dmjcYmMIvY0KEvlNnYBoeys7/I8ZrX1uUZ5mjjbrqsVrK1Tx0XLcn1mpqN+
cYQjm6gmqOJ4RhXPXsAgJolYAGXhjvuT8e+rNSWhdSLWfYy5Nwlbgmvbfj5IG+oKk0FMHWqS4ghN
8EDN9Tz8mZt57u8uZ0Ad8ep0I/FJ7GujJglEIpsCLBrDdEr+K841i0BlL6MqDhXVi6bYO63QJqfc
MzJw0ODpWJxYDly0Eec7ZGMdXfYuC79xYId4pp7ElVNXkZJiM257YVoiJtjtaFHH9vq1u2rVBCxd
mxqqsGFYhhhb2U5nD5kWMfcWGgQM7ccGEhvFbz4W/xCMX5zi0TczhBHJxdaRQzxhkP/ZPojQp271
ZTHkJhvt0oMj9bd2uMfzeucgMIApxr2jTfT5Bgq7cRw5XL/5HaTwCnCJ2tJp1MCbaJAxZrgggWip
HzaceW/n5vGDBuxrxYBGtqudKN8OVt8laLxswfIjawzBhAZjgwB8RF+6Py33CEOxdc4WMvSn+5ow
zd5DGPKHAh8Ra1MOK0ZPDJpnZJ9kIoU7V3SSjxxPiCYV2kvaTqCCxFHhaBi0HZzG6aAG9DkD+wdS
9F9oaQv9Dls/pHZ7+9IEj4tflujtzyyJhmJ88knM9Iee80E585G08VloJoSM6k0rBHiM/erL90Zs
aVT/8VTSueLKAW+zOV9uVR7kmmcGpciKl91OTtUCsr4Rmboy0bejLI5+WXm25NswVaQQvY989CpG
KdByDod2r3CqR76RuM+iBcKec8wq4s/yAfv/4K65Fa7jOfPSWmVC82dJ1AZAPhEgSqFsPB0KYfhX
f2RoUCutBu+O3WUr5gDNaH2MdCLJflWvn31hgqvOnnLM/ZuCYYK6GciZsie5Z1vwYV1oYTdWXc3v
Lm1efwfxA0NiQVTclT/Hqh7pFsvdubEj1TBUNXCAX79LcN1xidLJHMIPC/9P2Ln7aPxjI6VAObTn
0Fa7ji9XOM8iFnaXl2HANHGaFo1xJ4WfDC7GN6+Ui0BCek2Hpx4N4OyFnk5N8jxnmH98dtRgjOMb
9VX3uEkzuKNKrid6svrV9fO2YQB9VC/yl6/batXLpiQnal8Sn+tSsghfawPxbemFHCYFeZob4uaJ
arm861IbvyW27JR4Ao1AC3iNW+/DGCXz17Mz6nN5QWUTdp3/5L12MmiDqPeeY+Vh6yPtAHBxyenh
NthIWWAwggQ7VRmZAk1vud1hEuMQTpx5CAFmhAaa8psjlTPVLlXOElPUMp75mQfAw05JrcdcojA2
n/GVJcxcgnInVRHp/wmlzsJMuIWGxLB3NT7dFN335SQ4u0F+hyV9cpr6ZKVeeUOFoubFOaKKDQOO
uHD5PUzWFZ5zZRliIA/nbmoeGHfvJ8OdhO5lsV9TSZdvA0ze9YSAKcq15lvUPggd9B1XxAOlqgWO
JZW2NlqEkbhbMN19Ns7G3AHLnBgmat5YFxVYAi+9FLiMNY1PgkZLsYYBe/HrC4UEM4STJkFv9sze
sU6Aq+Jb6Fh+sTIyG0uv1FV7ERXTuNm8C9+RskWTpqAFX+o+jqkXPPAZhI2ZS8fUskEik1NP297Z
2oiSADhIRYomjvUckptYeF5Cg4UwsNHxwLQaUPnhmkVt0Kwcoeb5TiHPCdKnqaio1vNha4sDX3Ku
mAI3kPKMkyDDrVkBzLkM09McbroYE+ZIJLof8I/2rKHjknfv94n4ibdC5M8YJJ8Zr06sf3uoda0d
Y2wB12LhQcZSRIhaR9xSARwnAk/S9EtxGh094zorBTYT0KoVvEzoexMLZBRGwQp3i7o87RvqYJ3W
LEr+oDOBOqp0LYwCIU3DXGfGCeJqnqphHHimw4dqGeuZGE7NtbApHhXxqLUDKaC1p7Ztc73Rd30Y
VB7Uo6G/D/q3bDOJsrz2fdjQW7pdpy0wifXF6ZpZQi7zmYx9jveDkPM/LHaizjOR4drd2Jkt3RT9
w/WXT91RlaB2lW4HwMjTeFVroOCfpkTOg1it25I9IMIgt4CkRKjViicvOeLbFgtdHLWA8EHYh1Hi
JXELoak0JLg+53u+kmE1+4Nh/FaTJc6jiBWtXtJUjK4Q3hkvLHP/M0Sw+Ez6X8OujyAYtSVmp6cE
v2Z92t8Nh1cBSMXgHPbkDrXTMO9S+ku6M+MjAWTdD2iExgnWC1CI+GJbEkbBLOhmxPZZIJ92Q2mP
s5I4no9MzjGff5G8ODisHnm9U/CZvS9r7wTL2AdHcODAPbiqBsDshDQO8pWPpZBvHAXHl2kC4UDo
rxrfSfmI2IqHsmCoXXFNPtpLk9gue+1j8C7JIBKhTKYc/Rh+cgoxVG/7bDdVpt8MmbCpH7XzgHJC
Spt2kXz58kVDrOy7HRJLnlJz4oFBXhAbbQ3oGE9PK8bkhTX/LufTm/p+U54WnGYM/vDiU16mVMDV
S/AFBnCOwGFrKxLCv8/IbdQ5z4GuBbPQst99AyhLzggQ8oc9MZNZhlU3BXkfVzDA9ZrlbSFjSLPP
F2a3moqTp4XKax9YLHH4gPHO+iKeYtQ1JNX9qorVvYMLgnK71V6a+fIlLMVlzh8CdyMW25vOZ7oI
3+pcl4OvylA5IhQVlf34aK7H0ppRsroIAnQAvUS5+qEVgQM4hKI8CY+4ewlkhFAMLsyXXLb/jRRo
HKrhTnFh6INVWf0Ou8+NuMIEAr8VmAH1oN4atV/x3fsBxuqdXlNt7Trqt+z+SXKxi+HOpnfM4Idp
DonICe/EyKEwGSQ0bja5lRQkqrwE6gtg+iFKHSA9+bTU0bPVnoxihFmbP0QDwB6Odu5hTa9iSg+f
ToVFVREerVBrw3ZydUeY8JeLwmPyGdz6tDR5EKkI4WxMEZ5aeTOKb4Fk0F76Ty7hgVcoKIcZVznt
pqKQcP7NMR/tx8oqYSsi8m0QXM0ByC6I6ox9UbpORU6b43ncup5MJnIuMDYo0U+BLldgXPXrsl+L
08iUyMpbvP5KJup+mGtYRT263ekmNVmX/yhTvBJTv/789K3mjXwX8P4z91PgZkID6h1BN1LE7aG7
CUtpswqRuk4Sy+0RpOv195cnRTE15Lf4nO5jJmFrbwF27lhxd8ynRYbc+dJpSAxVl4qX8Wb21ZUD
Lh8LBz4e4dH03eTCWRGsQpBATNo0SBLd3dkdKyZqdyzfCnBc+ovv0UwUUc6jZcDoBlOfzcIHe6dR
eFYtCencXvRUAGzWXdKQv1iOriJtmFkmmdYCyYLXB1ntnF7t3IbrRb/npROxGmka0X/AxFdcUTSL
nLNCM4bQ3I9SPozS/B1k07wH414FLuqLVa+C0Txd8jZoo+nGp6gTKic/Ih0G8LKOkffpb84uMAVV
SsQCyy6+ycrIpFDCrKsA+UuLMrb4zJT2z7STFYioz9kRf2HXE3p3kxDaQp3H6h3AZDDuNTpbR21g
yrqUI49y4Ud3YnRevfR5N6PekCy61XcJiHY2Ll4kKvHzhSQez0+llYyvrzdas5b8v27i697Ayl0+
I/k904HRb32UJCTTuIS8ZgMY9s/4+66QX9ZYj30prPY0g4IsHc0R4YtICvXist1J7fqoXtrB7/D8
ybOSAPgEIcAThfupMVpgeDzxSQklek7QOIynGJ+GgMqMWfEMrdkBD6hlvxKHW0JgZsZKQFkSRCAz
7nnl3x9JaBFD4zmY8Ah0YVHMY/QbIPi04lQB5pk0GgiIxRKgtORHfbBelgGI28sv6uYrxCzefsKA
EbF9ozhyeh20Vgk/eP+NGOYZN3f05JJsYUHUo/KplbNbWxfAa9X7Umg/gmUbWuxLX3wGKIiYUndx
3Q3oaatFBK5WFBAsi+anxG6EbMEe3d23rbS29WvksvU15xybDHDe+xdHbGEzBlc80Nl6lel0B68y
fvIozwljzj38rOatHOpfrmtCDPje8vJ6YKS5y+6FD2GrxlyAy1rMG/nnAEmMRbRnNcOHVAGvZo/6
QR1FZnHfyY6QzMxZbU9qLahhgzzKfRHTNfZ/wDOyIB9cg7190rPz6ycfPRxbrBQ8U9rQYB0vvo4+
wcRc+dJ1FG5dSjk6KJ0FrX8ioNAKvw7COZ6BAf9R7RXDgdh/q+EbsC1rLkhtMDSo09u7uZGNb1PC
a6lPMTBX/z6dZpZksLb8T8ZRUlShg/fXyPU/RxnU8SapcQJzmkEwOBIGmIpSS1NC/JzJHflUQSNr
wu4MbHOC2ZoMObNFsmMEqhwjCelogHLCSDyjBNlLUCBkmLd3X9eo3YuHiOz+snT1Pmj3Qjp5KG3i
9aGnFbqp6nVg1YOk2HCHUVkmeoY4imUFmWF8EB8yhjmyJLVxH49eZxy71iJTTIyp1mSX2HyUOHhs
P/jhZfdtwBsULuJCkeoCrfDwlSA+fz64WP3oJh2RmKXRYdOJ/hkD0LJiZ+sbbTAy41chZZtWd+fs
zPQ6lRw5me3/bhx59l9JbsimKvFbFkbQ4hj8zd4B/exHgW3zcrjGFtqOEpper0cQO6GI+ADTYdlj
PvbC7MwJA2PrGJTr0JJzjalZ0nPKwrSkn5SUxnUlWKyDJVjyjtEp8/mwfzA6M34I9SlSNsW7F6DH
UhSJpmlFVFTqYFHmpqn16iVZVpxbFZQSWN5eXoQY8XvVbCURTu3lOWCV9pRTsbAzQyORiu3biP0i
FK2AJwEO07cnRtMS9ZzdYKLnKEgrhwNcn2EAWFNwFkk9/IIO58BFZi32ZXGs/l8QaRDnKsC8HrCb
Ende9K+xaTWyEMKvHO/Guf4r+i8ZQ63+nskxbcxvCv+KWLDj/Mf6CvwXFAaNWCiq3BTscbVv4q5C
6KeDDydQYZ90YE2lzE3yseIpXSI2wY3NMdW5NMcLrmtAYpS7ArH7gtVKc9dJi9VlF9SgobMu4UW+
I0QCwSEGmzg9P2hxuI1KzbsLSEeKZsMxxGO447qv4iM7ERHBspNNWN6y+uTs3M9CfpV/h10hmZUG
gk7h3HtgzcWzf1Lik9nku5IHiMUiWst9fduHcPoG2NeSKRwUleq8t1PBchfsJXeMHsUCtdoW7nTD
B0BKHesaXxVCe4K5Bova3LLk37heavRoa/Wb8vDqRQ3958KzWnsI3WQDHDPQji/5KsOVDq2qZYzx
sBLlzfyhy2W1Wsg18/d5fIqO7GxPk+PPgCly6L6HO4EU6cCS+0nBcrbyl4rh0On63DqDyUuQaC0o
/nWtVirD3V9Njk/ZqR4V3hVRi32ePAu3+WXxJACDIixWO21n+63ZapsHznmnYz46U9PQs4CSdCEb
0TUirLtVlR7oypu5W5Ok56JQ0YMN3qTKvb/8MKlqrN1SUvCvC8D3LnyxFNFX1hHC+P0KcVQo7SM+
QqKcKUQnAe1l6CEa/gGAi/1eu1vdCkGPpmN1YstJFDK/xV7mwDNcCmx2pmsPa8kXfn5kTVdQbThB
4NuBQQ2IukAcI9OE1xNR/o1mFe4wG2zy217A+MSpZl/zRQzqr0Nwq3pY4QaT+MVCxoM1LWwUpoAw
OB4ECPoBbbMD/QjZyjhrZgPIVKCHsYkMGqYNnCGAevQimhZCTJWFiAd7AXcx8MP9DQLWIWj8docg
HLHX/LtsV9ONYhaw55dyAR7aAx4pf2Q6MWGCBAAFKlQod+fMEBYfy/ehYxbnSfkB9401MwX1JJmf
ukU86UZq0cYtC34KhQff21OagnzoNDLWIYWhGZzbUmxhtAgi3QKH5rBffDwIxcljWO+L2HYgU4wc
lyBEWtBycP3xWh859Y/3JI0/ICa2TbtoLAuz7zIdorfjjjlihA37aWe17MjageChSECDz41ppmRP
+N+YlbNOSP+e2XC3cU8YQ586hJ6kbSFeR4pqzE26qLhXrDYXdVMqXk2BaiGQ5u5XAPrWG9tkAk+I
MapjDwkj2FPcDcub0AwJEwaiw606R0BW4zJXgp0YkWTLWIlXpVCRQJy+89aDmx+m/O+FQMpdCYk7
h5ppqbJah2manJqV4Go6SZkivKC0s+ImyEmtRr606+RSEgV/ywLwRA6dAKUvq//0dgmB5CBTGJZs
WFU/KOcjfpaoKitLFtDuON76V1ENfQ7U/6q8hdIODWOJTvPat5FBBLndKHxhO16JCmNkvoIusE08
6nmRGpBi2bcfPrrCCJ+hIU8qEG6C/1UDfZiW7rrYxFTCFjFG1UN3ETrZf7CVy9VFIzPCK05fgUou
8yFkpyKaowsx48I3KzCL9QXtHpZt8KHau0G4vFWxWJszNZjb/xhcrZl0gARyvIg1B+M0CWOsn7ic
ol+FAktaKTCC8tvi8NbkUVhMLnrFrONJXApUCzj5cLxJiZqBYphPb4z8jUPdPsY/0ShjUKRS4I/C
uFtUGJ3NpaoBW1Z/HebZqv/dTJXL3lagF+9Hz+ymKTMrPmLCpm9yei9WbM9XN+EQH8oTHzeYa5kK
7SWWKGTgvjJFGeID02mgujX1yPTM5LTxfVFJl4T3jPSYdg9bVtCAOJi6SXIm3T2zrKS0hkffBu6J
1dW6vSh81nxwOb5iI9L7KcKil8fC+O1vyAPWgSImRAHh/YRY+QEAojICqwkqKb5zEbJZ5hUmwpS3
iK2o8DTpvaotFMyKRXs16o8bTSK1d9e6q8rXRvEXKa3g9vB5IHus04PWdggFwa32c77spQqhBhaw
zrRhlpwyGDbrbGvS3dPT4OX/quMbTj1d05pjSVbp3M1LFBfktBcNCnf1Hl1aqboJt6NecY9/EU2t
j+cfHwVD0ebjpSBiDB1ODC0nN3jhZRDs+ejTdtS8MkF3r8l6x3UE9ANXg+R3u6qLmKADSrD/Pn7v
/xQRqiOPkbPP7+qlX+olmDSKFb8RSnYj3KAu5WhNBUYW9PNKF9N5aDRXQM2RhVsYal4vUHv2CwAh
jTfAPf6SpqvJhmvWakC9Lz0XYX8roVZiVIorAqZFjMlTBVo14WQgZeDKGn10FVGigSBz9yHwTKs3
NbvU7jLNCq/QoFrmZL/ritUTn2XaWBdXHq8c0i/rdjPN0C43dS3yJFYuQ9VN0q5C0ZL9bejVgNgU
qPHO0eKsfvB7/AJacTaAJ8RhMPKT2kE+A6e0Oo1EScvG5mV0ijWsTwJITZ7clNtOY3o9rRloKLlv
GeLlrrUZqiJcx0nNo/QFxRlqasD4qsOL81KY1iJaSlWtHJokVovrXWIU2wBBsiFIQs8BFrblgUX/
rLbJj8yADyPw99qcK0Jkr7QSdNwlCpS2shGDdmLCOhqF+edoLoiIowNL1dcVop+bs5I0R/zxbCz4
+bezn12wzSdDro5AOPskwJwzmiTyNV6vYyZmuVOzioT6znEsX5z6fL/S2glaVTxven8ytuIuBMBU
XKWRMNHV2kw8n/dv4JI71UGOY9IPbg9D8u9BURZ502g7HlRLvN98lxkIeEoQe6EpOv+6CBLP92AV
BFvir3ibp6SAfEAQ2ETv5BJqpadyaaLP5NbostWmnhflRYenjwgHQh2jYpRacg41zKGv8ig710hT
YqKdXOwDxJOPilMfnpSW23Jx1mSUcnHfVx86OmnrZ5AbTkHgrlmvRW3hUsISIubiIfPafil9HLxQ
Apg8dmiOWixk6PeSO2WCNA0AOEXTLLRujPOY5UFh8L7AgZuVR2FlH8fd8naqi3l7Hb7VPNzGar2w
3z3nxdyicC26208FAIZBmzhyjXihfRnK6JKS/hBL4OZpGBU7r4moE4SOlTLxq0z1S9aKeu44AH4P
TTvOC2Af6SLhQYU4dDdWZLwygjj7tjW3XE3s+JZnbxH6HT5il3UO4B5XAxr7aImEEWAG9t3ZpGqR
9y74i8Sj49kABfnS6IlG1ZLTsm/KteRD1NXlOaPhJ9pvVaTD24ZBFohuz4CFJQRL0ur1hp9fe9BZ
JCU+voE8caoCVacxlqRMEchaTfq/XF8vK5BBsymynz2kcBVc2nvtlX6b2qjnNyVN+69WyQIRDpRk
kSvNDV/q4R7VG/KuQVGw5331VbXaYobi+hDLAJmQ++zpiXXGB4Z5h8myZ+KILk0LDrP2A9qDThHf
HBetP7i9KbEwKSCgJykec4fgArpkF9D2ObMMWxRMCFRZWatirU1fnM8ptITTfA8iL0roUPBzrl4p
TYNUc44Wau/CJoxUPv2WnKx5sGMcNfEK8PPgyCJ4WohQWHsg9RCe2jvo5ujJmHTaOFYOEVe++a9c
ylpCsYweFHz1fzFV7low8a67ZDP8YdHpL9ri76koVukJNMc+ymjVWlhh89ROS2VCVf4vUWJpRk5h
pj2AjZKlpIgjAzubEY4syW5Ip4wK+UrlDfGea0l9/eE35USrcKa/mXdILfRfazOWZEkEdYxkB44C
BgoGtE3VufTSCBT8OfZ4oibZx7LItf0QWiY1J/CnlQUto/YBDKbYkh/13ZNFfS8j/xFC49U/BU5H
1ExC89duAcr3dOkXzdqFmBOpruvgs5EBFBWjD8QP3Fek3aZx5YVZAhI3hSiR7QhL3vD928RmoGqn
E9eUgFt3DAGhgHsNEiVCXEeSdFv3Jm9V6qCyTFYFD5TWMqcmp63ncidMti35hMWqiOJaMnUt2LTm
zDWd+gfMGtSgwo5MRyIGPuqLjmMKeOcs3Y8A+3WwKWpTsMf5anya9AEV3q4Ci5NUIPETUdq9o8xP
+uNh4R0sj0IgM9oQ5vLoImaxNZL1+E6GrE3GVNR0ibySPUS9y4/wYIjxR6iBak+IKQz/Z1dK0F0i
x5C70AqySP0RT8yR01jB1Fmnqhe+LagM3GVp800s/zyYXDvRmJUe9lTDgTknPSzgwr80mJ6TA5W7
CBsOV/gFanfa2wQk3aOMYmWcYF9mU85GZRIJqVvUArTsTPWujoD8ODXkXP+Mc0ndGLTEF2q6f1JZ
Lb5Q1QbyvLEVqcg+aeW0J/qrCVLf2AsLBv1zKsW3EHIHRiH4CXyXxjMBgmZZhSYJFeaikJ9Eu9Dk
2QpyRID7S/HvNtT7qnyzfRS6CZN0LwWpdmwSoGMVJ0V1yOFD6jzAhywoZbT/fzLAkzK1FTTOJF2R
XvD1cXswShg55M0HOCs7k9zvJincvBxY7Fi/yKT1tn5zowWCIcCs8hfNKCcknBvKKn0b1EQ/Z8qv
y3izH7ifkeIsJJZGJp+0rgOQpMBtEI2/BmKlltBOducjCO8pTUvykkOWoL6sUcl6IEHuB1GDVWK4
xPf8lOOHUhFGdjm7m4KV6JW4B2kAC+IhefAZ3/Iw18cSLssdZR/PBLSjStGnnhgL7SD5v6hKNhsv
cPH5+ebawyRGqeEJy27nec1B0P6MrOPIPoWJyS3aefzLfaJHJ9T+++MshtRpmg+dyHdkmnBmNvtF
1yD+FFUBiKVCGuOwdoBGmCSV1tyY4Zbf4kbfADfFzCWhP0x217VQaav3XiWmyC1qlKDlofVtVUy/
6dv5XD5XOiB1z6wA9OhIa5EM/Ml9q8Vge1uAcKmeRq7u/P59GrsKWqM4BXGm4ELAzK5ADJgXK2fb
MEXv+XaB8ChmjCeFHeFAbC9H2xsfsqauwbcKOFpRO4mfncQ5dmBWmGzUxSAm0Lu3VN/SpouyMfcp
x0R4Q0r9yCrwaGzgI9obJgF/E7bCPYX0agDiqEPoG/+7MnIRIQSXOOhINlBNCkMW0IIr2JM1fUhS
iWy0z33SfWMt1JJbPiaOGzSJ2sZNfSL7BeBgiNCnN7T6KIr2uMx4fiw7yi7HSisvQgRqN+vvWf7S
GhZtzkbfpKCWgq9o37COEPPFS7qMhD9FFz1rhrpsgUCDFSKlPD52y/nlaR+4NbyeEM8p0pHpvjt5
2utAboU/6wzqAUBR2Uu4MNsHwGddh5L/NeXn2D3QwsbgJ1Pg870j0ZKrmTbiL6lSXYDUaGl+kFv+
p4OW1AXfxBmzxpl8Mf4N8EtwdL+dEQ0TGuRto1CMhEoFKnLYVZwsmP+EWFBEcTzqiaVkr+pPmmHp
zRCKzZNOQLG3b0mdY1MpJNf0DLh5J0mbfBz3Xu6UVIVnpJR3C/1wzHceSme8rXg+2oE/PI0mePqK
AysslfxzgabkerF8AdUp7M584hzFu5NQP5qrt+PP6oDqdX7BCqEDnOBaaVU6ZwSODJGv8xUrK60c
x5N51mXp1fBSnZCssMMW/ciLu+jNIPJbeZDjKalXNeRzTNEG9iJxsevQEiwpZnTffyxK8NY8Hsvg
9k6Bgrw2SkGe0yhx4FwUVpCVaXOoHvkZEr3HTzlCj0BkLzhC/mSavigWbkKBe1HRQX7mDqDL3Wg6
Kylk1Kql2WSSPzfB22F1/YxsCz9O4hOxrkrYthKywzmjRxHDA/g2fWVVLkkXwlmeW+l6Lgd+hiWM
MWG08TLPlLz3PiAjK89hkHw6CilzirOJULX8V9LdJ443KAlwiXq554XZWnYSALzwKfzn3vxeoIZt
8nrQX+CKYDWUHEW+Bqj0EPZz5GpJC4AQmCaL/2/keNmUBjNwu1Ddk2dIKADGX6nFBd7X8fPNZ8F0
WWXe9Z0D1Y+RKLQf6hy5PY2Sqx3XIFZqwjT10m0fFLjrGkfm1XpbiFoSyeK/LgXRUojCCATnNuhw
Hc8DunfEDyKCXtIqDVeQoFaE7ARASl6vthgUmaYSFfTaWJzaE9O+kmSmoJN47Tm3HbWFeg6dzJno
i2czfCq20eHqbBb006QAany/YzzxX4IKOxPqK42xgz+TFTs4a9YvHhxw/ri9lSgkALO/g+EDqn8c
tKLhMROUmswWrwBUPtuaU97Af0bIHpydMneqC+CZvkjH74XDapSqyUb88z086FyUQPhq15HkIFNm
ylWppAlFphSsMNy6nDTTa4wKvWh/x9qq4MDfV//gCHPyuTTWMDYiBfR696k/QUdxsemxeuJ7VFI9
vTvDKlWKO8IshSnhze4Veu7XNM4cbU7DRlvp2/GW0xrGvfO7TS6UiWMEFcBk04nz4ou+pBlTK+sZ
JR6gPkBQsNpJ6/j8PC5xdLkzEBk6mKs9ANNb5JdbaPd1aHeoxg28Cj0TMl/Bk3R2DVt2WqZX3KpF
JhlSZdAiX+fCBC0N48yJJfUzSVdso6Xoxm62FosgsQ8YNPm2szLyZ/BENQvFMyqma06v4Z47G6Wz
jpUQFDx6JbxKGbmr70CdUsjIsNF4NZNbx6kaSjaPxbKvM9QnxYOfRS8lVZZe5xyCNSN6Lr8GeYXG
zfwTlE+6Y3/omQokV9ARbMuGe9Hn56IdUwm7EydOo/fRLiwQu/WQA7kHo8A/IPTBnqPYr+9ur6Fr
ftlLao8dvanlp3iORBoejod5a/PADsSirfQi3Xv17z02wccgQhFcBf7obzWqcaV3BKVlY3/WTdJb
c98w+yONvdgvPt6h3br7zb1Q8/Ep7LzsW5aAp19ItKuZjt76uN5Gi/ldigbp9K4inavZM1mk8Eg8
4lCFCJW/kUWEUBwtEt6qB1P/THOWE8lK3lwVpTdQiW9ApvKDdcE2mGajgPWy5sDuLuBCC/81N/0j
TMBGJrkbGgpSfpezeA5cfKL+ePIZV9T/SBxW9Eh+XX8ZuVgVqIS6C1ZcONLAzlnU5Pz+hylbh09D
7/p1pgAdW3KfvC7S/O7wXtqJGpieTwzmDjpGagw2TmK/ViziH6zJ7YutTdP/HX5L+Vlgv4QhnD1j
eLJ90uGjmFBJwzskuixCg5Lc/fZsoAZ5eYADfVo5hJQL3ofXruPtk7tfL/IEDMO5EFovsS+yGwrq
BYdmq9+3PVhe1TmhopSdX0uLW/4pkhFl3nltgr4RSAYb+Kkf7EVykdP3hHhbOPwkHzUsnEIWbPtN
ZmcxkM/HAwgVbRx7WFdy/aGOHq5pq0n9r8+uO0jb+WiBy5+Zj/LGDnXnlxXOYfQHau/syz+WyO2n
pra2t7MFjDM+m+iwRo9+GMlin6ntRNImI7TVVykTdvOLEF6xA8P86YXHZmWGCfF9Qsx4Ve9Y2nTY
PKy4F1nlcm9Ccbu+EzZX+kQoGzYvlId7a95lTiRjjHFTrAs73MYjWoWvyr1UdtM/c6KbSFVqLBne
RbBsbl5Nryk7Y0SfhUOH6/MZuZEl4oCNPEFlNjD1V7xrvNHkBVIOeeQikHs6rXok+oeigANySYQn
4D1Lt2MnKjYiq79xtj0ljnvyW2uRnTuR5hR2sTYnioLmnfY8nuBdoXOnBYp2O3V06r0+BJt/zR4o
iMAfHobTKdzSd7sAj5MQdtjRzOHCDJUh+9q3Ono7crRKGqmeQNA/VZj1UawOBOTj4TzGwjUAQpCb
4H0qZd+se+c8dUOAF2WaCR6M5Y34WdnXVrzYuKeqnhrr/Geyv6yTLvLx8/+X1ekIh3bh/RQovwg9
/iBkiXcvG/EIPsw4o68BZ+Itpm5r5cxZVokkvd5tMhGvL/BeJm6Nw3U8XIsL1ip9gEHVmGIICTXd
uVoUuBOS3nMnD/msWIDqrJixwV8T8f7yMWuOvYhioyEeaDxn17IZXb0sbbWCGUpoZbf/5DruLaa3
hupRhCKX0K+lBDDg6P+QeFf6960CJ2b8azlWihQSeyLmk9SuOwd45kK3UG7MzsjqK34/wngqEUjQ
PL7D5usgsmeKiILlJqWz2xKnnQnI74EPJQr5UbJrKLKityJSIayntzhNvo7dCJuLA97KZaJP0wZA
1KrMfZjYcyR3m3udDWWtN+aFzV8KwQxp1t0+45OChoGv5rVCJcbaK017H3th8UnJDhnBjYG8WLeJ
Kz9JUgid0CBXGPAiif4zmL9FDEvCiltR9bXlNN1kTs7KD+k7aNmerlzKvAjYPc7hkTjtWa8kQq56
NQrLjkfVLn2+gKKj3oYSzM/uOsTNs61ZjHMd/tIZOCzYKfSo2wPe00ILln7AXU4wUiV5bt18WRw5
EwhpgZAbhvyQlePSRHtVav+1b5DDtRZ28UjT4QDa9sse5LpJbWwVcRhdhFpXyB3S4dexuD4xXtkl
m6plhW+jSpYxUwewyJRLOvyUFRsZFaE0EWsRW/HrmD/kCgp98/RVEmoOHrqN1Y5ybaoV6BBQPWYE
cCzPRFll7Q4kDoBFAk6HtgSj2Cwc+fPP0TYA7v8QM5NAuc1yxkD6PTOx6oRDIqolMP5L0PMSbD7n
7DuDbf6L9HOLkLQOJvPHoHqBM6OFAcVaGgXeXAPHDc0smIRYuSJzbkK/IF3vbAvnjRxmb6KW8DlM
CXxYOx11thvRSQj3Kl3TeS0/GfY7vpZwiWvRHccUktUym9Z+r/bDoT3puzDrfrwa31cTeK84/OOZ
6paTZj3Eotu2icBQmb7lHgxWh0rS9ex7JS36sollRUlo2TgNGpMLt+NuwKo0b/sEx+70tEovDOlF
1kffBn+EkLROlO/ibV/q/uFXvwIzt2QYHn4C3PhTmmUjX5txl2cY+sr01ZxwImDHuqUiL+S+w1OJ
+6VCbZpOTRu5F70fyeTq6cfXs0BagE785ZGm3DK7OuIlWG2EmOC4pdHyyX7uaoos1Gd6L0ZaFhFD
cweyunr27fjv1MxSHoLmTyv31PyQhfEoDrUiSnyRF3AqzW4djZfrsqhfHUQWeuiy2pdDRSUtYuhD
XqJLHTNLgilX+KoyN+kk4gL7WpcSJ9yS419yGaig5l3YOx+p9DEogG/eKvrbYekIX9eCFbJX4aJy
SrPipy2qL8w/FgHPJknjA80MiW34t/N9RcehHqqANxZgbzZTKDumS9VjHqpNKmbtd/xhgxOqflkH
U1ET0DY0rv5VxocmRBKVB77wa+fu/6JY/R0CJ4YcIXenzYcs+X1A4M9v13z5dS5m38bITpDnFGF6
nTXjXaRPBnYylR3CaFiAp15juXu5LkCDchsqhop68ulwLIyIyKZpqEEO4IsShQvcRR98O1ZQ4rNQ
l6unvTew4VzNoQgCJV67WBEp0+edrzF7LLjYAiaHx3pk4HNJTLhdUlSYY0VW5HcsNlXewjTgXeAi
kSCQ69Z8WlI2fGvL2ngR6UuNMy4ztjZSiTUVYoiHlBBkbg4D0kpHn0O1lcWUy8UT15s/q1c+Lxny
jNtmdoCQgHPp2uqBY2QXJAwNGWInsx3rPaCNzd9X06HBkBfuqbaj7J7pNCrYVVfbe2IzPfFqh2lM
150vvSA2bSmYAmZ3i6+7hbuDIguHsmEiitesrZgH40CtJF9/+cacHW0eHdOvGZWpWU4gDTykOAcV
v9L6M6meN6ZL4j5oUJuMfnr7WdQTRSHQ3e22Z5bgVsUgy56vmnfc7sKv8o7Q200t8+9g6Nq3/hS+
Lm1zpT4K49OzrdjSfF7AOpuw9iugUD9XPSNbnFmeKk2Bwx4zYh3Q13fipeUvnlFLtB1nc8HUatXC
pjbE91gPvhwxmZX9NVg83scpLBazlQVn5taWqGKrqggEHbPiMdHRCyHAmwgVwV3dcpF+mW50w9zQ
K7OUG6wnA2EuH7H23OA+RgoVbfs2F0d2X5MTtN3AjTBqM7imuPB5iREe0XLfcXWToR9837Im6tap
1To4KhxljSmJhDn4aqrqNCWt1ZAxsZvbkZo5s7AQCyia+YsDIbASYjgTJ/NzLIFfuBVXS4W0YJm5
SAh+2luui5dgoPgZc5r5oWdoZ1W5vRdtPE3Dmn2Tlkz8/Vxo8faXEXMPw5ubtCSCab0oQainEyfI
7tMFHcFFBVJTfKfxFTj4Z5d5e+ALSe1GTZ7Yb9tlrHNcohtbUn9z4ker+0lgo1WsYdii+sysLOCu
rUsk7xUDhKRhpP1QmmTJ2x0CCx6b6LggE1kcXYfgA7V8tQgQn/rYCctI+2TkuNlV+yA0knwmH3Dh
JYs2bipNDLGjwvxSp5t5+ZzlFGFv3lmllNoF+gQQAIrWTBbvir5n8vnoVgXQOAobegBiz/Xkdz+m
RTMJNrkePjZWzznuIKVQAcoNnej62UsrcXtNrRmqLaQ2UZga64sgiqROAVflU17VGIaaLNv9o8DD
w07clT5VXgnZqpzvezM/ybWiKSrNva7m/eXycLYUYIdzx5A4c7GMW8sUsGsn6qlotYFPrx5SsIdL
/imMnstRnU44ujIVARQANbqG08ENKwlbDyF8ECXG+UKqwHVNpfHeLzFXrn+NQV1yx8aCrx/ZIbSh
R7i13WaTeaUMskeaUV+5SCrSaCZYYusxdxP2wW1aVr7Sfad2nEHWnHdLtRrOFefYai/ZnZuSEW8M
UoxXsi2FpDAvx+SMvS1ntwoy8PCRNS1Qi+aPOrhseU8ZvSOyPR8eJI1KEKGis7s2mS2+STarot+Q
4fMN7PLhxsuuhNH6lmmzdrSkhN1ogu2hi8u8dgAz2LfkmjTV3SqYBoT2k0eKCqrh2JxfnyQD+SOl
WH88lzHAa8wfdz+OY+n+SoDWSVH5hGNteh/Y82h9qHj9gtGsu/zMPVenUOtIMY8FrvOuuKo4Yne/
1OdJfoCxHxjMKCT55Ai9rw35QimbVab8cCF1/4viCyUAozmo3mO5vdyrzArvdLO03r3bEUSgBtgz
g5ToBNHQF25HJryG2+KCmcKtnAi70kKBtbgtyOag6Yf/IR9oPgsnOAiIR7EfHunNSMMNS6bNViBs
sdPaoarmTZSzI3AwOrFxl16JXecAbF4JrKPfmaNakoWmlh2rwUmd2JkflAxEB2QNHMVFU1zjkd3U
+sLQFWGQYD1gTPgBWqv6rR9JVxOFnltnuBDUOmT1m4LdAsAPdCqe8J0vmQJBGj+mGGOgZUe1uqmC
4ljbxVCPLRYTm1dHVE5ew6catmT8nLjnBI+57usHmHX0e9ejYykJBEzs2y0tsMduUMciJ7eHT7Rv
+x0uLr4scZ0aqEY/xO6eNlRs+Is/YwJsMQdhMt6tSNOZF8B+8EfIEDHmkfI5z6TuKjjeq8+JsdFA
ajbYKPb/kAwUxJaOva3aIvSIyoKB+neIhsUxrwilOEl9S7SCm77X83gVgovc1bMD2QBzG0WTWxHe
TDPrAc0RX1Q0t3to7Q8eCKcFE72hutRweTH1yfTqQRVl2JmOqhFUIo7NBUnU9ztCiXdLUR7e8N5A
MxGh0lkB1gQP3uWJRqFu5Tzhw0sD4uPompJGosvNLimoq6ZzBI0HPKASGKoI2ibr2agRjjVF3Jk2
eVN9riN2as/g2XzKLT5yi2J2ypm9lc5S66vIDdwcByfZxpx8tUAUR2eAeKb3B0qbVd4Agst7m5nN
jEQw4NQuOQVgCXu5GVU64kbhZn1fPpC24x/freJGQg3EALcLkOvAKgHJZpMdVqDb1Txvj73xQrmK
bi17cyrzANlugHqiex5EqT1WfxMERcQffuo2n3mzEZlMvwo6E7Z2nbjvF+mCiZCHKJBF5StPCXIG
zkqYE96TRYW0kI8xP0KW40sTkabkHAgW9UIz3m+FynrE8onrSSBPCQUdLQZ5CLT0OwtkjRZS98Q1
n/BUcq//23LDbOColm2RFVN/hA/s6vEhuruPW+sX3cEitwmCWOGvexX2uHZSu5TTa0z20lceg2PH
VlVld/ve/lOd1OjGPJe1BTN0h/zGxlCBVFkH/VwPp8crTmRCxmJW0g33+kA9ARdTfVBHY3duPV4d
+Xg8XshkAzeiTrzRe9RfrPkvNhtI4gy2UulRZQzD+LDQyWnJeH339i4wNWxmpQZ8kixNl8LadMyv
BBBOlj4aR8424xQUQcRebpqN+q6wvP4Q8V0wlWI2D4W6ufYm8HeWkC8ypj/dh9Wnimmllz1pe6x+
rPr9m6PVBRx7yo3lAHyp9RpExw+Ia7UOzl6Dd/zgEnkp+f7QNlh0vyM3Xg7T6wFXSGZRUYSGvCaR
h/byd3ZuRU0ysMnVxLw/0rPqCg/eh1uWSE9qVgyp5MmMJYIbTmXEGuqZYp/TXTkfppSv+2sMtO5+
UtNtJReUHi2LLWxCMfxqvyExXj9D6XfhA/0eo9+aF3eik6swSW6H6u7DtVIKtr4uqhZacvlJqIBB
PLn3tfMVtUpWJai4jkUaXdAeTHcgIFGRGLc/9aYW/1aNloa5OLpq1r3iePWCDc6Gvtzh3je9UeOO
sDzuiEltIEr5WSwd67tJHWF17OH4ooOEPDav9OyK+qC908yUCoh3okC9mo7NiHhSZiERjBhYpllu
Y2AQC3e3Ks9YD77+eqjYmiJ2Ise0bAy+A+ZZEDlR3OfP2vKh7UE5QznInRTHD4fjHfgYzNmZzr2O
t0iPaEhvYkUDWpDNMKhtllW1KZQeyK/uwUnvjXaiZyWIdQv6b5/I9WX68HMTV4mO2JLqVyoS14Q9
qTW04aIEhmNFp1lp6HD3H42p97Cl+CYG7tGoNRr2s7/zFiMMXPV7JR9SHscJ4OVXKsP8SX/jMVVC
1yv2WdSA3fJHsXBfQ5rsi+JllyoUn+zG8Q03MwsUyWIf3kl1LzSMzwN1pHKTOY/aAJYIshkBqEnT
S/9Y1zrmEpr7yRixypSjC3NrUVzO2UxUGYSkhzgdt0p4BAlkFAOvKuKry6N8/gnf0AQFnYdHlxHu
ZTLb4kf9I5VBSWJfL8SiqdSq0t9wlYh6gAo/CZxm3s4Y0XQFsbkZchd+hN6gGOgacbjN4chJI3ie
tXQqwZv6LmyyyIf+AMtA26pPL12ELNlHqJwbzpeel+/p/fiuOSg65ZJ8XmjbFp/d7e241zZMUUui
QfNAv+8Jh7ZLKv9QiSoT6SuWkM+E3MYnGk/NzKhGo/h3h8/GYCFU3S3gkpnUxKVIpAQTu28laG40
Ml2x00xgfGy/kMfvIokRWgKAa9JayYnwCHLH3HH1HmHj0NsbByRKMiN8lJHW9mJQHP1Yun/RZu3R
gVeLNzYhXGOc2uqvdfpwWeiiXqWqk/4/3onO1hy4KpCFmHxWy6xMo25+67Y3RFPKRRVRmx855bdS
vjqDlhhkqcniuWIvBLVQ96D6uxSpp81CmuPx2qvsUYYXUFUDx/pPvB1y0IT/XhJpMSPhjPkAXV0b
0pjWPuU=
`protect end_protected

