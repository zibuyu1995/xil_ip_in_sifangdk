// -----------------------------------------------------------------------------
// Copyright (c) 2014-2019 All rights reserved
// -----------------------------------------------------------------------------
// Author : hao liang (Ash) a529481713@gmail.com
// File   : simple_tcpip_param.vh
// Create : 2019-04-12 23:05:57
// Editor : sublime text3, tab size (4)
// Coding : utf-8
// -----------------------------------------------------------------------------
`ifndef __SIMPLE_TCPIP_PARAM_VH
`define __SIMPLE_TCPIP_PARAM_VH 1

`define SRC_ADDR 48'h5a0102030405
`define MAX_SIZE 16'd1500
`define MIN_SIZE 16'd64

`endif