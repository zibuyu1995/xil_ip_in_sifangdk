

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CvmaYyJzAT4gGJRlCkE1yXt5Lv9gJbr2gC0wBzixkhI3TupXRLTg9s4Z9WVWp43QDkUuM3VRZjAj
RVnqESt3JA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hHyS2uxRkJ6sHR79RwG8dxYfMwySDoNzo0ZpVSoiAp/93R212I5J1LxM+7EujDw/cO/x9djlyxbz
erzC6/tIqQ2nS2hUZANmmER9YkiA1RlXlIqDOWo8pOFHNj1c4jf7Zdq7OJMDPvKF+fLgmk5Lu9Y0
15oIyfQw7L+gXpW1qEU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Cfhh7YIOGyVJiZpd5j8xa2ugbHZdDDpkNcw6vvVCCgnGCfzlen3wlGk0omzzJqyVapnfg0aPFCVf
eH/noQVGu1bQkowx0JKcNE5x1v5DKH//UNI+lq09SNF0WKlMcTAGlNSUzO8kgVv9uNbKUHDXodcD
5iGh6bHMhVPSu1QKpTfJlIMd2CMz0JfDQiVbfTaAGKvrQhaqVte7pYpnqiXM7povPwt/ntWHBH4s
XSF4J4eDVLMuQmQNy3vrqFdEUqmQFtLWgNRpG2fwo19Y2lRzT3ux5SiA0Iv55uR6x7AG21x8BZlD
JC102ufirdrREfWUzlClY8zmr+TUHpTF/SgPMw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UWceDgHVHZAg17Yudaw03bncVn75AJ6y0RYlYeqdZU3kMG9E1W6q5REaQAI7sMZSrC2g0zavsx4w
utskoq80P2avoebtdvBfjr/nBCQqUN3AvM3GSk85froboZgk4fCQ8UtEj2Qk7ob+ox/md7d9P9dw
2YULi+eG04dUc1g45wwF0ZoZdARk7Ml+fXMnm7zxmvqVieAEsVq6ETZN/P0pwvIpAakLTayKriGC
qcrb1S28bOuV+Na/FX9rxN6hM5aK7vSdFqja5GGs32r9UVRIkX6i7uqS9pWQDR0Qa31W3z6wrRrT
+2wzEwNMDKYuWVIM1FQo/Tp0NKa1Y+kyjahSGA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tLsJPLnIUk5FSxPTGLkNhAFldHrP7oFH8h39nfqyEmnC/AmGzR3fePfCEcee3I4TYySABpWhyXIf
m1jGiCuHfIpFkF2EJqjWmBev0bD33cbw1av2xtJRFa5gaQjxChO9URfjedFvCQWWwjlxejc9nD0N
O0V2XUDQxd573YmSBuByzshlxt3bujEd6Xeeb8N8NI8c2ZsfY4693LGdb3k6gtY9ZEoo4XuYVt6n
S2tNFVJTfQjyBEXbuCPqpwGf6bPdy2SKvTE/s4rSIVTO08J6bXDaEOBUGg13XVoJJqrayiJRVuQL
LhoiPzgOqS6ude1uUaMHE/SN9X/vt/6uOsOl2w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jgk19ieS+ZYiySHKvgAHMus0OAx0HPJ59p64LMaYK8CyW0wSM8LIn++sFz9tsOBdLj2gb8IKpSVr
SOX9XXXM2pQFSME7x8q0m+EPg9m1+ghIpW4bU/w4zVq4NBjYydZCI0Hpy+X3op0a3+eENVEw5SoK
4R/zOL7aV/2nZ//wkaw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L/BPRr/PHH5da1O06dKRr5ST8eskM6lzR1UPuTvZQ6RCsFEjTD1HgyqjW7/ypnIq7V5TYDC553+Y
rJnEENzDc6RSpzenrYxw7NrURpUedIWlCc/PEf5Zq9gu1ESkpND7t98rc+uiAz7zsn/pHD/K50NR
q9l/gcWkOCgArmADo1Lw9usrfZ8ECIPKY2kLxeTYbh4fsrCpPQsQUk4NxX3N1Q0h3RRUCdHSFc0O
lvGip/vd24OK8zXDMaQv4fPmgToFQMUvLrJXErEUeRlkpxkcX6g6Zu4RMWwwmkNIfZHpc5K8Q3RL
MMc5rARUSXbNbpf28H3iyAMZ0y+EgI0CrKwooA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
9Zmavc6GF6DAbBhh+BAv6W/bOKWXbZ69i4csJLutdVXWOQNj6QzDivFqFre9TSBBrcL4vV+c4IUl
JC/Zd0BOlhyvUIMlgKNzOk2v9bDxPaTm5NIIW/56+ajlc9u8JeJt/0mKKoFUKR0hbACjPMD/aCyn
izlJWUuYLZm4Wv35oyFt0iJhwd+CbVak2zD1TE1AR8zZpQ0jh9fYXHhBn7nY1mRtMASumG5HPixk
ud9VnVwK6wqkD+bnV2KBmnAqddMh5FScgKWHS9UWDxYMlncy57X5XhbZ6ANI601XLF/uVKLziEa2
t38ZqQu66C1mo6ywomBXaUfB1o37z1nl0HXZgIGAuEugi20XeDWEMxf3zgrcQv8pOpto4xhFrJOo
OzE8mKlmhtp/vdTGqMj/nRMQkaR31tHZ2RhjeLNcC+x31naDzHoIvc9Ko5V6mJsU30jtEAqSw/xO
CVZzw19qil+8Iee8g+OTrGU1YPK46ADRDPoo0kbh9Z5EoPMmo93C7U3CXeUltAYZdt/a27bLASQq
gPwRj3haeuXXRDfNWrQ/5NAwWlyjszqcjzusqETGYknk9ixEDCgECi2vqXteouhv+HVL7aVEJhpE
h9Q6bbMjdwnz7OUHlfu3Iv3cIDkJZRpW7zgVU8Kj2GaXpTNYF1b3m58vCXH0eJsbuCsQugyf07vb
H9RsVdMKQzhPy+zu6oKLTUEu743JewysE0K//pUtfAwGx+z1w/Y/LalXloxpXkBj4I4uvmxNqZKq
z9ANCgC+QsMXCc8aRyCKRi+E1Q7gvJ2cb1oN3zI7JR8JLtUbVLH8iaXA6t4hdbjG1gnjrN75/Zzx
l14+hpeoqJsKVfHF/eMhVOGPc8txZ+EmwdZ9cXXxzDR4X4ljwrJfSZggN/dEIvBs5OlvTGXfct9M
CiKGC/HdrRukY78YCPvOHE0I2nvyn1ZUZEu+DR4AkTpYs2SsNXd+gPIPk/q1imq5Bj1AVt/x1ZOJ
s4t2pyM9ogeX6No50m2A7DvGg5xFFpVE/tKi1Gpu/FdeXzd6eTc6hITHfim71cRd9qtxKmDVQJoP
dAxmh61IotnOAY9thfWcL4L4eA4F3OYi4mG3jbUFNoJD7Guk/LjxyZmMmaO0rmDWb7mYlgR399gW
rF2tGVzFe1r8CrNxwEqUfQinIR6AejIhwcFaPxk+SLw4JsVhezk2xd/6ak0CfQBmVornRTGkO6M6
8fRkRT7VxEGsCj017ATIO8d2Gol2GqZi9xAYZvw9izK+ONPuBTGbEBor9VjOiEx73IXNyWXWPjDX
0RgoRj/0RjVvZXyU7713oefrnM+m0PuXde1qiYIzkreRXPrGZvMHfCd9BYyfkSbnLbaov71s7Yzw
dUg0DGAVWy5201KaK9+n/S0G+ckkIDq+DfrZRBfmNaC8uw+CtjJhAvrQrq3u5AJv6BuXd/2p6F1/
a29XqywU/kI61WZp4x9oZBX8X+LGC/bk4fuU+yijhIX1ZtnHqexP3BsrDUF376bZ9uctLlAK38kK
ZCHMgdjQJEI7evFWAk3XjEPX3NEGm9B2ZddRatYSsu7Tuehwbols0qiOkxaYUvyFV6UkizX55N1R
lIineFY6yt9xrpWLP9KzSLIVxq8gb/OnRA2lojmF2W1+uVLSOBFQfHUYhYnXpYqDeuTF+94PPSZ3
zqIR7I5oDe5HzdK2/jOWP2xQjAXUy+fxLAXA5MwXYAhgtAJvQ+Eihldie/Hd2AjJkz8jErG23x2G
55HOEKsul8BtyrYBT4ecON4WfJTQAFZJsorqSdtdH9hY/FWtNHSe4Sf0nilgpaSbIfchWFF3YIhW
o/jlo3VuZpzMKSkXpp+NMXopOWZ8tqKnjGaUrXFgadXkIo96iXcDUHvvttu9JkljHAaJPz56lLXf
vUCJXy5YgqGqoLqdN6zUGw8lorLmyZmMfcNPp0gHWKWWOrRAnL/iwJejLq1amNiA9hTYuL+eyOok
nE2OAftUVHEaL+l+hq4Dvhu2bl9Nl+HYNk2dpK32GUDx/8v2nTHvGUpt09OrosTnQs6lB9qRfXiA
4IKoXSn//t85829/ddrh6zq73vA1w0onpOEeYgoI8L2db/IIYiLfpzaNVX79GK901a0gEPgKWb+u
cTG/TpOJmQRXsFitPfEKILe1OP2c+vRXP9Fka9lno4JYrlmQA4fIz6KtHa9s5yBdGHZNb0pHIyro
8PWCReDEnqOast8tP5IaMwzi/WVrmN3NR1DExAL/5BH/rjHBY81lGy/395IL95sxtBdyT92E/mW/
0vUpzPUL5RhtOcmbHc9xYFD8xjr4ztA+BNK5Yr+dA1HwJkK/gESI8xH7ESaDWDcDpxYbKFrSEYp7
5RHORVaUljlDKMTBc9XrwySwEYXJEypFwju2ZZuxfe0zRJ3zvD20Df1QeI9fKci+qsP/GHy2sHyi
MBm8aqr5Boi9LGfR6J5xPYQxUbuiXVyJLI67KMfdyoitfrhnTrbBM6klK4xxJfO2D4ZESacGOLNh
QKebbFaOPdk9Bvm7zmDFBKjafxhWIGqmhtwOlq8y2EP6aJ9Emr9Mk+15KcYWH/UNBiIrT4yzqzQr
mhO26BohcxmpMrLXLv45utqEI3il3GCIASuRo1YNU9kRuFeYhXZF6I4MCHnyPfI/kP0uzf5ILmeL
+m8UI2oPdSeVCj9K222QVSBmMsRxZbJ96SjDoc3WW+oI4/5C9d85cQ0vU/dnpZ26mLxv+tUHSgIX
qS0vE666awUNT7fGapI2HHm927m/BxaRLA6aklCpTCGS+ELBXoh62wA2OJ0f9hfim2sVYyteFl95
sPqMq2KwsuNx8ay6XJCHuPGrIUXyVGzSBlXTXguGDozJtCTimCSFfYft9hESCQXDVbIgZvzKTDEd
jiw8U3Bl/wregYH8YhQJa8D1kTrQhwGF2o3HowAoUKM6tgjjIHzbj6dmeZJA33uR1b4JDjH+MdU7
l02JwwJbZuoEmKT+FXkSw/DkecKYXFllv/sg0z2/a3g35I9nXGH0HQmdNoLAsE6FPzLOB3GFD9MQ
cqaC5MfxSsU8O01LFoKzLoBOXw+4bItooWHCNalmdHAooz27ABNXqJbpLxK/UJb/KrB8tHa8pXnr
+fDpOc5apPm1qhBzZr9LYjkwbzWl5WDcXyd7ocrTaZXZqEdf87K4V0ctR3GYOznnOZB/TmLk8Q5R
k0mQH2vT6oUJXFaJo8qnWj5UYR9VJ8n7US4xmQMtE87kAOPXjEBtwtwZsBoWk0LWkFtQbu04Vkaz
J2yIqScA0iwEezxkhHKBxSyObJdQtdb5Ncom8IHFgrMiBWLJ2CcSmPDgL4W+xanORvx1Uq/pAMpc
k6Gb1Y1Wd5vrQlYBFLKdrrBOARiA0g5YP3OHIL5C0KCTdtiCoCceMzUCQqtrMHvl5lXLzcf9934d
vUXwY9Of20vJIc1lPJ7ouQBPRj0KeNYwh0AC7SOFX2ilvEmf+GJfVkATclHTQ08DvCLRUCa8z5wK
XzDuuW+MmKiRdri70TQUsftBqge5fWIHaveX8s3h9be0vKG9XRIzpAzFXP1oJ2SS7aJ6uGDD+eUF
6uCvkV2MjhLzZ3iyHWJ6gG45RmSx4tuF4pC7ePpjCd2tQhhm/VUeuHt5Shq+HeTpmFAULZAvtI5L
n1V1wjFNvaqbfelgQjxgu69v4lN8+r0nq8E4yhbdNNkwFPoJwLG7u8bQ5cnUQ8X1m5NH3OyEZ+WG
f/gUM03gt1U5qVNuRyrODYClcDaGMA5sCvW0UxqVop+2iig4jTsUHpDW8GX7lusM4Ttzb8Qga3sX
JLHJkDei9IFqbfwewGJg+l+YgeqLv5IwaFMpzOHI7MSggnUd/Wd12CfE1IsmrZ/vAngskqAQrcuC
7l8ON7Otm+sZByKZuGWZdoE9V6SjigJ/N3pgicX2D+NRXEA211I/1DsovhfmUGPIxXfY2u6NZtf6
TLhhfJpCzOT3UOTNOeH+47TIo1BkmrmOoQ45fwBpIEbJGw/hIKKRK4QNNuXNftox+xI+bf8b3M8q
WYFL2o1N96gZGDrhvgPJi34WMuap1is+eGWTezW4KxUJqAI85loA9xDkegCSJ1/yJ8ZT8teffTTT
UwKLFENXynlH5thvz9c0glXv5M/L3JbZBTHs+AVr2MWjCR3Qbv80to3Dwuy5zz0wpdm/o8/fTI6h
/T2KhQBnTFD6z7iEUp8mbtOmMt99jttb8soqazniSzOiImf2t9RmVdwndcoYeKZ45HX9+pNRguW7
ygEbSmacIbqzHVrFV+xKSuDfhf0aZxewklwM7HIOtg5XMg4IUu7fJ/Uktj1U+LWNC+mXMq+GBE7X
OdSsda9eJJxcJrpR6wLKTvWpFMPCgKLLULvshJXCgPOEcgKAslCCCdNXWAUPLqu46D49yjH9Bp0L
FjkvrRIhQOcCB6zgE6v0sZl1zhy5fe8hadKNFBGSBadlBB3j26YW+rL5IFOLKXiv7oYULHGsXsGd
BXvYlTN+oHShj/laI24vsrY+fJRZckxrbhETM/L6gdoNjbZPHuhMQvK4KeURkGCcAVdlEvFvYA96
KVcFWGIMEdsrrO+QBvG2xJQ4yKQRr0C+IZ1uI6t6QfMw1QIjBR0ZY5HSZXY4OhGAh1tet2+FtV/v
Cc+rMyD6g40RuTzCOrgElWWng1QBsMF1oKa+u8tiurha9CVE/K+/pHAKoQ7+RBvftwW8m8amJiRP
5Ulm1rOr7N/PW5qidIaWd3HBLGA5jadVQfleKYF/k9veFwxpZ5tspkWgEze8wPbw9yoggQupbZQ/
yA2l3WDQPo3CzI5SlwPPxSSRvulDXTPaL4Gqaeo19v2j8dBhZG9a0O9AwJJXi/I9skpHi3iidf16
M+Rfucy7dsexXc4XvCMIHW9qlw/eUC0fiw7oNtvN3kNlU1+kSvrWkdP6LAyVrQ5UTPug3Yxg9F9X
hUUiTy028o24EqSJSc1XJzJ1jpgSkRstmCA00iLjE1Rf49Xy1PvBdArm559S7c0qfYsq7DoVnciz
onYDyYCk4adJudyX2roKGaDSDTDlhc6QdRA4qGhrG+jlMLZfTOuLziioYPoPDAmjGSSBGLRN7NLG
dHjPmetBVSUzcDw7h3WxHlD7hvcMonh8pCCf55pRq5Le804uTSflbmVW+9YdSiuNTj94u79aEK8c
3V5UHlUYyhhq4unOT1IcWMmEMh5RsZWm5vhHp/pp0wtY9/qJE0TsdNbWtLp0L7B9LcI91jXh/X6e
jCFIAyZ3re8dS2nEYxBzv07XYdeOX2LHyhzcmSH04AV6T64uZPkov4crzyJzll+vwwPhEEt74Whp
P+PGmk4fFXlxI/NRvOJgfGZRlr273PAo2LhawkZskJF9l6jPqMpmP921bMbKu+vL8jvfdHpYRXJu
QwDeMRHyKeYx0y6HlN0xrxPNZKKPKcp5n8g8VkrI3ML7O09cTC9t8TRf5TZy1rzhzBipZ4EVVfU2
9EopSND3ZLl43LyhpPYY5aS2UqBS5orSrAhVSoLPQcxabzOw0DlOk/mFFZzqPySx012/lzj/CTRP
dHTKQul7+8Iu3HxF+4FqQdJFGv7vMdetCcrwYPCBQLfmMDk8EtUS3HfA9dBciM/QR2+bc4dHEgpw
quIQMvLJWChDeHYIlQM2G3kggKshK+48eJw8K8vyiY/VEMgBdFfN80kFeWGLcx0bul+TUB4cnp7E
W8nV9wo230ViHmpGFP5+kTfS11bUIahRxXt5FxOfv0aKbKTWd9YmwY1n+3QIEalDmQNm7rtRVOPD
n7o5MBxGEwjK+mhcT6gfxF+dSFiQUy6E3B2fIR9lc7Uufyve/qnkN5rdNM6ki6GcDw4ukH3wdio/
/a+E1HdwJGQIhw6lQarISO2SoPBDxePsXDWmr5m5RLy7ulihpAj5eZR+UDVHz3klcIFQmxIvkTep
ZAfl5lrRb4eif8czI5OT/FpszFAG0JWuVFcDXRTiK1hrcAegE6s6b4JveN5aruU2tqGwQA29+ddc
SA9ZVsx/adx6k0d4RFwz2vPdkBuzWmVtTLwGpOy/T5RG6JXvkIJ5JeSrOT/5wXF29ZE2HBQX8KGw
bMECs8cO39cc1DZf67nvfn1Lw2TyVp/nzyYh2IpZZYmbd8PZyavGKKytW628pQM2wT5VECn6VZ38
hMPzEEbsZzp9wbwj4V8HlAG2CwUF3jwOOq2ZH3RRmnTzqIt9uD67/yLxMKX25JyHtb+Iq+14COSA
VBBXJ+6TLARhTraf3yniMCvBADo1AYNicEYzRFc/NcNeYvru26cbjcTZwcthBXSlbcdxPHwb/+pL
Wbn8X7Sx6MyrVV6Nr/7WVIW249CeQsqrDreRZbhXmpoW9T2JXPQHvm+2yAznJCzHCcMvES9WiksE
SLfZP618xI6JBb+QrQ61c54Cs27TlpeclQd8wYa41A+j3lBVjgQvy34dsGNDYUx0z5DpdJo36tEg
rVNnlT38y54J3VzCPoJ8qRvi28BBeorCVRFDtni3YxwZHVODx2rnFJy4GVOu9u3Nh8Vk7aCu4tTy
4bdN93AZ7xG9+3FkpNmH1X1wzpzqCGp1aqSNIL/3IaCyelQ2QCcr0FHB5sRgzr8X1DyHiCBQoNGT
4neX0N+3+mcG4yHpy0XGiF4uw3bRfLwR4wlUwSRPGCi5lrxqpukQVDh1vZ+3lwaYutFK+fecsuUG
vEv+kmcRH472AcNhO8FEn6LYGJw+AFM7p8EErpknuOVLhcByfLJb6DcE7Xp/pPk8a8ZRoKASJZ9v
i2Bfw3zi1DCBACFdgrL54t8kWggRksv4pN+m38eMynwMfHEycyPmkUpUVM4/SnPVdFJy2mHFI+at
RlOkXR1AhB9l0AMnVF5vUX7ocU4thPPtSJ8GKyH/LkOXFWB4t9NzY2vWtVwWWWxo23Ui6E74fb1B
K+3Y9s9qswiKCfeXA4sFwwIwlnv2v0dYAWKfGQ6oKOV6nppDzT3Q5mQk+0at8zYJmh9LmS61J/rA
HeLQWNfaddsJOxx0nvz3twITbrZT2mmwEBYY0KOjDSAHuoLyQpE6Zp+Ktag42IGHWTRSxGti16BG
iKXGXGKmRnji+V1TbWXYnxud9wduS/VwFB0pQSaAR7avFhPgSztmpZ2xQyTw5nFsKenjxqKBCa5V
8QtY9qcIVlQu7gqSa7UZ0LqBNUwR+Y9iPZs7lln1yKis0e2PYfpPTgyh+4xEApTZqlUkpDOscFPN
K7wTEqhFUt2hSepvVcCMhnbiVLG9FWL/Cr81UHWj6kF6SBjD2xQWdF700DMH/xLQ1QV6nSY328JZ
oxRdyY86jDWxFUQACNz+t8GjJQTUQAb91AWn0BlO+tHa9HIT935saLVPF6ljSVHbtsBqiggoLBM4
bDSdElK4rvxckET9F6Xx5+NQp+0rM7FRon1P1eud7i3AkktP6a0WRK8MzrkA/44f8zdzrX+LWUj2
r7ZFZv24mqYFtMxGpBU7TClkFA+96bd/QfRbo9DgT+Ji+vBQG+s0W8Bld2scT6l6W/bOqnzMdSru
ayCqSb0w5+zpqW8htbZEfqPcstRrDRghuWjxz4P03mekBroAUq31e8SIVWNam7E7U+2pprcxPO+L
eB/4VEL5SX6en/jam1xoy6XBa7Ml0vjnNx5z1az8KyA94Z6sXRnbGel5dvfC0QD7xuW0aMLGLsPI
TGa8MmvsX1OqbVfn5hZ7PQ+l1JFScunFEbjm6CsjHUqIVsqJym0pfW7Qjb6wEkJ21DsL8zVwCIJN
cZGFr6rUnjo2OQ/mmOVBRtUITceBRSdtvXdKQ9tV1bhV6CLBq0ZXZg2yiQI7+1u4tRLoXt7gd3HS
f9avl6/N1GllHJwyrDiEmOxNaO5CpwiM783yHX6dJp1Xy/XCH6Hxu+SlQ2b0senWZYXB/9uW+buT
l8xZINEPIWYI5YjZ8dkmVHeOtVAzX0FT/rNZ34f5vkp3zoQVgE1rP/AVcJv1EACA9lfw/OrGGWWM
qBlwYzuI19UNpDtJOLZAcjhWD3k6EWn1galGqUi3IcSKR4wf+4ALcQSW7dz0cIW9lw4c11qDpOIT
KSkpnzm0pCktphZ/0ZE54/C5vxqYK5Q6hnWB0Rz0AtAv4d17ZMGu53OG34MRnYOvUB8cc28Ohi5K
ytvdd5otv3/pnX0IKBlzzhTIlErPGvUCQde2gcR9X42eGD62e44t//1lXkRkpmUP6Gzuz09LPJEV
aBo1cqETfGd84wCkFMj0XccWPTjU7KgJ7MZs+BrYNOqrO146TC3UJyYGbw+sWM9E9W3OHmfd650a
FBx8OTHt1DNkSE5hbnAS1lQcU3uk2ePjgSRPV+2gaJDJHHFIlbtaKAOJugSYsKFCkSNYn6ImaJqz
KLYokurjkY4PnbQqkwVIOv1UEtsNwxyoTg4yYZzpgJe5TQWawkP4X9ay+Sq+BfUsGVNn4j//sAiJ
IVumzj+W/iedZQRF6cNJZIDvPiwStfTOfjLyKw8gWWqNCcgU+POPvhYWgeSNJTLNo/butcCMAWLu
CMtr1AcjYKRB0Hmo/5CsnKoUv7rzjZjUAUsYzF/1rDfxNqvcn4wtW8ANvNZVREblHAjmyeW+CxQd
2NDciSiuUKp/U7/Dbyf4fANFKv2Jy4rpXLpb9JIrHIng2hnhlk+UnwrLbgYYXvlgaPTSP1AknXtz
tEp5kXnKLRIciKPEZOu5mLqbUm0YGDRdFXv5B9xIkGMEdgIKo0c7Jv/vbd2CPyHpmmjm9AtxSh+w
WyYcaOUHib8cqnNlTw3CB+PPcSJvOK1lChSQcwJnlv9ZtLONipCgL/AzDxVTFWqFWtYxB+n4tvKf
NNbbpBAoyv8cL+yyi5GCYtt5RMmFD7zm5UYV4e8dB0XKbuC2btoQNHGP86iGVQvmAo8fEnJl+xom
ZxP2+PxtC7JqZ8oFPiPLH8LHlx4IP/LtE/oZ69FOjJBYUg/l4+Kon13GWBgalOZn+eRKs9GwqZwN
WIIeGOSV38OkEUSxLhlqtwzAr4OOKmcslZuKd+Q2ivtD+n/dYb93Ti9t+tLYmDPSgQwKOT3cwTDB
eOasoNWLv5mmta8XcpryBxaLxW+jdDltzwdYdkRprnZdzK24DdbvAX0ECGryAmoGdmDsMg5k4YaQ
dGgJQsQp0C35XUSb+ioR1dJRIrBKoKujM+rnRPf/tlQEXw5G1pCg7cdsCoduu7vyeCsm3hopIZWZ
72l3urAyjBigyN8Ar1OUToX5P6ZqaJ/hVBWVyKF0NvjZIHZWEChniNcPDTQt+/+MVve4lSMEaA77
g/EmQJ5jFsj/mndWUV8dszFLbLH9olPt+2eZgQbt3T4lA3umoxHuro53nzkLiV2XrXxaC52PMmWn
V6GV2PMO22fGQPoDdZSHugXt+CmNKppyDFEhRoldc/IucLdz3pxgmguzmu2/I0yC3v+2X1TqIp6Y
GKKo3s0GbrZ0ZJSdIt5U0BVS4t7yqAa72VUZzvQ8HTI7MO6Oa022694w7e2gJaNeGEjbjGtW6nbr
js9rWTztz1aHMymK0HJsEFbF2BL+IcLMwtvxub8p2wcoKknmm+yeNM4BpjLuzWEhjOPVo+aIJEpZ
vkJZaoMt8rsNrjSxs3AH2/tw03rUBDWi3C0TT4K02yCxdGV8SxqdRl0Zyip128BkkdmxC7Jtv90M
v8r+z62omW73gxqFKprfCmamXnycKl01u5aIwpVYx/TZqv1ibtBEbyvLW5zRcDJ60euU9z7K/dzV
k9aPr51lbXTBqkMpdKrlNle3kaCQk39/cdTpPr6Z36OhEGAlyEhPaIiHmNg/UOrURvxOxdvlFTCN
+3MrBPDJDzFowNB9vz62iDfVcD0cX27DJ+eqBaogTAe6gkLI4T3RydZa3mfVjmTPMEgye5PLgfQv
QVKlWJuyGqrdzjypAQxYKtpvLDgtusLcNxOZ+9etqM6+4ASIoRHWpcjKvUl5T00DEhqNYIWHxyRe
TSGmOtWBTk/nymNp8TzXWPXCOmlm1jlfwMy68G9nlaavHMTW9mClNfpo+/DnBBzllCfrnK1l/Qfl
Y7zYdHxpPFdXKmf1vd1vgY7eEkKhGDCbI7Su+2Qpifj66rrCH2LE3AAJpL9eBwCk3xWlonx4rQLa
qXr+vsmsoIvQVqxvLtvJR+dDUK0wSUTkv6Kl/i/ln72QDkkodgPL2wdKyVDWd5Bq1R37DhfOECdN
5/pmalunwSDqJ+gLpI0n89n691cd7IgRUAUhvPIJNOzbggsRbMgwWjemvr+IdfedPmfqJLBql8HC
R2XfGwANPKtLWhw1m75vxLvX8VKoJBW2gate2BvlLj7Al+1Pk434zMhgGX2kLbhZgAnJm6gxg74u
PnRiqvo+Rb/+ERw0IB54UBB3Q0g0UOlaG9dUE88cahcL82p1LetVu+GiyGZPfV+ZBZ0y6cYJ1Plo
YFVN8LAaIZ0wUn3nW7FMwN2g+bsmMejUCaj1U7kTs2mPwaAsnMq3nyxUNxsxGr9vQwJ/p35fdKUs
Qbpb7Lk+Vn9T3B9Gum5mKilMmmUIMa4bYEU5GvtjxfdN8To/VcEtuLg2iCFG2ipogEom0Iwi+1rB
gp0bp8CmFLWhaM/lO3thlWQidW5iYW2n8C9Fw5WgYCiH6BwZqjuUYzo7QwycNV1CGQWt6gWYm70X
vA8eVXrYLktDBq6THyyh6Un7trLwAGIZeUqDpCZcckIQoWMNNhSX/bs7aJS3oBn1IZIdLglL7BWw
rUnPL7EP/K4O3WG9bJFabv6TiP3xMvVR/hJ0zOLvE5HdjJtGTe7arorpV5NnPhsQEvOxtoHPkO4B
IeZcx949xjz1gCaXOzYJSmF8N/8wOjzRDI0JR2gi25tWIuwArUsCVY4aqSOkIYItZwxBbSyAZeFV
VluZrWVSkCJwBMyiFGiFeidYW4bXVGnJNKar219rzEWD6NDn5M6HSriEbtcOK/k3FPlwFksN4R0V
2yyVkYcqgzbZ3KWCNb1Z2hosrVv+EYYhQleWGP6GnawU0f/NBDKFq3O9WIe4ytAOVNTNi8n5v5Iw
iAcUzNd+WhSepA0I9ImOaPLhTjz8WJmvGEDNNTelDgxld2AlxuCXbWVzVPw/9SJPThmBdUt++YuM
MJIn2iinVRf//G/VfU1dRpx83KUKHZjdUXXm1H71YpNKjCdS5MqXMAjlhyxp9MMOyoWFZhct/5Zf
+e1X71CE23stwRuTtIIFh0xKs2HxaUm78bnj8XKu6aGYre8cEGLUYid6z43Sr/jpvMad7O1d43rR
T0Y4jJHrmGEOsRRcxqZSXbcz5axiXKUVcqqpLSkAYkrzSb8gXvTPJbTESbYzZBT6VPkSawz8p2lr
KDIrd62M1PIsuvK4qEJqwumTKTnVTzjdRkNIPL+dkNXRtzsSZ0L9/teRQE5o+2sGDsl8K0VLzxy8
MfEniVKW3yo3Bg+FI+xbAToJhVcJaFj0l9KuWNAT4OsXu+MmE9C5g3TMUGSlzVZCphPuaQU8mPVF
Xsu4cXNAiZgVVvid9eDDxK337cXLym+8yRW+nZeAlZ2oQ6/HrYH3bb/TZyC4/cu13ulHfRE8ygpX
vzGHGpeonSt8x+lMVY13CfhN5evwyudcATpMMg2bA4PoQDWGbZ1bIiR2x/k18eS+k9T/UCKDp6fO
cu9XQCnTkrlwGfTJpavsGefq5rzrtqKlpYC4M0g3YKXHV6Cz+Y/0DucSCsua4jr2fXbtU2jO314x
4jikujnNYj/jgUfsq73XBy+XZ+K41x38KIC4v0e52SHJJ+mUlOnUtDySw13JxU7jIHxE4/DKlz3G
k6cM2q7LuGcxkrcKCzCArgWxgRzGvC6gqUsFJtuMUKar3DJuaqOFrD0bjRAJZLbrxHYEAGgizyNq
utof0XWKw92FlVVTM9LIhWeH/nSDHEobFMtoh1jIzIxxF/EKAbckvfhykPyJ1sfPzQq43UIE6HYI
lH2W+IMpcGeLa4U+Lf/ZdcH4XUH1llUGfZjoFpe+NduWYvogTAZ9OMsT3LKuKr7y905ef7aFNCZJ
4x3LP4RHyU6/2czJxC146Ml4y+zR1opsQQ6ERtQneHFTz4NmI/MAx+1XdOv6VqdnbQY4TO6lZT6Z
CGOYPZ0SZn8dvfwslUHG+mzwuiu2jp39Z6Yo6ekBOEMRK53N6VJ6vhDLmLfDyOhO7/YpYKZ6JgAB
Oa6fRB3TctJ3FLTD3T9LG/ZkiCHovEav2ags0oN2jzCeMBMRvupTjzm6u1G4oN2AnhGY7a2yV/xX
kpNW+gjPEN6s0tjCPQMEqV8UTA1weUWs71ptYXyZtzZrzxM05bggY6lr1S/lqKFpjrB3MtLvGccv
y+OZASnuuBVdlfgHltDkyDVkGAqzyfp5acsLw98Pftet8b0VKkag5AOz4K8v8ZiCyjAWZa3YYFdp
45KAmGkS6B0i7RwLkDs/tp88ehB2NgGKW/ks+SyvJ3iiwEmZI2oMeqfHJuzElaXr6xjmxYNSmVA/
EDC+Qj0BW7NbkrlX5pbDhXmPJ/Mo5JFkgKFFQwF41kdiPxyVpiN6H3nnzxzMqdSvIi1dxpeUq4w8
IWPGeKCHmk6t0xR4akKMgVz9s5KvMqWfM24WnI+D+yMJrproNo/hAr5sKehOVHQchm+ZVSvI7MjM
Os9M5ruJZltwmSpWihfd2zkO+PtuUCBZfF9+lwaSvCwUgftFjkoADKSBRi7FxNVwp3ce2ah5LopB
sAaFxuDE//KleF20wgy/pdL/7aMbYfgQiSW2NZSv2bEZd7LpfpM+Sv0ZtuTNEVRsAdBl04HrqTKL
cyMMMjOXlzUpV26lol6WaKXAuqq9VjQzODX/YLziy5JyLA1mVW0/EfJAwqpFgZecUNvrtO9Acx5i
LKiCpD55n2OxZo4YmNSQHEQMfHjPY/cqVk/KUB3cVbii+ajSOstMWkDGMi0mzAVF0uzojcTadVIq
srW8qtoaBTTacKg6Ttb4RIP8OCgNoOVYVZWGpA7nQwTAnCmBooZIGnVqkrB4sEmjJmSP5s8ojEJi
5gUfnhZMzt4mJt0W2llcFuMJx3vzK+jN1F4HcLncKM1HXDLXx/7qqmtEB71zGXMY1rs5kiKy/RzQ
IfLjKjv5RK5F5Y52U+dbCPvO5ERFQQAFjvEGsrQ1l/LALJ9MaHGCfTaTjTmq72oNIhCB1cCQmbZL
k9NdiiqwNilClDpSXMmGe82OjBTAMSlAV4LgnY/My48SITxxqUKdBZ/H1E5E3y1k0c0cZ92MQXQq
Xcqo/XuEvpnMRecpfijpNRBioTKLywb0GDRPYrWgX4Gk0Wbl6l8PNCIZKj6Pqo3RNQ8fGHbWAkQq
V6gNvLcK73EUytOiTgceVy86Vky6hdALhCbobDY6cC1lCzLPgHtHO8WH8PIGtQm3xN7RjbjAQhw4
Dzp75PQre94xCfRlmpSEsX6INIXRw9WJ4x1BCZFSl7wYIKRzICSmBnqzHQH7Zwq+vozJvtZnTc4s
O1+XFJIjCoVO7MRzvThg9MhkkPEFJE0TqsfHorlBKGhMNdCPn7b/3PFuvAgiTIsA8hPXPFSZhzMj
zHlOwPxnYhsWDz+0K4Tutu+r3tn9Wdrczo0gmfKhEsepGETIKHKX8cxUSJ5Gc4LgyFPFd0y1HV3G
/bYlT1lvgZs4SeZLvjQqENh2mrgrP4u2woKfDI3IznI25f2uiYtkUB92mA1VHr15eB5epmJx/Vv1
JKhQGzmVGINZpINpU0f38lbI0QZxK2T8I7y3hI4aGEaLY6M1VypYBw7+1Fwidqu/HcFVYVWp0aKM
nKj/JupGeMG+PWd398hoMo/gEXCRQrUt/sWNF8ujcjXQ1/yUoGDjsE3lvSebL4n0N2Y8bJQWtDG/
X9wNKTSkmxpTzbNr8OqKv/nqfr3WNPjY3mL2Wh5flVxewo6bU+tZ8jgDq4HyBSD6cQQhO14rSMDd
krsnnWYwbfDiGQOMpjawXObnWKFa5A1NXkbDfP03NAC4J58SV042Bn7XcCxKS+TKSAFz361Nywso
YZsFZXSc23cU6LyJCJf3JK/6SghXbzpVPjFcRV8W4vQFXHi0o5YCJ4oJE3cIRcgNBTEOf52PXheX
dptEm32Juio74WLtKf8gIx7KFazJQ6QeHXAejXJMHrTBR8LJ3cpVRFq5bcnP4Ga7RhKpacyujXNq
oZjSysZdmPdT1lnHRAEQxk5hZNOEazR4D/j8zUaYObssdtV+OOvnOAlkumf2HAH4z8T9fsPahxLi
4AMSiREXCKrMTfOjdmBilpfn9o5jm4uL+XMjHODhONEhPtPsSfk18Une3S5+1n+V0cFCga9gXh02
k7kdPey0XOWMjQyegb4nSAzBGTLhe43v+eV39PfCwkdH3dcMPgriK6LketgGDMo+Vy2s06JzFvqH
KTa9Osx8LiyNCPJsyIBX5htGZWARD9Omva1f8vXMZQENC75ISFqbkjVkTqeoM3qOKHRO/8RMZrXA
31k0erqaxKYjip0R9B0jDjrYwlPJXSp0kCRLqpkFWqIHFrUb3VVLN3aa6uKEPb0Sp7GpHHHXLQ/d
48qEPbTlDPYdAlntRzyPAqfHO+od1jbaCJA5ox4pBNwxBhwQoLDB+85JLrWLjvbkbW+e+dpTplPB
aHY3Y67BsQZyo8Hy5rivfeg0jdfzzk6xsxghfP1OWhkoqmpqTg6uJX52sN4y4HwUE1eOCHNOq2Mb
b5GXC/mzw1/0ISTFzQ+sAw+Z21cVDPBaZ0U3fJ+/or1fzcGJcsnPUGzSLbGPBn9aUgIgrA3xJY+X
fizcBbf09sC0bEcGlH8j2vT6xTBZr6vMiJDkeYEUsBXvxi4QgP8S4Iz/nP1WCqgrUSYXptTojiIn
EJ8FmBQmoVd5sdwJS6cmSQd67faFZ3SMFeayhNziwf6JibzPD4bQ9dHKaeUKKFIvPGlVqBEfsMG5
ExQgjEHdD+RhaGYuLnMjd+09VJfQfnONJo8vcnXvJemRcYmq0Sh0mMGrj0l0qaQ1bg2W6Z8T+2v2
hdZwgGCt5DWBom8KQ4RE9wFcoVbhqzt7N33NFPCGGzfEs6nnp5x97A91Vn6pUPsyn0boN56l8gxi
B3Nv5bPKSdswsucnc02/px/vUY+od6chlOgY0fuVn8xAnvPKotKy4cXhFT+1eZrofH933Yq84ToR
MZ7SJmIpJON0o7SYg8bx1zjt1VyphrxyYbW+Wr417a6u3z6VtdCopOyjsBvkTRvFRW0FWZ2j7Hr4
wd9GKYNTBw4Ax+xgZW9eDy64MWyR4kMh858hwnwsz4H65Dc02FvjZ+xxscrveCPE4u8cR2xvbUHQ
VSQZfuc77ilIfCzh9Tz+1YHeq6M4DTWUiXVs44jr6q+P5Bg5ZkYfR0sCthEdn0Ni0b6o0Z6iOYK5
+CRranewa0cc/wABGYzDENH/vDzQb0/uA/KoKW90PpiKX064C2YeBufVymOPddHXsyjV+7YeWtlC
BaS4UBekyhoLWCNhTJCDTSZmzWXzEOYj5xPlxNRt44Nvz65KN+Riw4wQEv05xPPLLrfgxsgj21kR
XbHTmX4BnsuU2bJzU1Vq4PU5tWEZj4dx9lYDsHjVflhtBO6NVAMsvip+YjHkSLf5VoAvpRPQiXOJ
1RFdHjrJHDc9mStDs2jj0ZQUurKSmRkDF9Y1Ou+0mQXRfE6dLA3rBLTn13YWtehLChstIbkq7FFN
VNCslpfl/GikpaqCmRx5fAgLlb01HwArqo5XJ8JCZs76//rLPcPhlxgPJQNfXj09dqfrkb4iLbHF
EmPCZgKYOH1RbR8yXY82bnnF0Qvp3cNmbOJhddm6nfH55ryWazDelVjKTwis58vVGZKE9+Mj+8kD
Fm1bQu1TJ85LlG/li7m1jfQMrG4+ilBlrwyYF3BvaTZO4GoE07EwD9ucZEp1z7c7HIb4ebTpC8Qq
3bEK5pFPKywUr3zCyOryRThmcEKdfjgQNeCbUKM00d/nLqryv2MH4+aVOHDdGnM9p9if5KeeW0gQ
r1xjevDAZgU00q4F0emeVGQNJLj0Fh6iXWkD7LvP/nZ2AHRouMflJEVd+PJqOh2SDO0CPM7Yvwnq
L6rEPBIkTpDGIATz2B0P69VYuTuXK3Xabpdb0oSL9MfZGJikHO6jy7pi+J6da+k9iFyufckwu98L
XQmIKcRjnah5PR0p1WjlMv4gu0BrVT3x7AXeyrfv8M0LRfrWINwIAEfGEXKOgLBRR5+Ipjdoz9tH
AxMiPKCMAXFdTiIPVxQTY5fiO6KAJMUBDfphpsiq+wQxdF8cuNBlsOFJMWu3bE5in9eONyHaz9OB
DH5s6BQwob2OGhJ15qBeHMHw/LYV7QbKZfHpWBpSxSzGntREleePXwQHk9RKYelmt24R2nLEyjKJ
jqTi+pYnpH7Eb3+GS+mRQTLaoKoZ31Uk50O5PMAH+oss/My7j827Y6G2Vr4zAfODxk79X2vEEx2i
AxOBIZFzVKCCBejmDkAi3Uc3ZFfhE3vUtUsA2kssj1TYLEDyEpa++8x9FGLwkrJ+uEx167Ucjioe
+AUl21ezvV69Gfk/CDHT5dJL5t0UWz+uxJlHWnoLZ4DpmYgs0YbxBkOLcpNwE21j8JpHDRLX5nGm
pPkz5ixAWTamkbAANaPaNDxvpLcU89LxYmG6E9WErUmeZOZu5PnCQh/DFnn73UU+I2HJba/DfsZZ
3+6fFNNhEJLsUHIe0RyPez5QbHR/kvPBPd+QPYPVRPYwkQLkyfm8CqpnjdJXpjzGbMyvqqEvZCCr
Zr4iVKYaGl36FLnhFr2AKV0cCfsshLGcDAvZ9w3sl+Jd7Dp0lNfolRNjsx5lxMlqNI6518z2Tyvn
nDZ94KKNA3qbdCCFzN4hKV+ZPQBYpRg+ylBvtOMxQTpJNGOXN+eNgptW2jxUI3Nu7dCwJEOmYAHe
JPJBUVoSB4WTYAr8fCeA2mQLHud4UNIM//emf5/i1wEYJd7DyIaPUwV4hl5ihTHUI8H4xNdRidF6
ki+sU/H0x+6sNRJkVm8NcvgFlQRvzoGjU2sUECykxUYtWWbXuy/VrKN2kju45umGHrjxXLcyBHLN
sqXwzG4VwJOoyLh8FbBCLYKGrG8JI6bYOGe7rgX382mhHnPDMB+qtk6XXyz5ZjU2mLDM1EFlC0Nm
/Z0TG3zGOOeddW2oBFRzW+cmIT9gTwL4jCd8awDDyyQvgWDB8THRnJfr5R0uM30SdNMg2Cw2wpxy
7UxsMvafytxH8OzU7Q8+nguThfFh6BCczJXzQMBReGkXyn4zSQlORUdiuVLTXr5pc1j06aB/WmCj
cKbiWJR8+cOvmBayasKZJm0c/3+7zQtbuQ3FyDi88kojAW3DvlUQf763UCHIHzNTa8+ge8/kwa6a
uWHr3JD3pVlpsfbivOoGqdeiMuXUpC5cBaNJPByghLA6kGWGOm3unVBPdkXYjPtHcoQHlf0vye/9
0sXFFUce2QKs6jBwxnn5GdoJy36cYr0Z4Qsm7vaA7de4u6ATvuD4XRXN4frsCPzcK0IXjilR5Z4M
AmKrhV06ATQ8aTrAQ4m15wQoSFsfSObKlHWkSj2EBL7koDpPL8Tfgep0CYZnSQmB8zRjpZpA1I02
7KDtISDrPZZdsNCSsFvaLVdG8tw613nXgrtxYyiPEA5d5lyYM6WYKX+F7oz2AgjFPPN3IPFxpM87
fgx4X4dW/fYxo02OlhyCcbwYZEeo3zchqFZeGXoBG15RIvnNpA2HHbbU2sKymmHVHLJEixnLhY13
UPKKO85avwKBcgg/JiZ43/NeUDrxLXGUWCwtrqMs44WMlGkNn5tbv4GeTYfqlnmB3RBpuxdSv9w+
NKoAxLx1E2FviS49DmBLOH7aYh4mmSvOOpUAe0SzA4NJvcHhlPeOwX+6/Ug4DF7OZ9vok9bFaJxz
bz2RQa2nU6bDs0219TrUbNFM0PqSY0M47QZBcl473BrIvCPxpFPeGHRJbHf6CN+vwC8LlEE9Bm90
FAwP4qH/NDpYC4BgCrKeaqXriAA+edzatbRGnvPNk80Qk5pKPEzdzjBKttaBzV/OnxzyDjrND8EZ
rPAl2p/fAi43G74RRB3kVfNp8cKonk7Sv9J93PqeoMZcUEK2wnX2JZaRKlQndKXB2J5OUyAtqy6Z
aLu57gOa/zcrUhc3QxB6y8c897A91QCv3v6m0aW/cRG23n8quQwOvEgBB7g5Sy8ZXlf21IdBJS4p
3AkFWYtnBf6rMnXaBGydc1tf7uB50tO4IeOnUjXVtCRCHMkg1Xu0d9VUKKpRmVYUfc9mlkMwODO/
v9f1pIFm7t6V0Y9K9er9BzKjsb/YnpdxVN+ouaYUAijpRiqJlEKhtfk3fvT2SJvzkh8+URUijJc+
zR1cZp03XgrAYKCaMZ/tJbPiWoROKIlgHamPNsoKF5g53KlDX5FxeZJsSYf+zTGdQuyLVGUubNX8
dOAOxZMMkXhcw+gzl0sqv86+quTanTpMJwDA7EZzMttZPwJI8uEPFKYrreiut8XbjhMar+nncNpt
1mJXaOlGi0aCCj/mczEOb9K4awp5GtRn30lzWvlPv77jYujM40SB5nzGXus1btbSwnRHXcvxZBB7
nBsOX+xfov8Yk/+CeN4R0bwTg0Tk7TirFDTh1vcHXEg+Q2O5YHRrCcUyP792Y0zwws1m0AfNNNrL
57yIJWNp/rM4HDZcjYr1LDqEkKKtq5eJeTrLOuNczdZTd7N2iLBfkGL+5wdcv2JlnBdz+WDdedcF
Sqe08UyE87qKl6h498YGh6fa90d0refCc7INhUpxEYsHnNeTtbOTkTeuZELBjkiTH5GRP0XWPVTi
IU1r91wu/L6QNTc5IfH+ub6GgotpU0u0jyERRyr+uKBHxc1uM1VTq/eRCzevB+83MnRH1d6xwMcf
b4G0EAmOJmOdae8eJuE77ldQGa7REzP8oWG+9mNKj6FP1ZPAW+YdzOuE0Hy6mCsKrrib5m2CrCfA
hiJl3Qaz3uyUmMEdMHoaULoVCmMKdQZ1926eQS0rAJZrJNMSbph8khzCiIWxn7hbSbRlwP96tf5g
9biXKICNl4oUnSz0w+GUF9Rgtr8nI1SLNaM5W95rLkQgRBRi9fxK2lw9yELhL6XtHgxLmin1NmO3
cEUzOm1kuE47kAr6MzjoEEwpAukSGuBqrkr5D0idYY8ghN7p9jZQmezMxxQFOoupzvqVw8bb03R1
kb9Fu8NiFlFN0INqu5IS4Tw1TB7R7nW8vfz79klsn6caRgvi4h0DQ7vBkTTPS0DALwKfoFi5rZVb
OQSwTegveZV+p70qg42fRfK718GwZTQCfkkP8Hcdz6/0O/S4QxNU6Gv1dnYpdVZYxQfBoXYKnmtd
qgexsYKUxg8ZVttbEJXVbJfbsnA2p8VzH7ZdmCSee6i4YtWcYLe2HYGfhlWFFHuAVEulu+ORRLEE
sjoA3VZz2uaSJnmktzERhHOu38wQUJpRxAZP9ZHSibtZN9m9bki55dqwFLKd4a+Oq+bmReDS6qMk
OcMh4FeGVzDW/i+CXMBSzWWjvmXWO2pr2N8dKNpQmtwpbKztrw9OrzV+LzK1dGpZrETJuQ9g4reE
j/soZ60wtKvu7DO8iehW9PzysSoDnNvspZkdhvcx+vsRES7M98HftKchEgjUXFfx6POmgYqwySFp
Ujpd3LGZpWm9tASPEVbjnumsEKA09JfHxpmqu8954dSAd5xxwmctkniTvwC6KyrvyJ7qRuQ/SRCq
OEDeiu6FJRT1qUURT4S9aQu4x7FpNwJoHhi+6aIcaENSVFrGgA7FFwPLk3YjwjiJ6tfqnpfskxkF
2dxnqw7Lu0NrM8JHqFe5xb95U6gqWot81hCZkKH44bAT1PaaHv2pMDJmCVWdU8U+wRrKc0nTvj9H
F6TBmCvhzOneRgCqlz5wbkcHechAl/N5GAs0B3r2XLVMNcI8MI0gxoP2kLFRqrCtKvfWbEDh/xFJ
p/4Ia1Qkd3o9VIYjFmBt+F1KODsFQZgmcPXkNec5Ny259uwztJvbFMLGO1d9Af3IaEg0LNRckJXh
Suf7FwmolEvC0hrVLtwfrBp5ax9YK4NyxOymQnOObJ+RBzkwfWI1pt95kpDIazcSDu6BVGafF1tM
WsYvB385i6QhOOK8BKPrF1OgvvNq6ROrtG2uVfRHhFcv1mtaRf1Nw8Y7QVGZNzuLwul5CCkQsLIP
VCDoSfewqAtnI9pYKvAK96NrZqUhlYqaIWWT2OQ1FXXX8A5PoVichNJ8d3hyBbFjXsXwG3Rh0Voc
gCuzKVW8esz3RNiU2lmjI+5DRAvnEGyrS0pVxDwcyY8vxp0xCxkmdhSoc+lePY7BsdUILALCgAXv
pNmsiwbdFB+LPNLiBgJWcNSxDgCAi4zaL8+A/Qg7xl0ehg8QptqGBIFZIQ/Xk9sMGxDQcaOgmZRr
BaPEMmvMGgV8owdPitbYK+28y3OMaLm120kwFcCpEpmncSNvSRHwFhYGlWdwWmKyH36YXOSBopNi
ANQH+xlkqIA7EcAm+sQ/R7yolt8NJq58Dy4o8aoyOpDHsOHPeCIkZU7t36Cs/Jfi+VG2NAotDcYY
5tDIB/k9HtC/VsVR2NYNFzNAFHwO/5F8q06NIAK5PKFBYh9nSzZUQDzWTcf0F2X6Yh/vvE4FfANt
DSpiLbBehh/xdOOTeOcNE9i1FOg/e2yjVdjRVf2D0pXuZrFtqivBGLZexRQjvrytXYudmzBigbVG
dnx9COPUrNb6DmCf1jb+nXyIBnvV365Esr1epDg3RAkG570BfCUcU3A3G3NGGNcLyV5/YYp9ep5H
E3JIWKFbRLiYApqcltm3JPd9a4yRZxpZHGAriVILqmAPNYR9OBPc8YT7HAkzrvgjLqYyfyGLvP6V
UaSTTRsxgu2PBPWjbQ4YKYp18rB9lzBy7/0SdWadFYEztnGiEvQzpLun+rGzwy70+MLfgvLfq8zs
8XKeUDp9ZrQ8ol8aMDrfdfp6pP8cUMGem2GOj0vV9wRX23UrnV9qmV98ThlqzLbFqbBzRmLSccK3
pDd1M5XrCDFb0IZYJ6eCqVRV+qJILR50yL7Qdo0lpNJ+oq1FsY8TKjhap8PyKYC9RB9LMTnklMxq
rHu2L4D3Gog5GNetilEA+38We4kt2NPA++ZigtRu/W1ZZAnQq+JqCp7gKJULYIB+v14jI/SMlevV
JptD3cBQQcMHgXeEm6fk8NBcSjlHLyYPBNEXW3rXXqHbcSSg18ltta8GZMoGKG20b74BYYwwSUVi
aTUX/QOfVtnuJmAmmU3d+xO4EfJ6UJ+Tj2UjXPcXLV6CoHqLrSLi4n6gv6A8KKv99T+0gsP/ZBbv
0m2ifrWcRzGlixD0JuLfBxzEAJ0Gk/4N3Hwr0Dzi3H4XHx4UXRsmPVtk6sCdPzLoeZxWxQo+943l
66YOiTM7/TB5DWt54dcgFbhqPzge8OhK55znHV6pjgCrRABUskz/3bRcywn9ql38KngkEL4LUjC4
CujEd8RHzk4P6i++yjW2UMuoN4eyaIBO9uGA1gOV/xzjOpMVIX5tAEhxw1P2McCkodlB/Q09uPD9
JJPLtRrQ/a2/gFYmbTxAAAM8FZrMbN/mL5qGDPDA5w22Fgt3yanVM3O8pn3XzE6DAPaZq/YfszKB
MjyBJtslc5JYvXtZfPQlY/WomfnV8hAxnT/I/pqoRh9seitzOXvGQcLiNCSHVChtFAvWNwTP79DS
FXPvDw0c0CG3HqYEN9DXA05Lf2XKAFdpEJaZsoxHJrGz49EfCo9G5sg9cZLkdnottEzCLzA/F/Y1
A0dA6wPM41NaVgTEDRDLIgTC1SwvyLFWcxo7vxfDiwYVXVW9VIjqb+7fViY2WVbd2osYXNR+j38t
1poRD4PtwlgZ3WWRHWNZ3DsT2mjPb8afj4yGJe2vNIl6/R0ylC3Vp9Zkjxv/NtLXZ7Zu9y5QqXHi
CEH5wlZ6tcA9FxNCN43339GjTtrlcpUyykjR1R3eUgViOC3d1TGpHHzaZIy8I5NXY8cjWtSCorAD
V5DZ90/rg+DLBU/OOOD9X8gjSDKhtPJZmB23WuA/QaqYJ++so6sVXJw18Xyz+BzrOcBbvS03kBZN
DTLlJCYhWPLM8uw9NcEI2O0C69vxXr4RdEEPniIwXgB0lP4bbDVPJLodEZnBxOR9W4euEbCE04T0
WScpNwnPH6RZq12RZsEAX4uC58dRnpYU0TRjXfdIdV4zfMhoIMu/nDLA9BQAimoksG82Ms0XQw6I
EncIMuUwWuoOEGMZGD2l766+WERiqqnRU6Nv/is0294KfuqmGdCVj5ZP8X56e8s+m/1DZRU19u1f
zkwFxtpWHtvU8Z8ZVbwHvCED/CjDQDCIui9pg7TvdQo+QbDQF9O54kTrArD4ywyQKFknmukDTPKv
GuDul2IcTRPq36udshFI1V2DEVzPgNcNyJ8YWfdsGznHV+Wejxx5/IlafG70H575+P3PkxtS/9H+
rmHSgmvhMDZQkMRduAV50dutTREgDlhLovXPhIEBkSeIwyC0mo9z/Sa48pTUQrAEndwk+3SSEFNZ
u4JEGF7mjVCpdZPBX7VgUdiSjyYkMi/vCEscpX8NuF8/IwKdfYC6/v4dgC54c4V/YbmqEiTcihUP
oa2DkwuLTdkJz+vPjDAwLOISwG48lrtiEZybwnBQmFlu2Wnx/t86dpHkEyj079Z+/M2um+XCq6/L
ptcVFcOfF3JINFCBuwXdZgDs6zwOAN2eW1oddq3eYX7oemhaipLEsp0zn1xldlqTt12zPLRWeQzv
bTW57J4BCkU77EIcAjK/Mj7jh8E9jp3JrBVNnVB5UhlyBTtWi6vQWbCEZbbivzjWaTj/R5Qn/vlK
/5XjPRElnskm1VaMvzTBAXzo7P5CEFZI7ljbq70Dqncrbc9cjNSmg67CpQ8TG4q70Oyt3wgZrAdm
P4pGSU3XZPdcG8EkeHw7N9wTr20i7xAt7jSZdEyiwVviLi6jl1rH+K1ZgFsJtMSJXYHP7+rBVBMB
v91uMwxQ/pjVnrgkWTGZThR9aoKC1dQHUj9bSkKU7jkQbwiD1x9edZ3SUS4cbRtartwJctgTw6NW
G6BWgQi7q/hicU9NaKhEqbSK32DS9HCik0ORBoGLH0SmAbleKlpUbsl7XqfmVLD88/28G4zRwLdF
qEDp69nu5H3xmwK75Dn0hB5odhKNafUQ62mdCncz/emDJN2lKxic1F8n914tZMHOCqq+V4SrKtPh
0oWuTbCYM32YSb3rPgTSbLL7QieMmdNLbEdbpPWFTGcKmRfkcjHSidtqILJZSYfevlj/cbLZA27N
Qn1DXQ5kmMtxmTRijG6XyHji9hJu4b2AjdcwhAb0+Vv3x7RHrbea/JSkFSP4g+GYgR8pE6i4uoRD
OQ75RFwwGViZ6MtFmQsxBTRIxFJxbe2yyhDusoqiYfdRH4JlRHabes6uzmVj3wgLFsp+Jkq2m2eu
yNqFdUeW3JFZvy/n74/HtX+st/4mNLRJYPgw6BBAFdnuuxSmLayMwafysyz3VWQZbcciR3ZvVspt
QkBLpDBd3K7dUNEG6ukez6zf1rPWZ6qfla0KEfIYi8+1XSC+7CcbJito140j1OxIz5+uHBoIsuY9
v2inbg1D6cg57S+DVQFKAbjRHSBLp2eAuk/8mTsvPBxNuGLGVTL5TnLWewbd7jjR0yvnyNs6rMY6
bu9jwDEmzusQ+qHsIJcuvrPSdfejWzppYckWL5gDgdJKHJnJ9kh2AQhwSjkBZ6hU3E/mEpMEaXgt
fzhCiniQ45QSkvJmP62tJaWBfth9kSQUP0RD69P2nNYx3UL/zQHLDXPIA38xw72NNEvkGUd/JtwN
7hutePD5Cv6GxdpeYVAknxcxUq665LazqHwaDr+lmze7FWIghw7/MkYcMzFCyI4od6Bv+WsDkgHB
rCs6LOb0NWjHzHrxY8LyR8nVF9Z9ATY1fW8FJLi328+whoNAhrC7Rc2HbAa7MTtC0W+Q+qKG6+uW
B8dLtY4yl86/ytjILLW7q95JHZ6/VU4eQG3fDbdo14GtMDrIDwGVDJJOynaxwXc2AhqrdIoQDsk2
VbGMiWMtGUx2SKYYYd+5sqAfEYu/Huni3AGV8V7mDI7AFDT2awJvUwTNMgiruExSBi0+5uXw2nev
bvDUGNYiZ3UlLVUmP9Z2nOLLYWXz7RgcjFpHbhVkA6bI+EMLq8NY4iLxAKNvAunK+sgDkw/8Ozs9
gDaWBrVzsB2R4wJjQvmnb87oZ83gnf5w0bsaILLjAliDqNC5mIeVw1h0+JIqFS4kkmw6p2LoM+Av
sY+nEZbPvlEA3+SXDLR+NqxRPwOupLEPHUVnhpu/vq9BIP9pIsNa0mLXM6+NQPDpXNzY6q8MKGGN
EFsfprKun8zuB5Cxqv+XmvbrDe0vb9anKoSuuOo/jeq4IsNd7Jbg+QlyjkltRSCFRZ9ZpK3scRmn
p+By54tM3az1xqyW90AeMRILYvRPqbZ2iMp6DvWoR9HHuXP/efuqipJ5LdCYnsoDHphrf12WqUep
lTwLW86b8TBjzPMcLr3qbuup0mWDjFnGx9CVNbb82q2pUrDBG4+k/7QUfv6HYFmK3I+TovYJLs97
LWcLuXbOzTUqv0YgcU+FmX4j7YuAd0I08uWlqEvvuu7JoNARPmhTE5bU5754z9VzepzgjtX5DqJi
4Bzl8x/qPyF603ipO1AP2UXhFUEW7xGzeNFzne4Sxn0JkfRYRNivwGdZL0Zrr5nizyal5FgmWUs4
+1sDP8m5+MiIK7trP85UktWCihyToh70t3gMw/aLbjfvxnjW+bO6X9fMxDeUvNcnHwCQ+cwvpHC7
YZlokejEy/lJlhKJnoKLhl9lJ15G7+J6S63vAxubuHYzirNhrjDLpoemPKVu5lBLHDGX0XdVHCcn
m6P2IsPdZYFQglgkyYN9jYigN1MSiuBwP2Br83tUtBr3k2vX6g0SpKqLrC/wos6WW9blSEBYjBN/
3An0aq9Hsgo5yDpejIsqHWI9IPgJ8pnvqQ3c85S5uWvygzXtLtHKCJB7qFpTVxRhddMkecCHtySu
A8tsT8gch4+9emwPIbk57NWaL6TVVh08hTJKa4YlXaxsPnQPyA7nlcIq5UcwD+TM0prTf/rMt8En
/Wc08rVYntuWC9Ffnse8wy0Zv4Eyrju8Uwrjq6DoZ3oolN4ziyN75mx/diNs97kIjJErYt0BBMbg
wHBYtO7zfPGlRmpfP3vsPtqwWhWLX8z1d55p897HRregnFygHFlHtXgEjuPfn4CW5FjRh4DBEDDr
77ixZjFIGhSLU0NQJLj5xZblPf19zyZDUyNgfTICzb7KCWY3vVAvQDjWWRT2NCG8xgmOfxZ9cN2c
bhePcl2Tdj40rXDttMMpr0j0UIoswysPHirJ5djxovYq1UGEh+EyNiFWDzkd2mBiqb5HQaoOz8z6
U5I8kyk9cjO39DQxM+EZALkFqgsQaHxiJtojvbAG0+VzJqA8JgxrxabtPnea3tj9rfPKYHdEf1aA
kx8Lo0F4IR0KdeSLJj8/qYZSXKOTcNkk3bYCdnmUawO12NosCLl4dEW6EFERYyvXijoaSVt2aLap
eCyn3bprSlT4N7LRjmxezVyNiOh7P9AaJQrv/J3es5fRRMf4DxSsZVHKxa9UYK7SJGAkzndq+UxE
spopNi1cObBMOqPjdiumzW28z3PoIdvmWe+SpnkKnB8VmHN5Czio2vdGITeTLJWD07Uw3SY+pkUp
+S65HLsixfJIUmXhDn2EU29sxQ67PWQKQRY+7XQ3T+kRlL4q4787KQ2nOdEdgjExKXG5tLb9g2G1
x2JZ7p/QRXa5YEmS2ePbRSgqBlankC64AY7UrqnPqDaBnxdXGGXXG1+fL5+KipfM/369HCldpjjJ
wFSsGVG4ACiwLnVSHhJxMEYa6lXkJU5vq0AKk+H2B3zmnrOxfQ9UifmNzjOEQzpzL920RfuYJ4HD
nclSzjP4DJ0Ah4DciluCmItL/UvAEs67AiaSiEgU9+qMY03LjVBumgn9SH/7HT01VzENcFqibKfh
bMtykLZOE3jZ+qIhXBnVINsd2bS4KWg/fXBS6lkehykYW5E+Pawnk7Mv1ZNeRBn6/3Dct0MLl1eN
0tl6IkrbS4Q5e3bfl7RAnm/go32cwDsBpnIhGd2o9GGu5C9Cuti/tygCMwbs0dikNJTGdHqAT/d5
QPPXVOhU3YPpHWaaJnzIcAhyCkNymDR74p1Cji82FCnqnZPgQjZQNUca7SirazcRS2AS9GGaJySz
uE5zn/0H1emrWm06AGYkn5PSIUIBjizRVo5HV8Ph5Z5G6XAxmKXs57N92AUj+wp6P6yWXvGukD5H
dVpfsBpkac8/T//rEOvKoxFq/nN58O1KgwPgMf1v/kun+fIlf6R+Ogpz03aTacqDFwh+AcDnrAgB
b48LXpU+bKmEGmHNyA6DfKBGGzqXqYGX7Yxta1wkkGI31itGj//dW1+Omzs0U77R1bI1ey4QV+PT
/97mEoQ1dqRAhIJ9wjdBQHmexR6RIqa2b3L8AKoSozWJCBKQLImF5taSPitT1112TpND2Por9eKK
KR0MR1TIxxRHTQhKg685Pw3/IS1TaJ0xaVNajYVf2gqQJerh/WZDQU5uNfiTC1yIpzAeiVLbs8dr
Dbp7rVHhiWWEc3nejSXmskiF0p/5Z5dJokpU1wUd3y96dysjnWDpNALklp7Ij//pjHaYSylEvRbh
Jjd+nYgqxd2tjh8EUJH0C76akAvbvDsZi0jyQ9qF0oWRWTqREJP1nlqdv2p3k5/qRGzsPechnHkE
qBow3v5I7nSTgaFRDzApPRnCpncKwFYhr/RdJszLbjvnwnggOJkBz/67qkSdg8OD83M1l2ApVoH5
QbHVJ5VezxYlEPnuMktTTSmQwZrvnRY6689+fD15rQrlvvB23zi4Z/XDRZzwqxmR4aiXqwUdzNzO
A97B2jce/mTYHKfF0dszszrB/sRjMno4m8dgMmgk8Q7lNGZUDRNVr/gY7Su9Zx9yXdOG+v3fJueN
f+imHAj9p0UbsSQCv5EuBGHhtY9lhu8w+NNe9QgMHJq+rRZl7bz1TY5rKJ8nTq1E8pfSjhqo3/75
i282wFFnXPKr9S7q3g49XrCNGxztA/EYHMaE6/j3xamyinrYfm35zUmbeIkf/mdQhYv6Wo5qqt60
LSN5D5R+eVvE2iFyMHAB9f1K3lbU6LSQkfoDrboTDwDUEic4XvJVDGUVVSrOEsXo6RMvv4s6Y5m8
PI1fLwO+L6JcGWVeQ81sG9W7FJ/5Tx05L7mYuJFXzqXQmzVGFO9apSBECw0lu9PegGsIL0J0yrAb
pRHoM9OoNEeasS3zOeV0e5/rhY5hOa+WePeZzdDwYoc1a8elwdNzCgZ8pPcTtvis9PmCc9vcR//Y
veIG48excNFcB5m7vkpMQbkzOnb3Q7jlFMOBiR752BmU9t1dFHqadLw8J4Iw9TjWt6g9kv8XFk3H
TE8a0dqNi6+0qnQ4efrzqtxYikqtyxihyUft+rEUKoV5NKObW4jzs/EOJxTT6US+9GtBEzia9E60
0Iu6SRXYE8w7myrn5kwehWFniqPx6j/3QMlsmdeWqdfWzdOMt5XNwaf4T9t9FY8HLju+KIqeYUHx
ljw7sk+H69XKmFRE9MZhrvUC0Qn/iAadrcfVmH8C5t3hSWitzO34fFhT6XrGJHiHpU6laRVpRCiL
HSSdofxHXWe+ySFmi/CL4RVZXpNRbYRojHL/GNUc2InCWLR+YH2zaDincMyEX9iGgtewDMg/owdi
R/4f9qe10OGszRItQ0dUR92MBsTu7dZQ+hA1yUwaTookh7yT5eDTy3pWjDG/gzsP3K28auqz4Kwg
6ModYJEH2IRJkxgcxsATtzG43kVM0lJ/A3wnHhMmTOc7yWNMcZRSfgLO/dWNPY4Zc+w4z5h7+E/o
/5rXd86HcCd2Xw0lg3yCm9vTXy+1rQVl0OV1QqnSP0asbXlpLQAgAeELuQ+qH/+OaH0Nkd/u1MCf
bugc4hl6/Fwp3SPbdyz/9xszViXD3WUt1iPvvQYA7Qlh+um+uEbfK6+vKXxdPHrlAUtVtO6U+Bgt
JW+ocTJiP4z2IvoFgAYhaIV44/3I6W8W5ceEoN3fHBgOdXsk8Pa/wYYtBHef5FS58Mqicewpv/p3
PqbsrWBxF/LVmconHGPE2Khf9dlL9sIm5QzwS0FkkPrA673S45OvcT39uMNdtFBUd87qeXBeMOSp
/gwEe8FiyjCDnY5UaNGoVbUuLAcG2IBXZNx9le2x95wrFNo3EJMjiufEfIYliC8nJ/XUfXkwCYw7
U8SWLcS9weHknhbt1F8/A7HpiYhNOG80xZShFvwenjzzSsi3pzl8DY6eLP/Rxs3H+oIF3oQyRaNh
gVhL56Bk7NCaH9A5xVCtyVUr8xdCPcoNUijMJJh4iMVaOqKeS/XTQ838TPzSwj5WtKKrpDytqqq3
WdM+SON17wa9HOLuWkmAJ+GqaSPQVdfF39jhpyRFDldteDHRP/hdL4N9OK5H5jKLNbdP/lrl7vIs
6sSZ3Tjlt3sWKa4xskkkDL6xs00QsitWFCLgh7eosy8AFtvF3xEbkGTmJYpFu/DIHCcXQauzkEwl
dVLIXQhEOdGDX/HUh8Opo1ZaXiIykHrgdyBew3LWQqtKRMuETwJIDM4nwTfwAaRqIVkiXX3cfdba
VdKkfltMkVUbY4izufKBWxjQpi3Nl8L61V5wHLUPamSmhHxL9a26Zp0Ec7OVOhSqc0FUFpVHsDtB
OeVpEB+nEqctN1gm37WBt/Xbij4sOZ2a7gUm8OuZcSe43eRVmiVgnofe4Mia6jRj2xSig9uBq3gQ
AH1ZxmJWJ0fFstb9u1xH8gZLhKMm8NncbOveEyp7xKgKzZcHLct4DRRAWuZcDXOiYtank7TmcMRb
YIJSKUnReFk0fKj0n12F8qx1wNsR8iRP/PoaftimEqjPMzIvZwNmH5LxBDzhbqBUITqmhp7b4+Pc
7OzWfyN1+JlZL92XoIit2H1lV3SGzp4qEILHa6PxoiuP1HOFkoAmw2u1ngmkTBsKfcNd9w6JPMLO
t5VUYegbL8nEVXAlpnwTzbOUriH9Cx9iTexBmiU97Pz350Xn0Fzrq8P1Vku19SrnY4C3VlXY0upJ
hT1SccOSVeEIKJUx/C8gPqRf5XCYwX9rvGNHiHQ2MvOvxPsVTrRNmU0HLl39YjfrSp83bsjY7nOt
vWa08nuaWoSlHN1sFIWi+pq79hRzzPkoQHo2cmocKG+1kcFYkyG4zzx/tSklrAEnvfuYXsfc7zQu
ODTFBHcuG3C2AbunXGC0P0zq/w3gYQd4EBGbKxQVhRfpkL12GpftjBaZLy6YLUXka/oz8Drd8LO8
sA55jznI+h2jFqgpqVIiYzbwLOqCKIyv82AyRLRz/0mjqqKfq4JyfhlXQWu9AOcC5DQ2vzqHVmSv
i+2ubne4rjR9fTgKlXzVPswxHmseZ3pCowTXs7UM6mvEtmDJ2eBcqHeFUe615I9N1E4+nDJk0g8B
s89HJn/xYGn1xj7JKQhRXLCMdL8Qv/ushqkog6qXigHIIrR3jqJPz56fpDRWVdvhKxxUBLO1RlT0
9g+ZuprVVNUTKz81LU702dyEEueOxWHsD+7AvsvSBobyH5CTfZicp4jeYpxq0gpRJpzPZVF0SkJF
Ao/hx5AfhOvZLcypmnN8byX40PDZT0ZTtnnm19ew5ZeQlk6Zrs6EXpqYQmKf218xu0hDF9T8m8+s
UIgOXeS5glNRlS3u4LoQOJBNkOD6hq43oHskNAzwTEJRgNXdIsdghFW3YQ7DP5X78u860UUkgOcM
+Vlm50+ENXw+b5prIoKrkwpOpi3gH4feCYtVvXkZ5SHMIW33pANDObduBKxMH4eHdOzrZPb9smq4
h/B9x02mqQsl1aF4WzV3wBv1LqctSYPCLFU9YtkTc0O/SJXPoFdM/13WAbjZCgTz9CCOYc+4joF+
oiZ2jlF6TdyR2TQFcuq2pkYOOQOBBBijM3HJk0DmYaMJm1Xlz8tN6SnOFhk1Q41kU6lxT7YeWmE2
L7Ff4ZDpB2jW0l/NAksWWFNoMqKNtzqdQpPsWzXUFANGbCZrWIhVkrcSTHTr72V0ayWfNwqqBrrl
OsHZoJMfBs9sCyOsFtCih5IEnN6QkCXaPYw92E0tgBDgUW/W3kOruxWH4/xJRqVYA+k7KsdiIZx4
FtD9PKHvZhQ1vWfLrhSZtyKBCfhNezT90gstimQj6C1EgQfsNLdQgmJkol6Ta+85ya6WPwtj+C4p
01VQgG0rjSZNqQmqh5ikhIRkeVoqUuiTdfTBNAWmhSNWdDjULONFVO5gqc4lFzLxWsSWI2G28IcH
o7abG6v7JamIRYqR9vFawJygejul5ecOnqZxMDJ/IHx1GIG1tEM0v2yqGmoY/K6OFMgsRLMRzJXD
C8vDjtHJ02SZnu36ZEXOVLjgZohzltMI0+FVsCWw8aRGtHaLY1MnyR1ikfgqJV7Cayihmq4UzP5x
Sn/xkm6hAwhyC2ED7kndpCvGdliTYflmMdybOnCVoUp6E5vgV3bPeiURt/N3BLwIbQDTZ/UOpa+C
EkodzsirffX4c6bJNxay+jI7oMMixRKfpFwBUjbqBIK8dRmnaUbEmFtCYp7lh1kEm1NAI1gWopP2
zZw1I2HL3SopCrnsktumRtIFNrKjLMdKoA4kND+qn1H/KEtalyPguRZ9WLppi3ODmvin+yiiG0Sf
rB4oT+D2R3/I1qAaLe+3D9aVwn214f2XbC7oAjRnMqBgxQjvEKdyOEEhykm9AfpqajJXuO4jmFi3
u1mBPydRrkme+/l/wRDqyVAOkNl6MK0X4FsYH0nNa/KKNhnteVEehcWb6FQ5J5/oXwjs8FRPnsxk
L9MUpb3nGfn64biR4zM3QrSRoTetPYd9CyvK3RgwF8NaKLvvWybDwc1DllgFie/aocqmPf8S+hb6
Lev8zb6whXI2fP2z4E9E4OxJ1bHlMxZbp9HXwLcYefVf0vIFl7cV1isuGy3ng5iw4KNXXm16BWcJ
izvecC7YKymM/wr9ROzqxF66kNOIlWObNTXRLo8Se34bLsJ7hHwKTpLGs7RhWAvoUAcdtlGwd3rr
XbZRbJBM8vZUozqy8T+2vdFYhPA7YqjTzcWkYdA+oLxD67ej+HERlTN4DOyWL7E1qh//fr6/ZmIW
gVnBnhbxQqBx+YZPRimqapviyIJfBarWn8DVZkGImSK9DsiXZVCCPP+XaKpUeMff/hM0thc28Tnu
tphUYdEe19sSsHaA9LHthuzBzp3CUZ49OqAdqDdDs533KiN3KEgJxAQt4GNFwRsdxKP3lp7FNKEY
IpSTQhbGQG5S3BQ6jsggNOcOFnAgwkmZVoCnRuUp9J4ajgg9ik2KlsOFRZ5MZb/beWBpX7VLe8Kh
9Kt6BRRJqvKhRwDI+rLr9gj6VMBe4g1xWM/xzm05aOfV7q8yGAIah3FF9QwlVbHZ9P/BIK+rxr8e
CExEDBAN2w3NOc91bJCp1cPWxA3kztCSe7gBuAk8pTs5iy3TXrLvCQpRiRdyhX1uVx4Nxh5kPsvh
+e4bTMu5+DV5GeQbl2LGuUY0xIAGSSa0rz/RYUpsytHKdy1fifeDtR6UKRS6jR/el+biLTH9G4Eq
tTmLuzq8vHrc4mP9zsCfcB6n6qj3Ja7YM/BuvacJjIQGQnrxpzpu6UY+Ha0dWLNA9j1EAyAJ2UVO
iI8Ug3+5V9Mhgry/VV9jPASzIIOqUf3PNDTMdbSu7TqrP6F/dKNmz+CVYf9a/n0IUL8uiEaJBiGx
rIuX7qV7yP0AXzK2pbqFWo5mu/vctEsGDc4y31rqMKZDJETZBHC0qAUPi1eRonlET7zAYadk9XEV
YRHTMoxpeFEZP+KYxZfQakqtNZBJRUp1M7/Aca5i/BzL1hPSEXOzudcZg9cKUDxERROO9mqZeGUO
49CNCz00vN/NqmAfced74uMblQoSmVekdx6yVCAA7bVVX1eL3VMtuzo/nWBdFYVUwvKWg7SWQLpi
aH53AtEtgnCYHZb5AGX9aCEjQ7Pg2xayC6h2dtnSVI0rqaOtdk2u0DOSDzbe2hJGmxhvvx/lJddT
d/EXfK/bI4CJet1PgKSXH3HDHdIBw+rc+24nIREhPICpDdWl7whkgH29wgzlDjnh7VKcgTrDAdLR
aN6q8D8dVK8D954+QdT0IFWaTzyVpfUPiKV7JFgoNmaNVeVLcrd8nNuOTTx7LcXurQxi6f+UNLmu
59NJXYQog1Ubj1tC/YSq6rmNUVRTVjtaVIBWNRp6KtwAUAdh2sJhm2xZt0WyJF8ei7aS2MqtNBc/
b5wxx+DVNfwo7vs8PFSeuWnkRPguQecTHpN8yKT/F2zfbX9UYyQI+gEMStvPphis82hTkLhPB8Zd
xdEnJyRXeNQ8gPhYQ/qzVvXCZTWn9SPVfhjCDClhEFUunfjaLwAJ8xC7mvOfJAfqcrqV6eAXWdn6
izeT4Y+lveR5cs+yPZ6fJ/AXU0qkr2Q0h6vyARSw4U+Koa/XjZvr7aFkFvBZcn2GXsJm7EygHLAZ
tXua3wASe3EtleJw37zgKPKhAOaVNhOriLrWivEzXhOK1lXkTA26Sy7u2cYutNaStHpNVmVF3/jn
mlXHI7t2vtXE90LTHru8kDIuMwZ1BkJStm4wnAsnk/6rnbx7cR1tOzAmblyINosybJS9o+peQ4sk
+8Onb8GkAQAl25g/SxoKUVewPdQL8XF/JCQ0oLihRAid2Z+/q7AowA5s2las1OJ/AMNkRyJzk0nl
FTxveN/bw0D8+hHpB9Zf+yUyuCODA9P+xnfEDoY+Hkq6OENedBqK7uNpTUcctZVCKHvZoNU+LoZd
c8ElVMoEdo7GKlGGtboCJRrmwlsHcW4KKLkrTZmvaDXyQJ3zu/YWzH1r6aNw1DshY0hfUE6aYwwt
nAPe64fAJBzBC2somg71EKOIfG116kArUWw700Q4etolB8XP5639wlk2exCMYmsQ2i/mFV1bUzzm
wqw42Ly+gZxRrEelnAcKglbuQKc/d4a9gwN3ijnJVaSh68Eih0IG3QdftiSV9tQfyDeePjrsnFGf
rOdMZEypv8zZ/hW1oOfc7vdWHTynMMN0L8AXD0Q+IoRHoRzf/CS4leP6sVmtDIe+3MzmcUjnwRZ4
sP/oZtsj7pZ3r7HNHNakztDPGhay1gSRES0izu7dIL95FSv6+bHgPaK+/PifRkd6BEl1tpfdbM+a
qhRvm4uUQHOW/8WwiPMdMi2VmTcoX6n4c8U0mK/JM1gHZqjEmSyb2JUH/lmKmIcyKv3F3ubXZuSr
9pgpo/kE35/SOYk9EU0F9U9hBlscgy1j93SJ8dsnqe9L8f8MtMzZrsbLvdMXrvs13Om2JWAZY+Le
LTpHmahuNGqmJ+OvQRHjZb8bUde3Ggfjg1L+oxWtIEaffHFigJfjZ5Vd+ErkiaaDClfg2yYhyWK6
i5Q+mxduuFWZJH+P3KE/GA5AyQ1MaVlCrvBvMebmpH4SIHVI++n5rfCSZZebdZGtVWqYmoPaRTdi
3o4UrakOWNZEpq2/iLBHDrsE8lguYdYkwOyb2LbG8dw8mks2GOHTNNnLFdl21QP/4Ii1NeB893cW
vV2aZcd8607U7adPyoD7FqjjoWr869wPViLrnk7J1YtK2prKacJ0TQPNshA4S62B7I8yME7YGN9K
3PlfEb7uRakaArGDDUDNCWwrceV4OTv1VG9WYp+KTJndzbc0azTwlTVw/AiXDaxcvVRrxiCXBJUR
79qVkbPivDyUcMh8zvx+m70a45msWqecK/0R9mliE9lDiSAnZ0qsHRSIXJt2wJbzWRemWvP4wtwu
uXBixpaAFSQETxGiK2DwyS88x27YiKsZGrIs8iKJA9RLTGjR4XasiZMdPcgFjYBGFVTKFyKEyjNw
VWAhD5ujUQezicWSdEi/7BBv40qH8Y3zwl8oCEgz5reWpmDwvolfDMr0E1O0Gofk3aPq9qkQbfIF
aobuhdkV+EcDvpH8TKfUuPg8o7hLSrUVFPq5TAeS9XBqUW6SoXpxVgIyOIXZPfrdkp7FA3IGhUQ/
RNs6FGCWaSM6bFK2XXcuOl0ebT+weqolV7MdqOXa6wIzLe7iNAisswRl5O18FXmw1UP8piKzFF5h
AfkBLtN2S4UkIu9qI9+iNQpz5C92wkqMXFra34sQ2NVAb8DIMxgBdDUTJqQ5xs/7Rt0HZS99bBR1
42ePqGCbcBRs+I91Mv38H5XpoRoskJRtnrnK/PVQt29f6QsGP/8FIq0P4O74nEp+2fcE05+vRUGj
9lRynTKBN1hbq9zhJLosMM56JLw4nF8KUnwn3N++ZUXtj72EF2umH/61RE6BXJfBgTqMiZskYPQr
aoUpUNS/eUA3zx5zppd9tqQ97Zz1iyZVxIfOZ7GK2rVZGZ1cDdeYKqkw+sNqfIlugWZ2kr1dDO5k
neLx7BwDTKFY+JiCwrX4Ho/7eWde5JEvmckpEnirUIqcrl7Jr+mzSZPEfKAHVl8Fc4hGYCWQapnk
eo9MB1gAaluj+0RyHc1sneU3oh1JKXZlORMWsFbTaq4fnOTuZLfzQJ+2MOs+hz2fW4yZLAQt+mf4
Xj5hu1OK6Uye/QIOu62IkbfSofoL+vH1zy+djMyqZasTDPjTxPjgq87M1FsuRUz9O0XsozSkzx/f
IeuN4D5u7b77v4PN/uCTa83J5NwMzBr5AZZtVt6XHe4f/gZ59Zg7KQqIp9RyWxZSabi8Y3aIaR/R
LQxSpnWDa4JxnbSo5Vd7gfgmM4EZxIz0vqL5g7BQmXarANiufydPytdSWJK+puA6AUJ1V78uMVri
Ssilk6a1mLipt9kZBzJibwksRKersQegzNCk/YO0uombfXn0/CtA5rU4hYPRIvAetFPqMhOaPwsi
UNDG57Vrg9qmk02aFStw64wSrEuGq+AFRlTP+9HemvjyxdsPKBUmPr/wvUtkqQzCHJqlgZAujfqO
YT7vtCsF5w6jet0EajwSu3Yp9qmgG0gTxxmzPmAwcQy5PXgAksbAeNNzmIB3yzqdGHrRMzgg0yzo
85z0BK25nB96n8j9Q+FvMHeALScwNo/a1RUY4MJkxTav2dLhtw9CCyNqPID3fPBQgbCe/B33PY6r
/iiRrx27bN1Y98bSTPxFAzRf+TyIjcnTc2fyIKIa1823ta9Ihs9v4qKJ0MgSFDqzspNOjXmxIYCX
lcTI/eg/NEqhcLhNBjs8LVRNJw0O+UzgbHDOPFCgrXmmKya3zXzAjGyZZhMvHuQEe35n3gYHS11m
OCUlCIBRE2C/a7UTHYNuYsMkksuWG4DFU+yl4jH7dWZc4Skh0iOoDUDz0LQ+sy1SJc5N23uZayuH
YPap817CWS/r9c5JQkYuF2eLsZTvkxr683oNt3AMvB4pWd0uhw8yLffWeJ4WMVz7fYXXOsgdvAiX
BfV8LPakJqLoWpo8t+JuLK5JEhWjHN+uxD7IAuwPwrYj2/tV6o9/1E+i69pALhV4j+Sks2efBWdq
PWp1p9x4oWw4ogLxhtsLhfLiDMSA9b82svb8VyhxV6SUtclFnxUmvg76fTF0OCCPF/xbPM/Gba3N
GmfFwpXb+/4Lap9aI2K8AJeXVxJZj7YFxQA76iwpllgSXv0bqtGvi7ifu7zR0flMNqTxKT34ELal
tSMmw9pLfyAuOoz9f+G673R8Vcjumo8jtlmh523wMDhf83CCUMvfY4wKhTteyZpy8E+dotwqoLyL
0TmRYQBi6+PwB0zL7rFZNnOWHVIk5cJTSkaIcfiJr8L4fhNKevbIrt5etBbRkmYBDKpRhZRZVFqb
vk/Dk6F288YRGlQs6IRYjK6TLfRc1csij+lQ0rNytWRCI5+qfnwBM2andBDlEFvJGYOcOnFSimVj
5Bh95AyFXmqeaM+JUdePcwPdg6bC6rEzR13e1I4le8SufIIZyONzzj+Hffvw/vv/K/aGr7zb+GYJ
w0riN080rN+I7rUh2DEVlwrKstuVudQ25g9SmelUV60Rj4+8ZLykdlUrbel61qpT5j5E5Sb0AIWt
Gt9cJOX37v+EsoH+m1SiNttor3nwurGKj5/UCZNSiFp4cVDmXYVsgHrjAQlPydUIyHeIeLK8dprP
jd1q7RVmOzgmX297R3df1DzFit40FeztCLE9hjEBtycziS99M/MinaWtdw+QE14xapqgj4j5UrJS
wOCWhJXEVEXGWDSdhCqQmtcmtZpuMyijwVxcsesOUEijsIZLGsDo9geJhzG+vJTA7Hi7VmeLtB+W
fOHIrMYGVBh1xNwM1NGXEZBXEg8BBaLNzJpLns5DLqzmmJNA0ji+xx3qzQo/JpZbh2uuXhssjzIK
lnPZo+b8DuNK2qJJ2Lglp4bD0un8asSgOPR3jWTlWsBqUhx2TE/EMjfBdfVHotgnX0pCx9rbxLPD
pYjALQb0WH0C2sziI2huNtMDGs2aVdeW65sZ6KbDvEn0jcPIU4UJ0JRqTdU8zqFS61lXR0S1SICs
uW+oMlNj2dYnnM4kRl4VCaKMoQc58D90qmcsv7vgalqg5C/lautSA36BEYSzfibSImd6q8Q+7hgA
o5THxrKBLex2Dl7A3j4PE253jY4zFt6Aa4j5QTji4Mm+2sIJGAQE66aE+Qu09Whvhm05ZdY1UN+z
CgFDcmB1LwG92ny+QljK5YYH5I4P5QBwELC2XwhYrmG80fEWDYOPf8i8/uoI1YEHoAH0PiUGCbW5
rV1bhNZq8wNCQIc3x8KT/bLQ2Z/TmpbrRbJtU3c2twHO+TQL8M6rXfEBc9/HSVgc6oapO9cFZcGn
FcwzL5kPN8dVl4KrtTblmGmWW7B9LsUU8gKy1Sq2RhcuZuJ10kxEHjn3KX0vHPmvbQ+EmsMpZjM1
tIHr7JlcAxoVhZyj+3sBxcFMzYJlTqAOArjx5hh/rMuOpT+M54L5IKI7O9r7rARSzRHsSqD71fha
67/41biq33PzT+1OS3BCOL8/0VpKjr1JyzHRN42ukZRB206YJCRVX9GTMRZOor2osDBpTsrIbp5t
rJbNIkhZF41/SQ5YNrfZPb0ILNRerrNmepW3g26eUqFGlOIyPxI+Lhtf5Z6LsZ9AuJpULQOi8DQQ
b6VHymR1oAgc9Cd1WzXmktQOlDGC/9D03ysHtKEuJ78rEtws14K/c7rrPboIT7d8eKW61gHao1jm
C8mnPAgXUcrayC4W6ZTVsD/Ou86bqgITIWICixFL2cNtA5kU90ABgfr297Sd7Pi9DVgGddGm6+cK
P5wJFO2v4L9MTdCJuxuESB9ekdwBpTTGkqZHNt4mowqCFccQv3fIW6tonSYncFbGzfRaMcuCT3G1
YTzy/N5paFhSeKyKO+rY5GBfQ8ndlgDpTH26gbZRrrbjgJYKz3V0caJZ+4WPoRyPNKpJ0m2KFg3t
xkQUR4gao1U2DU6htk3qjftZ2V41zBl/e7tcFB9XCdWRCuY8T/6dQYk8KgZ2FSnxnCVbNW2YWqUB
FrwKScIhxdWpVDseyOF3fhF9YXfdU2hksIBvQQyp5Gb09LIfG5HPSQAolAhDpE8JH6Ki1O6yO6WX
28/nVj9KQ9S6sP2dO4R3jezIcjBj3QHJon4LAn1anjB8GYXvkip6MkFySTFxmsXbUQwpT2UBupXb
49DzfXC24wI6YhGJy/MWhhJUSbl39C1e+jGOituXs9JgFhuPUQo3+nXJ0cv0eMgTkmX3xMzIZhUW
7gImwNA1ejJ3xt8denarV4IDnfm8/EpOdDNZSde2bbVPjJ6IFVU3Qw2SDV++hN8skwjB1oFkgCgV
CROlUQ2hmtAdjvoW2wHzrvWwt5qfSSAsNQomTXR2cA1Wi3Dz2cke2SYyhewGmuIjlByaz24NurMZ
u80T0FHVda6qVU8dWn6pHnzdasc1lbsyTQH+g2M35xln8CTNtM0L0IAucqS2SmKwhErxGfKSI/Zc
mIstxnb+pnNLm/KrogMBR63513CEu+v4rD5BBz4rf8XUQcli6TuXQ6E/Y3hqptj1kxwcLMFnK0R4
qQesnoYv10bZJaJMaf+wCCV4ddmQ6swZ3C1qu4ShlaSXayKNYvw1qMr2jzpB3STAnEHjbULta6TB
x22QEHle+jdrBiZg1dbPbFkJJ2M88j/D/Fqwdk+BxNC8LTL0uTn65niXT1feWtidaxaYi8D+8kbK
Iz/td0iEu82n8+gDEBt1mBbybjwa5mSzs2TKhZDlfh4hhfXD1IMQrtpXVHg6VScTe/iFgmT/xrRH
Fj7iXmDyebLuymnyz2xbz0JB5XP7jzdnu4O9vhHS73bP82L0pOG3T/NIaiwptMTEkXi4YvpOu72l
5UHBweXfyzcmy/ODKrYSVymdEVS1yo+VZn9m0Vs8l2KMGyENWQt7pB1bltONK401Ec2VHjMgp8pk
z4f7Bst732n/uH0cpOImfiL1ZYwtWhLc15/PV70tkmbKK9ZYwceV3KXllX3pp0+6F3FxGdDNW2U9
aIC3o0ocW7rC/965/EoGmMYukAAHpC45iqh6+pNjkX6zc0msk/Iki3WiJpJ6vsIzrViW3cSU+Iyr
ukyULkRcAx8I4ZQdWUN1qz9XQlNOjRQS4bWZbu/5PhO9ff3msBLX8nxv31kUJi1Z27ixmTSID+wo
1Zq7Iwh1QBnRTTJMCuge4LR6KHGiuGqSyz+YAtlbeAw6n29m5n2KOpu6+Az9p+gcNZuf2KiviQ7v
nbhfZpOR05f6kXrzVYWvnHSF2oSvfYW4IRow7UZLaqb/AlLhuTWB6gg3M1PC7yKWB5k0rhixB1kK
jF1AfdFDMky2pGTcyGUTdp++zuvHN8Cn0AgKkFY9BFiMnk15TmDF4Dfx0lkocEDNxMMDLJTrBqlh
hcRC5OOhOP5KHR7NQSFXyYbEbH0ldClWk8WjI9D4K8OOM5uyY9aYSuiS63FEZMQq/RMmMRjX3nEa
4Tkcq0KTe8LMKWCyxILoFMzk7z9PydIXHpnLxiSSveMrph9S8JK34MGjOv3K5HbVK/4d0BK36xqa
ubyzSAqszqytkas8f6bnNpqC1FzYO8lMH7IPIuHHmONvFP0hnj1sWasWdDcQmjIR4Zzyaz6YoqL/
XV+E4ziJzXOi66lkrRlTq6zFyAosaDKNlIVvl1Ch24IVA2jECI5UpCHpA/5sxO53mm4iir4di+4N
wQJAp97Ne37H7S5tp9ScHJTyslYMXtlQOwBXryeKH+nchHkmtGJDiOy4KXWPGgszx2vvOCpLK/+g
073U6/4wY7TG1Cq9g0/ouicGClAjRhKwbN09vDdpSh6Rvs/5wZECtXUYU05DfTtqLrYWYv2H6q36
DGv2KkyuYlRQibDqgxKqGoGfqzCSJkUQD22AYXx4bj06OlPHSrf4fBbxp0/gIgLUXd/Cr5bXOLHQ
nTDWYSw8qAYaJ4yX1GSs2Li3FOFV4JC9TsJhuTzQpphzbzKbmJBZ8kwZ8PusVno4DYthy5DUuw3I
XxCLhNGyyXcATXGby8SWeuRHAsgW+SxjatAKPQdZdlb+TlTvk30wa5Rz4cgo597r9Y+YBz4wjNTp
DIV/6+wjXSQ6u65AR6MbwHsnJlH2uKkbHTjiZVSOwg2EjcRBNUdWyLz0LDnXNj5wSzETLRQ54iUW
XyeOv7tl5xDQNlH6+17cd1ohg/muK6w5PEqHV69BbacA9ZypRtALsAugZaBhfpIiV+dz94wzk2TD
bbcfgMmBz0ZLeks9a95OP2IAcz1PVkneB8Jqt+mTP7SZ9i/KN5vSmXjhtzMgvCPCoAufCrXyRv53
8EvBsHvXy7IfT3Sd1X1QnBztag/jMgefDx5vON6s4OeVEOBPFFC5DyFrA0AqVZxWKmxjAsOvD7vI
hmIb2+v4ZNHDp1n+3ajSJHWMC7HO0h3505xgXZIbNFALlf8xXWkJhZxj/pMn3VtNQiefsuzOUg+q
P7v/Yo8Q5CcTwoOVL3K5C2/KYC62ezKJZYhls1H072A0xnA0c/ruUYarrXZsUdWXHQ/DOfhX2TYu
PdNFw+HYqi3eY+T7LO94hu8yEXTlfng74JD/e9sudqTZ+16PsKFT25TSCo9R3XzkC+3T970/2tNu
653FfMoijrHmsiYL7kZomGMBOu+XvYfjLhyVK+yV8dgtt4GH3F5Hso6GUUD94wMZNJwUZ+aLjXj1
sYjLDNZjEASz/GTB08wJbdQCmKLpi5McUNjSLWkwiSVHT09G35J7Ub8PazCW5Wdptm5fSJAz1Oth
/cfjuLFgLn1U4zY+cdthjj0TPoC4M2QpbCNMHWDGAmKdBAn5Dh8+fTaKtwbD+JO/c6iuAJX9LLmv
cbfMe1LZPo2+1DFtqgBGLDUvOPvU3xB/+PZhmtMK9HZLZGUN0qlvCboQUVWPUk8fLgldndwh/HtD
LgrUpw2hxNB198FKOgyEdgTx4ER1rstbL9F71gGrPS6ox0swDPpi+lzGNb97SY3VVcZiSX5nHQAq
BwAjYdhtrxldOn7gaD/6+jgMxAR181Ni7OkEYKfw3Bc80u+Ge6EcpRQxSMDnPOXj53+BFZgZ0IYC
5MU1awDAc83yTF4xA/sPgK35MXT6ABiqDY6maO5wM7gzC2GAAKeO4238NImYqeFSld7KoE+PiK0l
/VZy5dXytEH8x0wN7fKEQ8qpaWh1RkNzjkoOeRwViHh51yKMJ7sw9RF5RiTEdhBKnCdB2uYfXVAw
w2lP4Eizn60t+DMZzTxcd4ikyzlxYyIyXpcV++Xz65qtUC+pLPaEjXuqofMMfS6s1bW+ZBTrwG2U
yN/zpSMpoUyzrhYfichBq6iv80C6XOLlMoC5G9r9Gyl1jidMbi0J4ZPLyOkj/EdqfAReWA48fgT7
KKUSSEfIk/aMsTWirLLnWI0xpHxZEdxLigkflGdQiyWZctOHJju4uqVfmoVa5gykXVMHDlm+yYK0
8Mq+Qh+26yoWIcOl4ioExAeg1g6avRZq4DXS+7dL8nykfdVpSQ9Q7CnKd2MyLs2hS7dNsHAfTxG/
LahQY5FgEfSdVzutoQaTLOEnqq+0LoBps8uopeYbL8kGJHGQm9fB0EXKLSW/mDWopRX63T6tMEnH
zPrSjxZLCULggyKfPwfX0EnWPJMC7KVUb73F+RBzGEQqPzvBR9RQtU+WNhsLtAfXph16207hdPtT
WAzi9GaxIQ7MO2Q1WJRRlARAP1tx0xjX4JoEPaJTph2q/VH4LpsgfMFSCnosgM51KGINk52Il+m5
I+T3o9lSodyUQO+pvwXnwwz8IShwgjDGmGYVMLRdo2MKCgLxrexwA8EbU1mjMYoPqLQG1rW1/JWL
2ZrTa6QrS4pXDPqVsem9FhqkauGUJEeK77NUnX8rUf9oamq1qj1+XKaPJdgviI4z6AKAM7ylXWIA
JxxH2CEZSz++Dw5LzjV53/tkWtNN+unr9uZB0OslrDdTAq4+IEWLDYE20aW/sq6cX0+OAY6PTGUu
IM+n8NIRtwd+7gnVd4Xm+iL9CkDdbYTCtxMwD3RMIez303XQ/D73LQp82JYAfVQjuBp5u8Ul145S
qzRNmMx14Xka6BYk1GG+lN5de3JD6HIf3pvNC0l+syg37ecbUSBNIsCHaUCB+fFon/S4LGHjLc1e
wrAERYOCIxsIDN1T/1LCVYLqNDreu8RNnONrmYK4uwEK7n8XR4a3y4FkVZocIrxHNvhsMNjWghM/
eALAQO29BOgpgw9gBA5G3s3iaX0OB3FLzGAXFiJHZkzALBL0EmwL9MxEBUJKnSJc/SdeLTe3txeY
zhewvMk+U/OgE5s3rxIvPpu1gpgP9Suvy8CMeHB3I8/VL1uuAt71Csv3GR2DOMG9wvsEZsu5gmbn
k+pHUBjqLpgfrZvstIw2G94+6rBCO8WSnMtKeNfNmNFiBl6r8Q/EpEgLG9YjvDo86mENpdcBCF9v
iCeeVndwV2lyo5r8oAOxBT2oTlt9Qb8vin9d21JqHgbahz60F3sgqnHxRSco8PHBjwD3pTtg7haS
wM06J9jwGkrGWzLxuR5dUJX8OiwRnGIlFTP5v0961CLc8ajh5k4CDGR7aPkDupguWL9+a1CaSP4n
gs2iC7NGBnmV/6kj03UxPdUJmm1VAQV0DLPsf/9wCSuayEL5ogbDWHU0libqg9185THk0ALrcHGk
3xpa93DkS7wVEweI98IxE9qNtJt0XZGC+KDBz3gZHTIlfuPAaLMknKQN1ORofhq/PCv6AnhKHFfz
w9OBejfDyDU6XTLBH0gKjghO7inyqWPb6hkVsYjxgSWdHRduFkb5Q1IWUBqhVcuUhYqPx5ZxG+2c
MEzGgbYxI2vypUOX4apLxINR6yDi6RTlpl9Vv9NfWb5FDocqtEhjnCsXohQqzR569z9eaXX8zEUY
xpUCKqSIp4kUIcL1WKc04af6SkN5N5dgcCbhiaRezsUTeV6duVOzs6KhJV7PLkLKqlgdf9/R8unh
HwRw5gyHSpxlqF4QOrdsPfmVp9aikN3qHafTFSIgYkQslzVexHd+vEtLtVkj5vRyRYT4jqSrDdLv
ymLBngr0QZxEu1mUz7b2dcG6L10mvB3qHZ2vtN/IFMIJt/UUSual1TaSJ9tOMRsdwRkJ2CZZRDXu
bXVKQDs0zvwxTCbymjYtoY/7b/7y/z0MRF2hTugUz6CkYI6Ygv5ydwDhsDwM0Gq1VqSjue/MRn01
16LIT9XPUHznUI/CfYTpzxfOTOxWWmQAvxgFx3r15MHuj0Kmc/uExr8j/4gbGDmmjLeGC/+Y9oHN
F9B+2dcUI7dOdlJ9wFK8Ndd/mUkPSgssunrQW+BB5Z7e0GbgaEij21EXQTlb+JhazpdC4VuKyql9
7SnxbEbsgeos3NOZBTL0N+XRSQeQRCQmNBbWvuBun/aHA/FgjM8cJ8ihzEIh28VRo4pIgrvocogr
cD6t9xXTTLnO8iqB2tmNcBmeRVDhzqWmQDl1q26pV8bPoghMmE89N+X2I/Jl7NQnn2jzwQQAx/TE
rgRd0Q6sbOMdkbVBMjURCRG17RrHOae9piiGyC7E68THI/Mezxb2zUI2wataNW2+6kkimDGdV05p
hTK55fULnvq+hOk2+4zkJg4GsYsdpttSZLC3pp1dydrF5u/ctvBpTo3q+YZK/NkAJaVw5dRfuPGi
7ZQGnSJhTjluQ+e2h4Ol4mFIDD2s+GxBkjzw+3pf9nTBdoV/8JZzAdRmD6I9R15tzz1aoNgaMCAS
8zu3mK8/8rp1KSOwXtJCXeKafc845nHLPbGCu85HxJ7bcRkjwF1KBPBdEhthm5TuUHQokK1YL6cn
YPKRb2n041dptzuwE+G/t4r9WvaDuCbGx+ey18J9b8KMfysbezceQ7iWObwjmJ9c7Nfo8shQ0u63
ZFrVOrx/y93JPnEhlFsgbT6lzJ6eiaQNtUES+vEMI0wCCki3Gd1zQvS+apuaTlpKojtdOrni2jn+
3YqnHWO3Xn5gPRYCiT/51C3/+zc7wWNs5bcb80Q3kZMHQei2gVmHMLO9npF37p99+chiZ2Nz9FpD
tIilihYxOcRw/7FRqZmAIE22tHLNo+S0A9XXA9UtTGKd0OS4C0L5ootY9gDtBAdX3w2hgBpEKdIj
jmV0nQIPoQ3zF2P4jq1UCOP1gdUj1TOfs0K3Kn9aK6k8m4skuozxNARwabPEUns5ooh5bBe/+Me3
WzesnamgL2lNbQu2XvADXC0zmp9IuISlBTj7nbEXnjSTvA4RrmdwknE62K1mb5WfhnccnASqG3JR
W75rU9msrseAKx1Uvdr6xjuLpOcctIE/aDNg7+fWXp4DaJvm9s4QDkp4rAYL+ud5N1YyM3nFdjSc
XllHqvJrdXxREP533Pvf3h18qOQ09XHpX9F5YqadvPtBB2qfPDDzaZYf/5YIdIshuLqtVvYByw1Q
0chkS5IgrpmH6UJco7Y91UOPnaZ62lYq+MZN+EG56vf/Crb7Lh7XVm4etQMINXIPjO1QJaMOpVWp
8Gol/2DbwFbwx/3t7E1STbeZgK+36S1Ehunm/ZiucR+ZNn2BmNd+5rflNuJCeFLlheUIpiBhwj1x
hsD8lP1VzZ527b8/Y5Zqb4+Y7DAPBDlULaq29cNirBb0RLtNYPXz3pYLX8MZnHWj1uTC9qhvR7bY
J9hR1VMI+E7MIHXUaQ7W68lV1tbl9izF2zzHeaFtVYBm0/+4rVsApcQ7OzN3ArERHGlcYLWBFxfx
02A5h+NUcgcVpXDnOtm0Glktwiiqzo168L9kUfJHSc2hGY7kZh4eetna3WQwsdKT8IPaIJIuvYHM
TPb8RNMMmbbuozPF3PtH5Qbq7h9Pq49cCtF1AlHueAWAwPXcvTPQLBNM9KzVnm5aJq1KXJeRPQJX
Pv0c9c8YJQTFOCsjVPz0x+oR1vdOz9U7Iq06ZRVa4QUAZfUWtD/oHCWIOAIkEYmYi03uE18rw3y/
eqXC5kRrWdbAS7YX1OWycio5FPgrkNk3diotaOHvmr0zN06IUos1P4pOVKn/i4zlrP1FcjVcY80F
zT4fFLgyTR9mw259A3j+v6LfJUMk4wXyJUdY6E/WQRea3Q6Ehgr75Ab945t0SsKgIRJhEEyE5wYY
WaOeqIyoMgUy+mlU/axO6wwvZQ97bXM+pPl2fdP+/R/W02gjAHMKL4rqjhhM6BWfgpzFjbH1UaEj
Ba/RlrX4xS3RYH7NT+lMeC1qmPlwL31Gi5Uh4R0X1l80IPW+fXfa+V2k83rIhtOq4xX+CPRxsOwz
zjXtQedIJxT+xAX6/41d2cFQsNnpq+IzDbJ9g9QV1opWN/IyV8hpJpQi4A0R4Fg+d/8bwEayxakL
TGU2/FmOlrPLPq/xXriDvND99xD+Dmv+AaSeHpzNseXlwKHwr1FS+4EjQ6yE2dWl56HhTqjNsImd
brYdu7WzMNbAnKk4wjVYvH/qS890EYbJtPwNjkPysf+GH3Y7Fzb5IMKkB/XWFn4QrcpRa2x4NN/i
f9MgHS2eumA2j8G9bSafkVcVlqYtnusnYqqgHOFhCfzUlLm+OHPdLaSTjdTYvo4kNtgv0Zl9Xodf
LnmZMcbNPkmDwxDx7c7UmS5AOpO1msOcXHEM98zd7T4Zzn/eY5LbbREepA/OmpvcuMHZxlbM42Yr
LBOBR3YJJUAcXFEIO/oRt4qxtdUNv9waQyeWVn1Y31nsO/kULzUh8A+pbJH5N8RKh6QKYdcKQk2U
X9SypO9RISTZsf5klF6icSpaLmhSufSh+QX5ngjhxdQ/M87Ar58lrb6PvwjBQbNsE6Av4fE96GFx
aT7ElHq+YFfxeVeAZ2a1hgbp+OKx5QywsgBKxuQuC35BUx+FV2OCPqJsClGZD1NxIHCk/gKev5N5
SraNOet+yNfwp5LC4udr5mNofS9/Bb0qE96iBbw6xc/Ts9vTDcHOZnPhXepVoQIbNc3NYBJGmC0p
qjWV8FtyZBWLZlecbuTr71wHP4SAoJK17QgwCAQ6GpDcjFy/m+xOBxJbbji9QxAG/eWZIXUJfqhh
2q2to76C6WXPQM+yboM8qyRsu0Vpv218eUHHXJ6D6LCBEKQ46ADIsQe0U2ei0Et3affyQYdqChT9
v1VdOiosmJffNRvu/+h2aMeXTUdSFtgJQsJeK9v2dIEv+bEdqujsK9cMPhzIjf2u1wYcLQWlsS6Y
selIj9tRx71VCyOeX6DYAKXlL4FIZphCuEVI5kZOyeFU6+9p0haGDoZd6YzFoFneY/nCyPc9U5aq
MM8pmhaCaQYyXB/fUSOHVLQD444O/wH7VPRpVQ2VTXzrN/T7RZzbAJWzTOtyq1KgRGLnKkwcy+n4
pmlhhOYgWmrsKPurhmDuMb15oRn7kmAkTOpW3aQe6Xb4gMlbCdYDohp/k+qCurpDJNjRmxMhgNSX
Eo7pcky9g/hqU5fJ3b+DfE2rmhjBFEt41+iCO9Hx7NJphrBPowtH7NOjW4Qq7z9Nmw9R42h2zKaJ
kej+pM5M8l52auNEVl2bxbhYDKMRCYgnQSE7jWrkTyOZx+v9xezNDrQyvOG147ZyQx4gNibLLLJt
2gCC9GTEFlqzsArBRQii0HaI3wmQXPn0/oiawcCH6btfbFAEIkoeULaW+ePEa7Kay6v3ZOLP5/bq
RSXjHjzTTsknUQxL8ssMM/5QqyIcFBI1WUl6dpbCavM7Dqb2V3Lb2JsUc4XdJJRbFcVj1unNj1ki
2eg6Kpogbv1vVLXs9Ob9e8AgLmux0odPxR592E1i4p+0Zm9lU6J5Qz2L6qlbBu08iFIFYzX4Y7OP
mjqYOTgbXNKvtAf7MZoeotiR5UvfLbgqh0JSm17tGzZBzgEp7UP/OENIwFohbEz6JNKEeHOefkz0
jv9OKnupxdF2ma6/CZPJ1KA7LjPck8JVhH4cydMgv+x22NxxJwJcHIO86NliNbDpB7qwWSWFgEf8
kQAu+xMg57l+2P9HWl0Y+DjTTMm2OpArBTmWQNDGhRX6xthJXnKY5w97qLllXBQp+8O+IXahAGCP
WwjmHGSdB6g51mVCLDTDpxEKaoux8bGdxpJ1kfC4g7YQMSVK6cQ7I4IEd9GNhgj9QctpJyCmKm92
oCtG2CU5ljejmkaNJuQlpRQUNvXkIdVa3D979FglNGd6yvvjVDvOniqHpjrNvqziBOuAxZLBLwr7
FJObrljLe+34eSJ/dCK+WaU8oNLgaap4eoiSiruFVV5zYraAK2hZDb1VFSSgIO3gKWAqpGm2ezcn
604R5UxCn0Ksom1XTau0ALdp7N4i1PytO9OJKXSITrTLCnQXJWk1Mdsss9ps1/u+UBOxT06907F/
a1oQjSIV4VvrmY7FMuGWU9Hc+fjBMpjwHhJEQMJNjhXUqVWVeOCMJ3kC92buzSQWqgvwPx5jGjKg
6djkxYZ0BiRtBmGU5Mmo3YQCnQgK+HRbi5CLxIGGKN6VCB/E8EhI5h3qbSM5bu5EbIjsN9sbSfTw
OiXw0NtV2Z91dzMNeUeKiQR3fO/GWR/vQStQUmb5Ws2vHIr/Wgu/I8t/4MfnhrNNXNigLr8EluYh
GKcU+hL7Ky7m1Srzv7sjUWKeXIgp27Bmg9TBGjLPZjCPLDB0ZIFWrwV+EYIy62wb8a//E8hyr38a
yg/GCFjRWBmbIgraMOhQNIAbn7g7zltNyVqfx5wBECcDBosHX4QZcqAnOTQ4LHtPF7BMeYFHhVPW
hKwevyszyyNVKtrpiABDlexsqQnKQrV02LJruTK0xcyIG0KiOIVrRp/JVsdWDQoBUsfQx3uCwqnb
r5NYvB/jkeX1oAFN5GyS2HKFdDK0Mf9ei74n4+rr6mjLRgDPXvRE/wTehbo6pHiJMgFpA+uJ9HFk
ZSOIISaGfYykfH+uRQxbjo7VwlsFD1luVHKtRvC/W4TBJ5ny0FhYZoJtHMOZkLc0/opHNsJo4gec
xAAqO8UVURr2QhpUtvrdle//cQ8IZh9eYp0byDyJ6BexJbGAlqHTLefoOUB/LzGY1FcQmSuvxZN+
+su2j2yl3emGsToUfTiInLpfrZK+lSkibp4OUfZUBSMVstG8bVpoII/U6i8+Z4Ah265Qn9ZXK2/a
+hN/jTKuT+glQYPDJcxBlcUlhEbE7sdZ/D3o5CD1yeiC8O2cPUbeJzphD+5XhTqfykHYNnQOUWgH
giRnfR4DueRMUokpLE7jDfdMio4vutC+ur0eyuvQCp1EaMWQcZckwfRsGPdVIwhBedCpXhlxa9Dy
M50GTYK9e8W22T+2WP0eJJy8Fr6/lPHFk4PL32J11EKXmnG0Bwfzmr4t9dOHvaYt3rmZy6x6uWrY
n2JtM8AiwTx5YyWBJfkdO0v3V8kpg1JlPVwQwFhRkYBCbwxpnI6xK3e4qZy4jcFSxICgVWA6svyR
L3u5P+EFGqKaq5QJFYLo9rTob3u9nKZzuBXG/ITEYvx8f3+IALRvjQc9dEDmgaj7SjQYygniKftA
vTYgVYaSDoIIEZPs0OTspVM57MIHcASbZwpjdPSZI/hCNRcnkGvbLpbJOwlXesZXhIrCfVuUed8O
ZJZIH4sTtCJhDSgXnCodU/gjxvqvrgKgC5u/e2Hdoi9L8Fx7TBZVW7rkSckaOGGQ8j6+Wez34nbM
Trbk3IIQgxhlA9EpKolqd7GjjJo+paM+6lrdSrYjt9GAtvsg8WDw5QGf7RVOqYWXCNTnfICImjeQ
iAqdvOW0oEdQXJXSiHEhRsRBEc//9z8yB+MAyph/xtlctTmNObxSGee/MTQee+OXTSsBdTSxeQ6D
MQQ7/PFMVdQkrpuIVTnqBNTlM8dA3d99edh3sBxv5l66+/Ue02BXPHJ8xRL0BItJsMjXc0pfXKhr
9F/stqJAlXiIchZ+h3Ic2DPxLZQNc2DRS7NCjzA/pm6jFu08yC+xf2c0Fh6UtJ03uUlRmH7SQb0u
Pppv6AjyWLSODff3yy4XOtFEN/ss0SJhSBrCjhCIkLb3Z0xaeMCyT7rQpXnd4DgF0QcPA8UMS4Fk
kMNIAeHiX2mZitglkylfqLQKOyjcsYAZ1unfWnVizGJqBW4y+8838s1wEcCstRJteIq+Z1ovfThb
uyUkl+r3t93lPgG40OLWGViBGNykcgwAere0N44An4HLtlDKVTOYQ4pOimDQdFEJpX9X2dxtxuPH
KiygbqypAZHRNdPzpC6VX6GZBiUDo5YwHP9rdk95a9MX2LAZl6fu5dXU3mElAEaAd2ThxHn/MFmC
xnoe1c9sYYMYWVWy58SsyI7kFEcFrHWhiFlBb3Tpp13FRrb8CAUDEa/jpyHgkG1Wem8iUk8v4E3z
We+E+YKgO3mHmqni+bzy9aK6IuERwg0b2h1yyo8STsBuYIJWj1am/Mecf/vjy9LrAynXP/xRHVbd
dQ/ufZ7CmoI3loWgZxEoPPtYNW2oGfWy7L6taKlNZSOsM3P+ia+MYEbHew9nMs/y0PM/448UtbMs
/uKYBiAIgBBU6y7E/OCnkkrBagpZbJ8jt/oPTSaSw72edVHxv8wk6/8v69hAz+pODxCg0pdVZu7x
QnLRzwhS4ZvRabR4Mgtmp1TGZj8lrJ1t6uOsJ4QyiCMCznd9lO8x9dssRe8qOY705IC2kB7pE54T
oGO+TeVL7cMKMVixCuaTOobrj6z8H7ch9kEHQ4TLgPVYaHE7hwFV8nYe8U0DxqgcU3bjUKp1c7A0
ePCjP3wcQtWn4K4jrRuZpv7FT9ODqe+V8o1tX8gU/9WG8SZoUULFsmxO/1si8AEEDb9Yu3XhbMr6
lWHsbJPcf8TsKi/PoKtW/Pk8d/aZ1aiy7Wlv4VW80GOWBCkRoDowANUZDtcFKZGP7zYk9oFIfUhZ
N0M/vYK+O+n3CCTLgNgWzRzy4Ze4omyavMwSuD/PWoaSYA5+eWTxkKErpto12p3U6RfQ8g/9P1np
NZgKeQRgTlQTqD4ZxkQ7hdayudT0pr51T5lrBAGGWbPlPCT3+QrHP3pIsFo8l9XjBBy9qFfYNg+b
tVh+g8jlPfl/+vbo/vrT7F6CQNf1e7OScvw48jFriLB31GbMhLattRe9UFgzXUmo4m74n0/m8Hd/
bsZjNEujdG2m6DVxi4et/au6DKIuiMP5RttzmJSP3xBJBNgThlSebp2/c+XtGgWeNfkSDfe6/c1l
wxrBUvJ9u1XT1mfyicKfkM+HsJTA0syLZw0LbVMPFeVlFYJ5LNN8uycnW/DUh8TzX5/RyWtVfsw7
wuKpPQMbMCG0g7dht07xNqBZ2W7TBbGSjEqcENQRzJPQM3w290hxMu7RXH9ZI7ujBvzqjmny0jcS
BuGS3upSvVZDEke1GB08lIcSFspgWBJumBMjMciBW8prcQCcw1GXYQLDYK5UnFLmtEEsDftArqEI
1FnJozGgofXTwo2E01H7dxS5wQcfNGhKmqtUtgoPHkGXZRwSx0SosH2nPPo64Pdh+ZFF46izcsHo
3vKRXI9FBDn6BtvBXOstXXA6TBL4yRHB7zynfwCkOvgeha70YGnQsYAwT3E6nodhPeDpMn9FJ/ha
Xe7BEZXBHI9sFlH+YMqdSpxt95AzPSvoR1CkxqSgBdjFaseGNooO960YGlr1YrWwMsz/vKYND8No
X0LI/La547Qf9CIYz+NYu3QbaCxlIlnmks6eexE89Hplfklz2/gmfoG+paC1zo/EaE0dsoy+2Dy6
QJMxiMurfv/T0m1WeAOfEgqwMGdt+wWrDCpY1bMw4rdpgc4BCNKEt4FHH2jegqv7P2toExdRRU78
HU0WA/WHggvviGzXYNXrly2tFpu5nMJHLgq1nfRw4E//dGSeJJzolD6/T7MQ3rrY5WjFzwdwlZv+
cfERZ5xsl8jqKcg3T9JunsLi/L9c1VyXzBAb9SltxP/iJesiiof+ZgqO2SKUugn2xNOgkrfO7w2A
rNp1rAcdHSYXEDt8NemHJH74OVChYxm7kjBH+7zcPZMo1+RG9t74cN6Jpd87X/Hobuc8nWJQQT3I
CfeslT430cc7LqxI2GuvzH4uNW2jzZE/4UmB9gUSufn6CdD5QX6bzEP/YZEs2hcuBo1tlJDA2ZB+
eIcL5e+tzlSRt4APtFR1/JhNB8jv+zTpuhHXyZAGaYuV03wbmi2FvFO+WNBqyDMa2//zQkPevst4
VHde8B8TkkspPcVdNg6O2tzyCSJ4BGHUC/uGzEYqSljcuLiKOtHbvKA4uw73dwZEATOvlDv5NsKd
9ge3lwisD2utxGKx9hVPlrU8mI2Z/qKvAbrVtBp7po80RqqwJu6tw6EA7V8VCEh1y+Xup0EDRvLL
cwCrduryVgTRPR5fs6YmnGxEpnTm2KvvXIoAk8iy382XKtjh63P6C2hppyqxdgVbVto0ieWJRjUf
lUMWcrFdxwwK71Wafap1lA60HTWLgBmXgzl/j0allDVnyS1SjCJCUnJxVj5FjwH01e/THz2xjjWV
1sDTLoCNpUtAbysEaG0Ww2tSKK+qDrnJ5sMm9ET3n5H2v/qOclJd8LIFgKkCbzNQMMsE4KBB48D2
Nzqoaj1Ve6H06RePOY8a0kafi4AEE80O5qcNxGAvu6gqH4USXUk8xWKHD/I3ENYKgF1IwsB9+NFo
HpEjXs5hkQYf55WqlBXWzoIe9w2hT4F58edc0K860kLkVWlhGE3FMRkBKDww92WhS/qhG7ceYQG3
E08fyQ7ISvOTXQtNjCvp0JcnYeyahQE4Ncn+2Q3NK8uJH4j9uh6rzE9aOKgU+CUNOCmR5kzSdCj3
wus22l9CVe7sl6zdB0Jlgn/yHkJTZB7rA3IVXOjnPmqV9PA0t297xjPme2KhDT3szEE5Jnr9+3Di
pZmgq9S2ALV41QHLUybxZK5yM9iRJNgbiR2jzYeqiSIFe1WMZEbmxJtri0ld7LU39sXvDCSnMtlR
EAnr8qJB1BlBQuEe7lQpkbqZPKA4p411f/ShTB2hQDDln/6bASXssVgebzR530XdSbgGPN4gPYhQ
SBVAgNtMWE0RyTU1Y54JJ3bnwZ+QwIAYP5z/lfPCHgwlHoM1Cf/w70zFhSkqjprJ1kSJMWhPc81g
cKAMiIdocig1dFRDHleXMKOHwcZKs66sT8NI/VISThxF4HQJ6ht9edXRhPrPqYAO00w5PBd2Pf0A
ST+fqDVnnuFtMBrbvB6d18tI//EeL9vISjWi1L6acwIPopIzCg3nHvaGyNJsV65TMoPBUS1OYVIo
N4RggLBAYTdo9geaun12mSmJ8nx3+biXXNRdY/Uz6kukB0f0I2XLkCiaisF5AI5stzd4H/p7bzgp
SKxwdV7RvXgkteqcVw52GwjsUvKxquB2uZ7NHy1FIfzgDkFx7yNF0Bkd1VGOeoepTHtCVFT0069B
B5M0FEOtqeoCgURFfdqniY7mIGG2gigk1FbHhXw4Tu/ItEPeoNYvIiJUPWfnCuAubDoCeTgW2+1O
1NkuXHs6rfKW3fqIRQQqMbxTa84X2LDFE4SZG8VxyGvTexKnVXN8nVs8escUbEIRlnYtCZ+NFKLE
YvYwTmlBo5PgXMrl0tlRxP3NUt/Zea8FyyoKXNrUkk3ltVRGRO1WDOg692mRSswFatqpOtKCx94I
cE3n6f7/RdeD8HAAX5BiQZ01/lfdIpmMYqLY22V6WOhwgHDlmxZXTCm/032crK85KBdraYCzRzEY
NwfPGIWrAEbKx30uC/PkOsiW0kIVaCR2EfojqAAS1mdif3U5dNJuV6+H9jnpmZ5IRqMjBs11VFuT
T3pksrd1Vik91XSGxWzNszhGktd59HoaJiOyR1c4Qodko+HqPnVFrTRazapyANXRwmRNpUP/1Hr0
j5YfSAScxuLYs4OnDx/mgGQnkfqm4ES/nSGLnWRJBrC1hPLM0ww2cziUrWAp3co10T2oIbhIEd+G
4mYry76VhYDBtcodax4cgJPSDSdYjNraG7tCRyss0fhNPRxtUMPluGIqjzmMDizeAAUwU8FK2dNt
o6ekhPBxP7DwcPLGQATUG64hTRbpQU56tJ37GNBgEMivHE/5TJ6XiR689z7n73JAsIb0GNAWhl/B
mU1fitSq7Hg/wI8OAUdgbgHoigXNXGtXLCDiyzEEK+Amby/pwKdAcumvNf4oJsRyICde/APK/LvV
orEzngnGeuzyIYIyatpGjCY04ML0WQeYrFtG65t0UQ60BPbJaJ8zhkVDteap0C1ncRI2IhnHV78N
tEP2LscI04OAvP9yyxKHHsNYa5l3vm+16wsZW86MqZzbGAtb8R+SKPdTsMAt6waJk8ffB9e12MQU
lUhwaNDP5vABGZR3mTi14dtgT/KVM0IfRWxgFOXUtS9vh8kzZkeJhanaaioz9e4W4D4TX+MwklIT
R2YLA0tCtF9Fnur9qOahKtZM6h04gZB1LxurguujmLx/6b8+JJAcHAP/dqTjEqUT5ilFPswDBLJo
eLA/dfcstk9/MmkgRGYLVkFCw8DWChuOHlyb8cvM+NU+DOnJ46xeBZ/0wYOts385j+NEPtIw7/EQ
nsOHIxxLukcmPbs+mVvSZcuY527WbJP0j7r5gKzeH7J4Qii4lMLsj4uUuKswp7Jy5SAqvftvcsyM
qs4Um9MrgVsKM3nEgqKzaDW4wkmC49gKoh+bgUu5P0Hn2G3Xbb62IbJroD19acT6UFz7jVzclrAH
QaDr4A31+u1h4B5Dv6EeFDdRVdKhLREEiwOq19AEQLqubSi1Nz1HGec799bVSU/dgt6BynrCFQJu
7AYmRsLjwlv4TGKL+aZm4lK10KpV6Ajyd4Yf7GwosQ35FAUTG4IE3muDqXio89ihS0QYk3U/vUCh
pB+X0Lgg4L1Ev7pv7S7rpoi4ZzJT/ep3VbDOAhiTK10bneEwYYCIzHIuMDjmJ+9CMDLaLWZ5D+P2
yV1KyyYcylNDQychIQfLu6fvsySfqEmegJWSGFP3AMDkVW8OF1nDB/g+eERbKbUnqMe+PInS/Q/B
AKvbz17WC3rj17vuFOZXd/yRdltQI52kMC4OeEiVod59KsC6c4Aqtd+UeKOjy5H7BRQ7qFaXg4cN
JXx1R6dF/3kjbPRZmfNnZvSJiMEizYVSzxqLYRLYum/7fYTnKZE9gcFTNkNDFt5l56FFjch596G9
yGmzYPDYoieEG8dPxC4UY7Yww4huqp/2r0H0NYn4OBdfqeq4TC+FDde2Azn+57PJefl1UCxbzxRI
GWB3cikRnwstMtGa1QG2D4ycXL/4/Lde/cvvIE+sRCECbAEE8tvLeyM8ry64h3qXoP3ghWmdvqEf
tySvY2zLV2oJogd3PMIN95O1bhVL5HfMvZ3RhggAMbBcB/dElbNRAVQ17EUiHngL3jEzpuMHuK2H
1pHJC4BlYeke4wflZ9rwW1Kd/VEaeaiJOMZj1xKeZwANLco1TrbISsE27h9Pzr3vtQRf+Y5JfkFB
hN1BUoK/qVq6HtypIDkTKXS8YYruP68QGxDOTA5takwh8lZtslQTPNqGQSGfc5EovpZagov30wis
slPttxVCWkQjOsrDGYytj7cTA8j4up00aDmizB4Y56x6qWvpRjX8ysZf9iOOtalrwDty7J82FeGg
BcbAAZaWuUDhy8TBsa9CNxz1z1Q0caEjangnQ14AsmDNrK9z79c4XWVAFSHMnwidD0P0OliP8r6q
+SfmO+3UhZeheXvnJLH0Jvve6gvkcrKa4NSOoBq6NZ2vBzYOvTNwzSso4YMJ+0u4AP4czGnqvSWp
GlJGVohdUyhH081sLjijpfqtfkevGcwJPh++6PmvYITrDrOcKRaLXrUp1WeLhLtkFdQztORd9xfr
eCRW1JD5xdZeMvvyg2ZDvJAgz0aNWS21RTrnihn2rSxEHOOlfdRFolfNx+iB3+ltNsIpE4YvypPT
0UwZiclR9GgvwEoCbSWs2icJ/8I/Lkmz/BGFFvy8gEg9RAChwPl4dKgGkztpsGF1Lm3Ek/eRVZMn
k8tyZypW4oM8v8HybYk+F4mvoJj2eRgyQxS1F3oJY91KZI4Dvw+KNaAeYzzxEtciLIvlSKsH+6c2
5HuX89SenJpRg+Pm7wjSzvpJav9UzDsp/7bJ18zdkvULFlmUuKM5EmAyICqh4ODp7PiHkkHv2JRE
6L5lC/YYwKoXB4JIo53Yc2JlxrROFECRLCcjQ/Lkbxaio1xd9n3h6P7KtjH1GHnKtXCqOZyGREdO
BUR/JMjUZGhN5js6FiBC5Rr+599GG0CrqZ38aChJT/6y13j7HnIIsftclp80G/4kKNBao8Zvx45l
oxC9OGeXyOgkLcY9HarsldUuetw0wX0W2yCvnYb/xpneV/SRTCX8HEkyrHvWFQ5J05kPUcgL+Fjy
YPuafpkcz11M/9/gpcAil8g6C4u61UP7Wb0Uflhot9N8rtWy05JyRGcaJ3uUh2J3RGJ5LypZHv0L
DZ5T+wEpSgTX+ic35hPKNv+YlC6ujQ69a8wUHoWynMnu/Tpn/4lFDJkY9TnejxSvFRJBu9Dw20VM
lrhUmseJJ1qsXvhNKQvhnnCtGhmvW3xU+EDxiFrY39LbsorHT/v28YbCUQnh4+iI7TFIYfiHpXie
X69Iv3DjI7+3gjgUgPIojTPQmE9uvQ8o0BPGfCwcsY1sSgZF8gRrHeG1kqZciOb6Pdkm9mSHdZsC
FKql+fulIq5EXhdIYHsUR5CevSbo9NFJNtM/d85T+VoCbpvIg7cklzs+0vStiq0Tdrmp2VMII+lp
ARaeXQJJgKDGGzwY1uDql5sFQvYCOykBMF11FXevymPsnyFKGABUOeiunEOeoGFoxI+GuBvsMtOs
+5+g4sBM8WxVDiQUWCXWIKfQe+X6M6P4/NAoqBPx22Ayrw52LIkqWHPK+8xfDyEozvehmUXX4Yiw
ZgA04WRhe3VdpKuLbwOH2kAeDJwG55RsoSUrHBY4YH1VAQ53I6xLg1dkew2/1oKOHGZn2eGgL/zN
ZQPKwUfGdgv4LW3y8LN6ixIJrzdftqZzEJsgRzx4ccJvPIxaeytpuWeZCte4Js5s56R0bn/RC13p
OXpzwjneS0QsBFXrOMaT1rzrJaeiv5JBlvvlLpUulgcjL5jKrcLkhE6vXQ1YXmQTFGSQyOEwtPiz
SdrRGR79zRQNJvXyu4IBtDxt1SE5NBzxhfXkAH/MqXCkuXNwuyw3fQEsW09ldb/7DLbhiUJGTyS9
QJxRHbMr7g3KQJfxKcJ8nNttPp1ZYMaOIVtDc5uc3uzZOiX6EHAL1LR+LVIpUbFBJl1RaRHclm9E
iEA59cFgCGY0JkcWQUFlizCb7pabKRHAYaX7xV4M8UNgF64gDza8Z6BIRE07r8gBtyYqxv4gGq+2
I77JB+LqaLtkyDmC7ivChRm6TaxDwO3PZz8Ss45vMD28pD7Uakh7NoBJDE+BhkjtDqug+xdIQr7u
QY/11vj5C8BKtgTCFU4B+hG4MvZ8gO+DNd8zcMaZG4jGlcdre4pvBLM3LFnnveWLHhN/zKCerXn6
HnsUK5gXWYwyLoYNRg4xNjSbz4IcUnUd+3FDvp2iZO7GE8M+s/6MKZiZGGir3DYbB1Nb9ZrPCe5V
jCzWjnvwE3dVAYmw6lJ+gfwsrnbSiZs1HRWttywP267q5lTzNjmv2OAtvwW5eOgxTEr8sxukSsDz
/sw1eVAD225Q8xJgOI5gPXbLg6EzdSR5PRHhgvQ8Q2TWJxrDpjjAj6cRJBzzcbaRWFE7Xx1LacxU
acuyVKeOWisc3MFzybTcg58qkUncrv6ueo0APPcKQEYptwcUW468rPJS+Prm55b9OY1Kxtr0f3P2
zOtxoCoul9AHpr9WeUNvKWOZZeyg6ktLQvinDLKUE8/trh7HR1Zh4s29AwlF3nB9QSbZ3NAHejkc
Wc39u9fedQxNVPGKyYZSTbZB0mj3ADR2glhSR8CMzDaWVJzYR5UQTR5b8n/gZGNo8iIH0K3QA7yC
A/Q7L66UlNIxKtQjadxzZGu2gvCHCnc0jY+iR3h9l18JSL+BnUKOMNIcAt1xtfLs164UXyiX3n4S
7lU5kiNA3RFisH+9N7w1sGIIJ6iVQkNZb/jfhPRlSfiFZUep6g0Zan/dQZTXcfGuSVXEcrOGjtPP
x2hOnDfrPeto3h1Ec8pth9AAbJFW6z1qY36SWVd+0J8PlzVn12fUOJ9g0D929Ndmd6NwWsNtx2LB
j2FKrFf14Z1Glb5MSrjMiYPcZGZGKVrIRhN1kP57bnrX/tXEOqsXLAlV7Ca6o6bFBwlNuoORW70l
GmFkw7h5GWnjjyTNc7D6LT8Wb4UDBk10b6eO3aL2Mt08X12/ChhWkzZjOjoRHKxP+97fkYqlqblv
KmV8trcvSwyLtX1hUIvmY1uwRZNxl8aaYX2IxnG8FGe98k0N5JW8a8MMqQ74M4jIr9opvTT/pXEe
UGAVjiv/y3hzBO4b1xA2CRoVsABkIhcmHGrBIX9sGoqe4BLixt8R+SggskTmuHdqqIgXVf5dqUlH
Xr+vBAneJUbPInb/wRq77CPrUamdlpef4igOldd6Q71ITmOevd2vB1K++z1BDgg4ChZCYyx5mTyw
5/0P6Ug7t81aBL2xDlM69E9BFB6Lz61AftmgvMHioWpqucaXstTJS1Y7Cfe5ASFLcWUEvVWHoH8W
JIFQnxWjt4fOw+zILijMHIqNA5Fk1YEJ56q4c49KvVWLNqkqgJrMuBKkhcC+GccY6fNALXB8UlrK
D8proGm3ybMpKh5hLNEpVIZvXjvyQ4hLTbR0NgdA+nbt4YkJohURhF6xTuJTQIUVmVVFa2Z0qB0B
5P1rUo6Ue3GZvNYXitozF9kywwG3Rwlj1/hMc3/wiOHyO+m2JaA1kKNtZUP32dTZEWOUL0y0G0mz
R7Ri2DhDa6uDZHWIhr0u8znBBU7SO+BkDUaw8Kvb+w3q7jRtOBvWq2qwDbjGIksg9E+L/MtpOBcj
L/PZg5XxNZZnBXa+QhhaPQQhG9XRU86FqKHwbP/5ihmCsDlhyIbzGUjRFQYC7tnPnUofoGytaTgU
lafeX2aRFs1HNl1lLXIaz8+h38MHTVgTOFDb5byKJXJfwJ3jelsmZCLnjFZLzzFFSHHIMhcxcASH
511nWbh3sU5h00KzfF0pAPnVqkHJn3R2KORmz9KZQnODOEnz3jRcd+6PF8pz2BSPxCGvqc4lT0bu
cd1JWMoZhUj4D0t6xNgBPDIz6tz5e+PstcPN+XqNtaElVVX6HKphusM47GL+0nS0pcleIRpYbUHM
jImGWLRctcwuYPPdFlmz2mPNthKff/rijG/GC9MQYIRuqE/RF3pcYS1dWKqFAVrHM1L3EAf3V6A2
j7Wk4K8Ypc6RgOLel4+Dfu45RESlL8tOwC6YK0AYn2r75zL3R/sebtnMYWzbk8r9M2dbMnDy+eLP
oUI5pf0BL3hEyU97nfVDB7eE3KYAzRv9CxsPnkXK/7fVf1dI6tFMb1xp2iM81bnARdB515HITsuj
pZBK+Pw6Tnr57n/3fxISC4N1YFSnD4rifI4lLYaY3euOepsmQbOz1eaTaHKOq48lWZr7foU76BkC
GszgKgn926ncEPbzv/MFp5WCvq4UU8VrlnzzeKvelUkX5viZiIuWa3Qbvbchyu+b/xpO8rdUj+fO
X76vdJnAKy6kMnirnj76JvUFiawWpWEmFXMM3VMjxWw5PTnTonn9NvIVwstqFNDITy6JG+v/HsLH
jtxnuttwjIckrpMl2dYOTTXDgiZoR4v23Dyy8oiWs0PATs0MiaZjqMeMDer7gxxiILi+8IP5JhId
XZRp544FTP8idsQ6QwBphvL9IpqotDfp8ZLKfr6F6qjXjDqO1ex1XkHeELFc2GUADcQGASfYhVvf
FAb8gsSOSyfUQ6sZU58yh/vrXz9R1j8TxgaMZ0v/UdI86FMU6rz+7YgaWKVqgy0C24rwdn+kUR/K
KlbbE3OeXz/WdEjQVUr+09cP06gBItuKD34AtJnyoDjOPtqP9QYUr52aDUXmMJmn+OffdSiT3Bxl
aIvuFwTUKTIL88FQjqxzKmpQ4vXJ2nW+Y5eFBOAqVrxeBRPUKe1ax7qqax3R89NkiwUDkhyqjHKL
VvjN/hJzb1nJj/xtH7cAq/pDbI5PghJkjc43G3DtLpvqLge9HEJ/0Vc6nQ+5nJs+b4SuDXFcqVga
rCjuL4F/ElBIZkAH+1TPK/LY6K17o+oW/TeuzUxGsi6mqpq80AnPrTP25ErTBBxKtRg1yd4PXYGD
Pfo/cEg7i1DfTOzs9l9a3/m++pgILQrJWkr1KDPWYS41YF286GqShr6kZclboy10j8lK6Vj1lYyQ
+1MSEKcAqTLGRtBFb8B9P3zgD3aquvkk9mOsyB7XN25wXnKPLPbioIZhi9VndtnEr43gniAj7ypt
zQp+dhbAW2gWGJTQ5PmxAuali1nObxV0b1BewGGqk6+cBgt6UpGEFPIC6d8TB52NOipevkA/QnZC
945iHzM1EacQ+ID+aXoyWvDfc0u1mgBrpLXPHBJct6tCV3sQ3otu/y9mzIKKvsKqSIAlIqnRz3Wn
pkIr+Lp27LHfzblX9R+bW4OywwphbzbKwbJEp4vsNDB0ujawHFUjz96ZG6vxOzd10dmBmRrPmKSW
wFVUKoz8+Dtt2cQX0PAMy0XrYCDt11vBrVOQac6dfSwDUo752sWzRJTN2frYREuKt1Tz41aNhT2n
6+m5Qs+FPtfEIKdPHZibt03P4V/qkavmSoSisCOvrDaGtY16gjLCRBk6r0KZrS/6a9jZIE0lTSce
yHyT1evWAB1iGkIsBpg+/+n5bwm7ntvVXbbKQFJPSTWqXtILyv0t4HBZ5+Vrx15NZKUcFoi0/NqV
cmlKPXFN98sB5+DjYcyjtRwwjZ/b1MLPvu0zDwYBK1Y/GiIhyZ8WjhyFdlFuHO5DO90YCgY3XI66
00wr8QAh5HzB5drXGPtXDCA+d0FAbDWhDzmSxXjpPvzQsg/hphT6fh26twnrlCGV7Rp6u9bP/a7n
Rtphgub+BFX1yIVupzRJNGn6dMGiGv5wI2s5PyWGgzAUeMk4HoV+w+/u8RSmYDa84kkQQ160XxQH
VZd5g+PhHLDGr/BCpKUMAHRtS6rE+3QUzXpdR8S/J9UZiHFFvc9UXuUeLVrUxqkfXpRPKZeLeiUQ
/+LpUScgX1uzwqLEHFMT9WPJs3q5eEsLH2fZPshGWtAOzJm6BeO9WWTtnYtzf8Y+5mlQ29N9lgd1
K4Vdpw5VnGXOqd7CU8Rjfb00o0P3TKTkLsHMznxQ0nTgRIxiuAA8d9rYUQoO8gjnK4D+rGSuZI67
bGagiOIuEnlsTun/D8kVYE+KYGsdbmZvagzpmD0n+H2u0ORdolIAWgrsreXNZYUzUxbSgoZPSUYI
L1kKD+SRSWC03RuBfQDOkCAWJjGg/xJms9TTrb4luc+5ea3SeWRDBPkUIbW6ERb6YQyR1JXjW/vt
pAfgTX59MmZgAY41ZizhbfSbCgEXgH1PdfbFTTQNDi3rNuzxAez07aaQYsrmPP95dJH98Qfty4Vg
m68cJ/kL21/zUolRRpU6TNhivunWcEQw/ljN3chjfFdog93Pm2WrJNHX/2NBkuW0FOeBBYU2OPCp
+K5pX1uDkuWYe4OH11Ius+qx9Rm/+y/Cdm++/X2eJtzDM3Ob+Hu1wosgU3hO17i2qfBB57mIWqOH
7vbhvt+ML95Oq4XKXsVU6+iYtqIpUW7QWMYaNxStr4Sw2KQCvG2yHxgcF//UFbSDdZ8I6BX52Q8b
NjCb1Vfz+w9XruKzkikpg4Vzn89p+zvX6t2tkWYWsTMX0ABnteoZHe4sAecj6XhrQ9ZRT9OjUbm+
nObArA1h6f8o83JivgANMKsjXKIQq3nMaUCJ7st+qaunQzXfgFQsy0+f2diLszhWrSBRTfKXuk9r
XFA4HLqNxcUw5IpktyFRgnHRLn+4hqVRTCAFv94/hef9+A4eWZoEbt5K5q9Rk+3w2J9zjoOZmBAH
iGLhBs4uZJNwrB0xs1KYgFye/j/Ive8oLouXnxB1PboyrmsXBclvMgx/PxlE5BW/K2+l4QrUAhds
CXvCcwAi78shW2DkaTZo5/J+9+L4QdNgTKLdCK2VNO5rH6MxhR75Q59El4drpV9MNrf+7k6delCI
AD2A1jq1An4ZO4D/SSNuZUoj+0ER7tYeXUHgzwREnUGC/yikdxygkUCfOa64S4g45zW28qGGjmXZ
cm0ep6GJ0IWATfowDndDwbw2W0GMwYmPxnKMMnM3ML9zApWNk66F/nOVH2twbeooOnJUPwwOcBq/
1trHTyW7avLL5qxmHkT3YkDe5FSn7qZ+yWdAM1407QOoY9YaB2mUYceCnWB0COWfpzehTKP+4aYu
Pm123s6rfvPcbfN/talbEXCrcbJRReaXi1gBjl71nZH2yqQqatZBLbuz5JY6GHq5poSat61mBTyS
885hV6nGS02IoRyzAg44xZ9h88gieytpA4/Ls2LSvkn5qj7XciaVjoxITVjK3Hn4+aszif2jFJei
PLfxUnf5hfkkdtFZHonvYNoPsryUfkPmD9zs03IB7NlI865KZpYDt5LJRTxxsT0/lXlLQLwY1QS6
qChAARJv3BzkQ0/lNbdByq2unAjV26/roUtY1M0VAd08vtju9YUBt0iqppQMQKoUAbnc6TyrNXYu
7E9OjuBsNBdODr3PuBCybGHZDfwuqIrSIkRmLo2bdX8/gNjIDwEgflrX7R/nA7OdB8KPvsFLdwy1
/1rGOmbArBX6CzZSbcONA12pLWYFqlazDl/Idvssplxka35qQDteNBYDV7rxEIOkfCznUANXO3EL
yi4JcE92CdNY6lncRT+cjYCPkpxnsaKBpXGOA8SZZpBDsp8EAL2ueXOG4BvsqT7gVbjflUovH19B
CQwUAreYA+xJlW/pA/vhovqWQ/0VujttGIltj5H7oQakse+ePrESb2rHQiaDDywmwKPBexMuDnCo
MebPprEPaW3GIgeAGy0nt2KQAvcGkRQ2mZDbrIjaoMewKwI8QTAOibdnCsATkZuyHfzcfX0z3cps
NzjH2NPjSLkAv8YfwlPZD42c0TT0W23AC66p1u0pGpqcdP8UfeMXvVH8oPuVCLqwQDwd/NClogyN
U9FWrrPu46Cmhhy5ESbvUTVWX+FysbdaKKGmhynzDQEdS5vQ0T5/dgIl/WJsgqbIXMjHmpOMwcF/
leKcZC1tbKOrsgjRSkiqEOHrVX+30IwVHcM6PBfXtZOn8zLwajmbmrj51l5rLzg7exqT/KWiJnC2
hMsoQmL6LrDddBVgV6DgpEAL0Jrg3esh63mgnbktgLVUEgGeLLyTXzJz5NXl36R8CHLVaE6z3P27
EnjcpGpifoaXk3OhwYNqaaqhibgrEZ4dTFDc/CTwprrolHfFlFokJ/3av7QTPdlmMSKx0G9snf4s
y7PdTsEE9ABgKxnJOi/JnmkUWXNfIuyxs3zeM7TM/lrX+e6kW9cdRO9OxJIBKtjUSvnyYcG9THEL
8xXUL874sh0OfxwxzhbtcWm+Me6ooWraOQ9RSPxzYwEItZN6DpicvEH9/IBjbeffp4FwtSXaKgvh
nVC8ce0E/hFy+FE+mBuEY8tA+Ej6vUkq8Xeew4lcceZJquauW3nNnVjqxec7hkSr6GsG8OgSQp3+
gUz/diQgVIXpJWM6ibRzMUbBKNCiu99WqChBvr3XOxRg8gNQJIJIDNMZYsxaPxnuXw6A74dPuO/A
+FBNizeNvlXnlU/znEa9Qoam6siML/qW2X6RBHPiuRbfQJAjYqo4wLfaUJWo9RX7roU6/AL1lMbZ
aF9V/yJF5QBe+cNbF0AR5vMe0s6K9FfSINc5Uej0cRp4HwgnL5UnmCytA66gcN9FbmR1tbhonp3c
iMSlUZBCwnpMfKI18aOGhitOktE0y2m9+9OH+/Jz7PkyaJU0387th/3RnZQ7+nQq/+zQBaL6rq0A
NDj/uee1WzolwXu20LHTJXH+51ve7pwzHSFItzNW+bUqgnSRMpx8sAVgwOJpLyKh0/hsaBisOLJL
AhAYNoSia6zpntLZ3WQywKLK2jrfKVsy4zYykAVfZ3JPafxBYpytS1XihgrR9hYfxtaTeuhNDe06
O16hUHvhHYouQCMrXwi7tJvyffB5nJWZKLCIWxbS12FIxU2HnWNAYab22CUJk/V30/9QQ8BTXjFs
OdERyUqbwxvSwfPagmYuT0Qr6g5iyi3M45eNL5x2canuMUIMR+O8fd9ZGISil2ARS1FBYPqczyX0
n79c0+wNRIFUmPbl1UAJI959cchynLTqrG9JFsGc//WNEPiMt1OH71MYJEnLUWsNv2Ms48rrhpLb
8XrsB5JcIu39QUQdZixtV6Klx29aZcUwOWzgN8EJVhQGch0C//XBKlUebqAaQmh6x6Nko58hWSvs
dxQkda3hW+AN4cVytWGfVuhMWaXn9W0/BMzypoa7x1pamOMuP1cn1vvYraur3PwVZ9MRakFzPC+0
khjyo43LeBhqK9ciaaQVItO1Yzbdp2svaLfe8Rjo1SB5GLgTqeQhD4kNiWlGPHRdwGUJxOf7p5X6
mHGVxhdWBBpCE5udGHPAi6/IshCNNTnw3VMkEUFB4x6gKKKmrQzjyeVvh1FriD4b15O8qvW/nKS2
zdjznBggWDXa3NjhdI0NNTGvSm880QmHEQu0Ennc7xncpSXKlLKyfwaJDL4HC8vr5TAuqCdfD0do
T5QNEPO3inJ0rYfqWpxi9suaAqv64/TfmSjzm5kXPuvK/nlq+RTJ7lLSv8tsRi8UA699hgYO36B4
QIx18XHkmhHAORsQEHqG0xGR5vzbRfKJz1YyujVFJowJAJfWsAtC591RZ9yS9l2uIKcjkOLKBBiH
FhjB+REX+uZ0/I9xG1FvTZVQ8Y3arymf71YydjDvf7RjypLADKMK232kaI0PPlgL+Oee8HzjBDCz
5m4Nm/gYz0GjPOLMq529jKFRtwH8fMEEkYRj266x/1QFtJXh37ayuFdpfGIII4E+JlIgb64oIlVS
GI4ie14sjB447RAXIh3JX0zJXq3wzzmY9YX40szPrtFSEN2lX/PiUtwxkHGjT1SbSXo6K50UmWG/
pnFuspaynNn5O3H4e+0/I2NEf7JW96D1s5fzh5fhLh78vrX7Rd82+Nvsa1vc2PYirty8h4U+Kq/l
BKE9QtA/w2TX+kmOSIC57nNOfLbEwlw+BhmVA2FdIRkWGeaO5pcaPyq8NvXVV0MlGnxwi7LjIutu
W42LgyMAR8qxf7/T+ofwJwct4Oxu88tMpJAXqi/tALUtGSzDQuFTCYkJmG1KVPxJz9b9ZqYfWwn4
7MaKvGWjCssnb5dmSkbvKVMb0wlz0Zix0GGF/qqILvuZ+MCXDAkLNnEkbjXOfR2cTfQgl+iEunSM
y9L1aFIauBPJtU2/2ewmbzOzlb2Ffd++fmtMy83Mslo9vjFldNihKoTSoJzDwZ3abHgZ35oaJJK8
/UGMXuLZmAr6X23DETlDR53Gy2uu8iGiGDMORYCAHsYAEBcFZ4pnp+X5T98RHT/56PF3xmWHdT2c
+0y6NzGgo92nc9ilWlv1eZeVH2ShjqsMLvJDO/7LzHl+koai7kbqOWJt2SeVYepFQ+V5ikAC9Yib
juYcMNANSTGtLGKzX5dTa3RbCz8YZzxvZdEu392D9uYmLjQWPeHCqD21EAVCwc6dzeV/3dfBU+5C
7HYdoM3TGJ08b3MdIjVrUt+3NpwG3LkXTToirESwMZDAF+t4HdMxXgpemsmZiKLp5eCPwjrVDLjV
BwlcEauuDrTHHop0uK0Vl1jSG52d0YR/Ml5nUUNuMgWi0pLbtN0TS/Yoc070ElBwwTaGi44GKwGR
fyps0jwqQHmI+NAtBzThI+BM11NPDvGOAmJj0a0t2thJeabypuQJ9YgBtR5SCVOEEHgoM50TsUh9
FUe7ZERtgi8X4B2i4RHwjZYWC8V9KxaZka61IGRxmY98Hg6N+zIUFoPY9x+add9Us/nSXJMK0VIa
JEKCctCEvz8U4Mw9y1FBRiKTLhYAx8DabEgtaaU6ODv+E5daMwyBG8zVcf1mR4kt+8rvxIbNLlMU
FgAsRz88j3dUQXU44RZTNOY/zudJBcoXckEITL2AhIsjI2kZvYBOS8v2Na4e+9A4T6I4AAxWxy72
C+60NyEs/hUsUAocdYjOiL8o7GCqtRRk7p1yqTzse8nx+2XH6MLe2mCm7Z2w8Llyvg40Y/D0q9tS
VeIc46i+JF5yq16t9QUhJ6yHYXYwDfkUmlzDrhvlJmwX8bt5UMF7ycVFdSeCfggDcI8dYq1mzgVO
zZcDHPMKGHS1gekRMFeoePZmIK1aAOAWt62qvvMMdazgf14QTC8w+cE65SCQqE+PQnvkL2Kua78s
hWHik07nmZWpaTOGJ1QbAuYOlwdWGKn1yAcqYhPwT8X9EfaMVDWa7GPNm51MyQEEfDD/vJ2YERi+
/GJ0h1utalSvZbiJE0nPe6WOVlXxSjW2QZ0LpA3HFf+cNluZOYHkewnB9a1fY4UlLzTJxZkOluDb
eyy6D7cRxcHMz3/gE4nlbsP4q3qshb5iKbFTAr5GzPfYJ/GwQ8hoij6VQjX4MZ23mNQ2jCv3bQdZ
txtWosxQK/O7HwYcw16c6Yb2l+uhWQqnbJQbQBK2EdkWyJYCwRrFydHmLujGgDJJ0zlffj5QV6Jo
DSqvn27NBqTQ7bnlaTZh5ADVHjwL9slhvW+ey5ym4jZeZdFbu4E1gTxSUHICAfnS2MSeA4tNj4nr
W8BBD0E3evbFKblLrC9sJ9eC95N4EdtHcPqRkMUoBJzIordXjqEB5z4YwM17z49RICFgSufSjuYg
lBJwLTkUW2Ydfpz5OYaqxxhTFGx10YaJZkv3DvJxgv8mR3gOjzU7m7XquH1oqsgIA5wgS3/a5ZjN
0bjzinVOBEgx29hy1QuhmfzMCSS9EmMDQeA95orImnVcJNqjf5P0GFLtNbSOiS/IUHGXw1dzwZcq
/sb8G+oCIrv1hkkKSM1QyL1ImxHovd1mYpUdCuK3x78wCYy5mNQe8POObCW6LkffXFcwynlCN1Dz
pvIOhSKyet1YCtH2F7dx18kVD+tY/RQCbg2VoFSn0vspL3FAFFPNFPXOeQzA8klSyLtmranas9Nk
+lbPnYa/1KSHEeiKosmWKpvXGO+hcQR6BZjXD9olmTCIMfMFx57qgbgQYK4TT3sa9enIxZJH5mvw
5nh369LSPU3nASslHhpznKtG1E2DBmhYyD+QG0NvQqz5GXvl2493VIBkxY/xGSHe1YasnqUt5Ilw
CAx0Bnegf/860FlFgqTjj1SAQCWiF5J9NxaQ5t9+vw8L/OE87cZCdoPQI6/joH46MqG7NCekM6yx
V2T2CBmgvNww4MqsGB54+hsHadFbS4F5QDL2IaqeKde6Dys6FZH/u3HhDYOeHhsHYuLwRYYP4WBX
Fk4MY3qeqmQKR7XGYkeaT/QSsMY9HdeezISkjyxNXas1FzTzs/cAua7LdZ0GKkbqhDwSlXz31AAg
nmq+H8sHmp2BH7BilX3Zkg6W45PQgS8GH8h/cau60TVGDT6xHjmfl4bca7sX/PEyKOQIbYZkXcqX
fEAaU3hKlxBa9lvNulh0JzV3uMYMQv3aiXZIxk94+8qW5NI9kER9x0T2FRAsbM5Sybzwcxx1dV3K
y4BFZscnXpZMmwjPk9PQVER4cSxQn4wFcgF6xXFXQa8dV4pBVE6rlxkGeuN0Wk62NQ+L0Pxfugp4
XM1A8df1Ioz6pnQlEGPUHOJP9xoI0Y3/ofGBuTJOmzX6l3xe1SpRKNthKyc8KCNlQksLxDzm6Ce2
OiVWyFSts96hXBHlBvBVxHG98WEgXy/O622t6hNaEoq1xTBBiVGMr7X+ejs74lIk0yTQctTWIiZz
OZxsfYdi12VMwYeXtBabWt5C9PI/9qmw25qKL1Or34i+1eiPP2/AUNquTPTPVBhjeipP3XsuFZ69
oX/SXSOcFpZM6eI68XNHFvfWLuVfv8J92trzJcz0YLteZHL7QWlp/u5WTvP+UGD7iJuQh7A0QcN8
JpGkEk8IQV7nnCAyhdQDtzxlSUGgxu8DNA1+i6oxgcPJEWlUqKnhzY3wE6VDqWnAUYsqXnQtMYuc
X9ZJ8xmNMmEqbazKQJvBLFQrEePkHbzz+sh+N7unSXbO5/hsCMOqmiM1a45ZXOUO0+Bf8N6IkjyQ
5FR8MYhkicAE2v7Pntiv6Rfzl6DFE9+LYqmwNxtRL/rxm/7jfAUiuRBrohvESG2FYzGOLT+3mVG1
5J1pqj6Z3IRXIj58DQ0ufQQKchG7TMfK5FIhFTBusNuk7f5F4ZPwBS0ER48PzP274RQdfkgsMXfk
E+UWRuHhPaAkIzbuASXwWh/Hxk1B+lKjZXgvD5+MAWgicPEW9tsO/YeeEvVPrLkr/iLGvJaqXKEj
iH6xBuMNBZMvF3NlQgDhfEA5EqoqBKtxzS3O8kn8dFmz5L9AQCZ1zCNu0mZA9GmVdgkQ6NIOcjPD
2EQc7h/jqejIVSwMOiMG4u8iCUPe5KrJfpsG46qJ9ewqZJe+Sh++KP+V1WiFh/U3uNL0wPa0y+Rt
anfLdt9edWrt2tI56BeE4f+HwNkCtWESZXc5tGDrSRGfMLi64dqeHjaFqbQt4PgdTOw8Zhx2UOZ3
wGGSDygaJk1bo7OU2lKE3ZRIdbOQGlWSemWI5ewNhVEjFVzPDJCbXhSZyJgKfOogg3/uLEy8rdkN
ayBNs9mxo4rFumFx4jeo3sFTLyCuOoQA1zN2C9ovr4XenthXTIAmxW6ehiOK5Cikvj6l5THZk7r6
i/9x2SbA0Nh5nGC4SFue7yMTyLo+TtNpBp4hh6l7nU35HH3XHnI0XA1jcIlQl8bon7ZObauie7kF
TEHRKzDlTxMJEm/lCYiZw6QD6tU84U/rjC5vq2fZXFLHWmoezGNM5A7eRbXCJNVUJHWXRB7HNlqa
e6I+NqdO67BlDlZmD77WqAi4VqO02vaMUecdX40dnqtbB2LM9VkeaoCYX+M1AhHxSPkHNc//C7ON
uB+UQYr/17lpKrNHbbIfo3VRpMJGoQpTA1UiOQmkQSTFYrKctBFNczsX5IKsxvxGa4qfhQmaET9o
szRD/R24x5viuZ4xF+eIOc7WILPl5L51vm+eGH5YbXWA6Rkie5mBb9/ZAjk5wjOiJdB/tTDn47sX
qKaUctePHjzjRsnvdyFOeFWe6qR4ZXTc1jKPxE2HS0YKDi3bb1XaLiKIoSFq9bSDDvG60GuCSPQb
hj7Ndhg0kC0jdwjNjkNNMJMQtyCncrcMChWxR9j0/OW8h8ODLXHemRmANIXx6Q0qFXzJi2RfBXXm
JCSCcICyB3whF+uHybTc5I8FdJ3XTM5AdvG5M6kh09siJ+gkus2vAI3DqF697Oq24MwM2xGvS6dP
zB3AxNPptEEomNJ8TbCxB1p7Qm+HMVuJQBCHROvuPUwVNKc7Ilk+zYBDqknjCgpjjw2hkXCf6eNx
+SLNtMaMZPgXpOHzWAd/JQH9C8Nf4nUU3vuOIKM18ImLkZlDNB5RpeMjTbUEKMKvzpKeiHT9Tdq2
DSwoMdpgrdeYf2dB0bVLsP1ap/u/lnyC9xRIEmyW49FT505TPeOWikFfyMu6bxBYQL+8md1NTTHX
jGSmIDseKuNLLAWkiprBAujgCGvYVhEnAFjVZcVNx6F+IB8eoFysLpDxW2zuQR7pqpjLWqy2unwj
yRJBzpX0NGgz70NOzt+gQ5Z6iyvsBSR3gJhsPo1KjfQjS4u6qT4q2e5Q8sWekcHxt7dC7x8m0A62
gnb7722NGbciLrqWiwfUxQGI2SLksa0ALew7rLVo+6jcW2S0m5Kd8rygCEZ4OeL3KTREkVGWLJ1d
RH9UOMIMO1BDQyA1JA2K9xWlJ/+XF7AIMaF9sDm8QyVc93HqpS0inP4jAhlfV43zzO9EGGeXvzQl
fmqz9BQ4EvC/a0+M2aUriXZ2ZothWN8k8wq31nIptQHSP0WtnouKW37zEdEQifcYiuoi+WByJbIn
bTl4f39jR7KSmH0KaHhTkQuf9ltjksYkWNGCJLr45GXPwdtXyzlvLMm0gnH9/EO/41FiNBkH5Woy
V3wfblqZcR1ZYwnuxlSgLANEq39w1AnyIcPiASkTTn79aOD/pDR66pUmTruaU/VIpHzbl/z97OZe
sebElCWLKWHb+IK9ZsKK3ey8q2vUShyJcp2U4SGNaP/nFztWxPIfPTB5EDeUicUKA3RH9lpYJpsV
YoyOaAwBVaCvvY+sAQRhJOKrgB8+/X6RN81Akg2EVoeg/23Fw1SN7ryQbj2cEtGXpMGCDiDX94JL
zcoQOluMNV8lK5fCMUtZwhhc/923tG1DtjB25cGauYOd6GZqz1JdVyTlRJoW7dfBnll0SMgpXyft
tYJyw3kmzRGZNr04VFSBIlE+7zFOVerEKsX4WedbZp7XtUmBPpjcNlV4tAPTRPUKZJPkX079PJiQ
t4Xmn5+M5eE1uKC7cVn9vyWI0+JtihOIY40Uot8kYI4fw1HoBjhuAlL2knauzMm+HXS9NEYMdGbg
CnaqoEWFZKN9IHoEcjXexmruk73ytA46mUsRFV6Lp+DLsB/RoZIKmvno5eGmUHaA5WUoRwlHR8jQ
Rwcfeb2E2DftlVoOqhjolYoNv7DaWLCxnqvlRCCDVJJCt2dBwNhopLS7WU2YhKkQjl2Mqh3fIkAv
/M8CDbweHuGOfJ2a0CDqR1nOkGrphbgDjgw+hrVoBQRT1Gh7oOd7QfBQp95B5jwU9lofejonOi1P
AZ01DyshnTy2mahp3VVuxnC0jN9kTNma4RmQCjLqEGCaDT378BpBTF0DQINPSU6dZEFBxejtSNKX
Ebc1BRi0fvmUtRMICdZto9Ot34DnGP0+BgoUbEh+2MWqmsR9Bp8j9P6P43QZGkCeEYE1aNAPr77l
kHcoD2k+ddyIEbCOdd9MguOalsKWBntB3yBlQ9/fl5/wcRLIAW80ztMSbOhdHq6Wz33gz3ex+ltY
JyslcfUtj8j0KDMG3JkGUQ25C0AXpXqCrzG1JTcrjbVq0OoAn1DuCegCdKj9YtQJkk5SxdiSYUFS
xbyBR06RSCeW8ocOShDX/7lZLqt6Ze9Sv4PZjfOVTV3zhu08S9A8sv4TkE2cR9Wfqs+wDYwvplZA
ohTE4j4u+iP4SJb/lhawJPbDDkPm8GkDZVR5YU3es1C+7ZqjJb1yuDKwUKT3vJ83gTNSy65q7mkJ
Djznunuf9G6+o8+FBnjCmO/GGHEuYenIC6+Cv00Hh3fCKMROM2FLWIAKRlHV4tZvASoRKwk1L0nI
+uBGPeUFqFX4gNJ2wFWY56+dODRd3wzSnXds0yklIEDBzhF8TykEkwzMbM0BjUN+At2Vzi/kEoKa
uXtLobpTVysW6+VUONSH1QWexAjC437WY29bTqLxgZ/6YuLpy5hDNs9Jo8w+pX8tsqfs2vUKNNvh
YAqLAtEcnl1ngfxjS6rsNTsWe39x5tGseUBAzt7ZB6CCkukUj84yRbBoRlC1I9K5+l/hhWq9SRy6
ULg3P6pAYJIgY6R+3Ky4Lsx+u0F5i47Xrnz2sussgYehPjd4tG1C3qp5zF4d2dirlOzJqv5cAOpJ
/gHTtkTmcitkW7h7eKE9uqNCFDSDlRoXu4r2iC4e94kDB+01ro/CQP2xKZQIkVAOg/SzXOjS0YIg
2V5sE0pkTAYExjDfJHRHQkOxYYzCamyn437YzWUxN0DPFS1bmm2tMLEoFogwjZq4H2bczP7/DQtr
ewtLcP0H4Y6X0xnlm1p793ejUB6A7eNtblosyB5exJivFKOZ0KU2QY6TFfdfohnnFB8+fTlcB+YV
iEy+u5t/SGXD+LrwuFILiRnt4WC00H14any1OF67qUtgrz1m3FtwHx5Sy5eDx+Nu7WKqWy0B6vaE
A4DFlDkv6LVfqEUp/SYvXoh1k/czQ86xcegkOVQiD6JmK6inPW/FPWisT/NNe8v555RvFeWzvZKl
9KMb8dlrFeoFmSW1UoEkXkcmH6aD7PRr8JqvSC03VSDo31e7hl2wTe2vgXrEaPzBV+rout63V+Ui
g2OPw2JjNmXTyW1NyieoxDOpLAFwAxnB35UuoBa72J70QOWkDFGeUzyUo02rrXyhPvvLLVmE1G4H
npQWyE5EDM1IAk7J1DXjQ28/j27iOcfItqPid4Z8/OYEQwB7olT9R3ePOSTm82+JBmtrymk7UrIe
CZItbmFSrPX9h1/TNwqnSHk/8vQys7yj+4ZbDmjQV2fOlKnzhPEzb9sbOJJMNfCSJ6sgoQiv9ivc
OxSq4FWoXj79ySJX/MKgSwC0K/GO2IRVCKLS9rxr7mnrFJPSc7UISJjymt96WhTs4Rod+DZHykwN
jBbxWn69HD55y4bugby/XJ8lTPqYGPMAgcb/yS17InH4KJ0Lk24iRKVF6ydVHjbLpunclm2qhe9k
39UYPXx8xZQMxLISj48/xjY3jqg8SLKWwGNvw6Dy8LrFI2qlsxWaNqev8pqFopx4pW3lkmeLtnFT
82PDXH7YfgShcLjia697c+2dh//oXQNP0tyiU8ZWJlcuwlzUa7lRGccpob3sYV8Y+rsaZ/T6yPnn
gdAIz2lO0ZemlqnKD379jmX4xharZyrD9jR7GiVqsfg3+8pt593difiya+47AigfeQR3kaqEz7DE
Z7ZBVwb8GKpSBp5RE8qfCnRjP7SyUz9PZh9pQkaIsVoJRO/sASU4BcvcpOs9UKu1h4v1iGUVpWm7
1SVg5FzxO0f4BV+4wXleM8ykNIZR89D5QLv9t/EHFIKVzzb8Qrp4gdo6ELwMLqNKHcvUrJnipgXZ
XHxaIPFWfEFz38xN9xDW5+weCjd0stRKR/SMFYFELrOClS9jTZhnxMuhL/LaW9X9LeKtwIFNr0Y5
k0F0KqnN8tf4eOCE78Pvju2S3wE/w+GHI4uLa+QIp+5uRANSFORUDX4g81dnRvnWq5kBds8bRkxH
XeO47gKp0eEPTTIafIt+X5FRpxG+/r2EuEjmMX3NwYnWBm3SS4DTU+jq93AcpP/qMYxl3agd/sZ4
HqiqB5pNU7zyppsGtR66MI7q/EmTkP0SUnAhIKMgJfXAmsXqS/LDEpo4Adz1Ppz2+daopnl8YaWH
kVHd/TMEz9Uk3s1JuhrDh52/Prq6SCIesOQqAdzF50OPIGqindCkwl0z/4ZxyMJENDn6CidKaSVO
1hF+f+9+o8mKqCC5uYSqY0GNxXqP03W+OQI5dS8K+az2eNJJzzWPtLJSPG5rwUdXWCXLhFVeXeLf
Iz9K1LL9e6KT8wN2ujpFk3IRJwyZRyL2qm8fKrd96IWmGcau/JA/ZhetJZSsX3YEqgcYpXSXLndx
R0lbepFqSD3iEl/rLRsUIf+y6tWVYP3/+h1qjk4v6pSeKUewaOYXIUUjyKGGs2tTCmZAnKwiLVbz
s/bfCBjgqtOAvdxPq9s0N0lHMZs9b/5L5O46nToX2n4f7+ADJ8gC6CC2i661pd0uhdlewMYPL4q7
T/lnMTLMtDdN3PuZh9gMWs0z20/bpu10YHvjnK05DKvPSsW9SO4DEwk+b9N52QcAL0Smgf1AsC5+
HFFeYI8RgoxWhOO2r/0/uQAzfG9j7n/XusmQ+ekJ1E2IsE2kWh3iHbooX3Pwe3rTv6Cux6OekggY
xqcPtRu1HvehEMM04XkAzakxnzKHEtDcIfFbFMXZRcrma/qx+LIcp4lmj04KswoP0ab/iX1zJDb/
OL89rvtxMx2ngjyVIPGAceiS3R2ZnimEbG1CfzvKLw402sVOyVl0Jaq4tacCReiNj6lXMgyz5d1V
VYhE+Bxey0HNadgXp3Km8Mm/lxoJP4UgTtpbPWZwomYg4F84VEMquCk7JOuUCZaUvAwetxsVz4Xt
SmbkWqm7l72lgVLkcJUnjBzLMEazw1mGUIY2i1pyhkknKKGNnttm50+t4pqIyI2jjrALY2yV84Pb
JsRXkfbKPLbr+mpCoYJpHKKFCyq3AllDuF5es4eiP+KpHMEwwPU4TAlCZOJMyLBM/cUArP2FeMyP
y0eNaN+q+VppPoyYUu0rerxt5i46dvHTa2FdAGRq01dzboG8pk0yedY10XeoVDvpnAvyUE/I0w6U
sikPvabXQJK81B6aOpsJ/4BwajC8074ah3ektU2HFiSbPARAbUq+yfghjRNns7zZObCSTUOwjKnz
IRgZhda/p9Wr2fy7xJuq+Pu0Oye42KidmIBbxEzIXRhjlLWt/7Lpm1f9vJQDtOsYMbN0GQW4Ox5r
d5OJqZY3xj6smRxNlAMMb4AxRVqzD0p1sdVW5g/rxLoMhqfFddWS/oM8A9F2ObE6kTXSakc6gyU8
Y2zIWW2YRITRqMMAVBi1COsjJBGc9juKwtMoPrzBjpGa/obqBZ55LcbLETzqjcvh6Yp4A6UCXVB5
Fo27m9hQiKMjFxbWBrEI+0itQT5ex3MIhV351djVyK/UTETjr1hc+NVujOXznq5ON7+t+svVFL85
adauhsSdpBfL6ubwB0x0rZAE03YBmcGSYCHw4ayVsTm2myKSWXM8CG9Gkw8UUYGatoSSYRCupFKR
xYylSsJ3hv3AAAsb1rUdfj9xdTPvycfxmq8zKqqMZQXTI+729VsgA2cnqMB9A+cDyp0DEHuHSD3Q
22+RQt6HdoPbHs+8WorDbM7I9dUZfqnk9RKs30lJ8qN0SqWo0zXTgRzfBkDzXAbKFhkw0+dg/ern
B5p9gss5/ovTovebimRjQUyTQWnWbM4sD9KcOfqItl3O8NbdzJ45hC8BCyPsNM6iWFC8QJwTctJV
yYDCTu0ncBRxgUDlHSC7IP7ztMcKxl/19slIVKwc3aRPTIruiKsOHiZ+5oR0UKEFzhotr1gIcjXU
fIikrVdkY6EQv0PzGxknh+wrO8/MKVIX0rwb21qX49WQfIRPSaCbsoX1pdK9VveDUopm7NArFF91
7Wh/hk164eqfh2tDT6Yd0D6Qqb73fmQRnTBDwMxBmp1uKGOaxbnFNnj/hijSy/uZu5SIkqvs2aOE
iBpUbFbLQ6mBDd5JdODOCMnDBoLxdRcUz6ob7OARw5AhyhH6JkBEXfmw9mlRVHbgM0PiW2poAsEm
xN1gpVaXY54edtpMG7VUMl6cXae/6UPJkjF6vjS0QCCSNMNJFlNN9p+Q1ruSxT8PInJAaGjahQC6
A99+Tvwfend//KYIadptU36b9H23YrPIPg/0PkpYNoPlxrcfnAWA9YnMrJ+ggTqkyir+HGEzax2r
9GMVsOEGyvOoC/cWQUqi4KjGIAIIbstega35uyMwvARWiIPZSuXVMhnoqLLgUN/bBgHeJtWeo5dv
J+khzaLzdREQoms2Hbrxz6FYWJBfKb3MXP9o9u+1qB6bHcYj8/u1BblHx6oQcWdSQkP9DGk8OBIf
knurl0ICfDwSKDReJzUc08JWzXPkZ4ujM9wa32n5ZyVlCcnS0BIbitTfk24gAc1s27IgCHSVIisy
b43wxNeDKkREAJ+3zS7Dx4u4tlzTz1sooq1KzsW+kBADGYMOwDSaCORKZNZFdL+hWL2igTBZJWHM
pAhh3SqZrZbZ6UIIpWqJj7j8V73dQy+6j8gnomj3OSIPU5qOSAS1Jt1VCYEw6fWkiSD8u1oMF3Zs
a4H7Mb/FMbPlyBJafdhXltS3ycToooajxYbSkgSHf59vQj2FLQmMQITS/PbtfEMwb6jGTuutKfdy
v5FQ/L6MAc4nAbaVs9ObZxHQ+9OQhH6On4mSB4zYpy5s2HNK0Ku3Np2JEilxCxb5Mk9Uc7s4eqnI
OE30ARLNnzeYnYSwDYs76/lYIYFDJqVsDP0K5GuUYLgC1LcBoRht9gN6sPfQ4c42Fo4UxxYxd6Ku
qGochdyrtfy4hmhcWXwp+E+v1/eN2Y753ijYCXPBp4Ba8+YeDug+MfoSabq1dhG3jO33l0cLPOUZ
xaTn72M2lTqn03Qvk4NTTUQg3e8NhGGrHga4i5bgL++p1DJ/qEllHdmzCXy5dy7sAVr22XyUsNGF
cCnZgzYFvWV4bypcyhDwcGzi5qy1zHDFMRLYe63jkTJ4jr1rL3XFrqTqbnkxlM58cYdMjPm0bnXG
ItV1sfMljsev6FprPsKiNERVpnob8X39+NM1hHnov3dzExa5odwEm8TE1mVEhJZVj7FmlZu3UpLI
kjfmx78OLiYDjK0RJp9HMx65pdwibd0QcP077LicxL5pPTlkwSj7h5Ii6uVzJk11zeaMK38kW7c6
p/xyieroO9kxEGwiZYdsCbcwQ4lUdK2eInjl5uBCMxrsNCRHXe0hbzr9j3+0kZO4RDGDlExigahN
o064195CQmq/zilZI2NETW60vg9FGwsIrQOGRnOwkiHto2M4uhmXlspm5RiPl0XwKOtpezcjk07W
eMcXHO5xCvLCLad3WbJZ+6vEjO7xHbQLHZq7BP7/Y2LmhoS8SyjbfuqodenqwMogyAw/6SnNWK6v
ns7qwHIW3eoHb2GcsObc+Wny3SGilDhuf/gujRHa4J/uaeTShnQS1J2mCXfmamKbSWfas7sPgkr4
e+IVXRkUVqV9zG4A6arN/8KKdYsSXrkAyJEoGb2Ml4Q1Z/X+sQRLlc7mXZ1NHtAZUVgVQvFs3WmI
LKzk1f3VCsDNqzMdnQlZIEgKWPQaCxejYXaKmRny6v14bDG+5FA4pR5Ji5nB4+eqe+tFv8/s/JeL
91gP5JqbBefsr6UFPFcVNxHGxuWwJ44+ockMTm39IW8zo1oN9y4LfFKdnRvtDgJxt8aVfpjZTGZ6
uzMtEOUae7Kw6pHk4rGq+T/jH7SaAfkkhkVX6uWJthHP9C263nRQaPcwKSqFmTRtncSHDFV5234K
+GouHA7irP6dwfNqoIeAYiI+e5Wg+RNWtv+UTnhTckczfhPPS/84gA5c+gyTfBw8nCLqEHUB3CGc
Ej4l+G9Ny8zeT9HUWQkMCiHduBgNQ6ZNLo/k18rkc2QaiGl3CLYEEIV2b76lvYDG/f5SaKvoAdzT
zYgA6+SjHN7oxLC0TYFYgZ2bpQFTx3y7Dc/gPU2C6PH0vp4sOPieWmwoV4JO/IWyprxCAwzNWGU9
6G+Bx89M8Y6i4/v2r7tZa0P5B5DqlJeBGHTFuY/HhHkenpex6piAMX8am7P5eXxQJ8MmOCQBfErD
O/4OAQErEVXyfTBYRhIzTp93RPDIRnikDv9f7CaWzxFlrPKcYF+xYK5emX34vsiHy/OOft/OVFzl
kvR4sWZhshuI+SS/g+CBqpNLOADX+nyK1Ra5pVoAxR0UmxpLW1fbCLodI2qgtEbG8eYNT8JGwooq
2HgtIItpaEwWwz01pQIpahCqq2mSEwoy7+43QNhQ3uN8mVpmbvZOOO5AFcLb7Ouo14B0V2PkM88F
9oV5pMCkDeiaLm9N4HiETjpqiXZwZ20B96bTS+3+M4WoEAoKRbnsdu9EDC6I+d09e3GMJG8sBwNB
TMptaCzcTMbMtoR0bkBnspiO/7ydHhOQq02Fn05HampFLVVXH3D/FkmeSLzs67yBtdnoX4Y6ShlZ
tP0VYQn/kb/GXlsDQByOSD+5hJuqWplER1LorcfdHiMZtMIYqqa2BOsJ+iCEmDq/S0WiMyihDenQ
8GoQpZHdkqpN/qgDscBaFr2gq0cKSPBCtrBeXMqygAb1jU1jHMX5gJW+qSbPXKEVLNOeK70Zhb+W
UZaKgzQONa5GcR6SY2zIX0MDTUYrO9KWsJNuKxAEygpTJV767o1OAg7fKKCcKpd0FWN9gqygqe9I
Yi0VUuAf5f+EdI8HnxXjyHKtiE2Goy+/mJXMzpxGQ1NrfMeI5nNweUeJyHf+MeDoYMM8ktmE6FGr
3oVZzIBj4zV39YA7o/9Teb/laXcqztpfJpwe/N372xeZ+pyOU4dPRrUqQD+jQd4uNnmrrh3/4Hlf
zNgGec6+rzoQ1Z9TUA9YBsllRRLP1s8PU7PL4SOpjCgG64+ckbc5tDWfpQAetWYsmkejN7WfYRKl
Sxh0Fign2rPjZxVWUfoVv4HX2XmoFBv7vVGfc04zvbqwDJM379o+Ef/PHaPnqgpnV+QnIBsKrWPD
emcFZwWo4okjiABf1NgAeBJ5Jghclj/SYWGFbOo+ZAM6AHcr5xRurNPeFGThJBm/P8xB4lPrFQOH
TIGMrFWaXH/+69l3y4iykoVkmZ5x2TtkFy1Z/594XWr2G4b3rR1y4z4U/V8jv28+bRjFnE+b6AoZ
Q4JKIToRseiz7T9yB9e3noulnQh9aXJQyTuabi5b3hVFc7+DnuJO2X/kuPq92Z5kKT8cSFNnhwkY
FcNxGcIsvc3VuFX8H/rStbZaUZM1+FHv0XzEH472ib2FaKImPqizc0pUvcve9DhqiBbK/+kAjqgp
jv1laAjS5z5Au+8GErajh0X7ok2S3aWI6p/sUKXV4DHgXFNtcriHy69Jo2pVwYtz5WYcg2m+71cH
lLdLL+F6XcjAPPAZoSwRKpCK8UEgBaX79p+OXBXGsnMocZ8bauukgt/r1ZJaQ6QrsbHmQJJ6OjkL
v4yPXNdLF5qeNsAU+b2AoLXcEv6O4LG1opRI6uyG69cN+rkrJm6PadKV4QlfdONYT3SfF2GRf0OS
7QBo3rA6/H3EVqqueu0tqxN/MXtl6SBDhTInSt6tJoEnvvxpjqj5IWdXusv5VldgtTxTLNU7biT5
wD+Ogx25KN//DFbxlCpIWCkxe+FFrB7cVryE9iVtq/vz6j7vBi5xFpeBAyJ+Xuk+us4Sca0d8XE5
BDfmy4HRCO82RGkSJwVAZyItOBDIH0P4DcY/at1Q4UvFW2hqrWP+bEs3dx67mwzDjut2vtgUtz5F
BFvpOa7gsDjwn916yATjxZ48sTHDSnSbCpQy+8IN939wyBV1+z24uHf4fR8jeeWD0WvZLasQQic5
9a58wKNyNQCBy22a3oMk09V05y48LLuXYSkE09GuJ/447oBwTShqRMIfuxrjHKWX4r1Tnkyjaa1n
ELYdH14SZsgVQPF1ZybcoT5u3YmO9ZtILFsRHevnbbe/bxlOizQV2hrzyothG/9V5U1wkrUyeIPh
S6QyxCUE2GuhQ9WhLBv46lBllgW6PHBY5+U1svM7+lPNfNiiiuALdwn2OBUTrABqObfa1p+kNygQ
U6q5HCDJgApJC1xXR2tui+Jgjh6FbbF9ZIw8NqD/0YvcKZJdilJU9Cc8XcAKJ0X7TrNpbuDLvsgq
s+Y1iB2HvFtcGqaopZPzvaAhWni7tNDZ0WBGY9U1wQydM76CaYaMDlJI556cF2TfJv1jVYrajrW/
H5qDfnC3qfmHWhJbTMu+Bm5yxrl/gwuUJ4LnU+c68VQTYgmCgGqVnv47kihb20Zk2zS0Hro8Fnlm
FibK9Dsu/A6a6EiMRo+A6jF3iR+jeCem+3UOCeUeSRN3XaUKT/upAuLQPDLMsvK8EAPKY5k5oEk1
iMKbQNL6M51/0l1RrY3L6iVI2Vuyuhz/Eg2kO2eAV1E6jS0gPQyVDTLpwwWTzC8Yfl2taJ+oW3lJ
eigz42ug4CFrDwwi5WOTAxsCv7ehm2CxrgfwN0kBUawWK/O9dXY33UxOQkjeLPATjZX5thdNiJSS
ke7b9DbwPNKXB5+9WxYYUfQX90j5BTs9+viJWgPGUHXB9ZAESovgr89F8tSojPfhn8KZRW0LEnS8
lbhP9udTt6etBVoZhs8cHo/kg4CXUGwt+lZfAJCKKaKtHlR+bsF3LlL+pZ27te1JtnJKaGDxFSt+
0Dfb2LXegoKLr3Xa9PPW7UjtPJkihPTuBcvBi+E76t018RM5WWD7mJdoG4zWSzDa7sukHpYGJ53q
LJPWV15z1KwPonCigxxZdp5m4VgwWHrUeBzhHs03MZ+KdRWrPZd3ca1P5mE1EwsoEuF1S++b0MCR
nnAkwxFrqBdJcyBICIDv5GM1yLdM1aHvRSWc97JkVQuqa/Z2ejiV4NdBbUK0IQdupe+6+KojRP5J
sZ+4ifNkB2W5d085XAn/UKjhuUGf1TbkeSZskJbo7HnC3mUpDb5hxL4bxGY+MbVEg4oP4MWBxKSu
kmf7Uhj+jKMY4HM7ykWt9VMzvtXTJTFmu2s9fODHtKqCjMNkjodGRySZkX8jYNX3W1/3Db5GI8BB
sRSAmm8/AxW2gaFh2LU+wBf0OhPjF4TqnOCUGN9mDyE9VdKJJqQ7Jc/ixQXhhdzlE0H6UKaKFjIY
EWETe9uZf1QUs0cYFEHez/TpNxghbabGn9nCHkfz+emfBZz9yk898a7wnJG/FAS0Tqu6ankYwGpx
5c/4kS3yDediol0NLx/C02FILeQgcZCNifNairoNItiZ6Zr8e7BQ7bbe1FK3d8wtHAQ80jSJSqCX
2N9F9Fr/vpUvwz3RuoNZLTp9qSHylq5Znceha9lERzhxKAtWJ0YA+DS7Ieto22KQ4r3omUllIO/T
kMqhjVnNb4/4RFjRRDsXog+C4v2eFklGKhR6f3AxkXF2hG4OEGXS1sZeyodMUSlHm4rRaNdSOGYN
rYmqo9ifUJXMTrIdHYOJO/T5YkLkCg8yiuXp4UAJyg4LbOo7ioaknka7vcIolgoDq/Mgg02kvTGu
Jv9/ZEwfGI2H6JtsATp1Ugh2RSn3FTPmK/BAgVukPYn1kFnWP7gU41TBG6i+nB6zL6n7PF0JJs86
muMmTvEGp9s10IL660Ce66HOzAce+3Y+oRKEvpTVwPmejQpyQ7/WlYC+iG0DSH3FLsVUmAhu1SpN
FESFGztJVXBTt12oOR/VUxzqQOsOC4xzF8WrSKWb+nU/7tVYplQ+F4ewGocAXv4pWa/yJhWf3clR
ulM/fKe4oObG1Ta3LTGnWawC1n+SZfXysJMOI4Yt/ut2mAWBHDp//hWQ+0lrSqgJxkrXrwGFwTCS
sYM4/9N7mXnzMO0kgMCCiojzNMxwjsgKEAL1Zzc1YwDzrfU2S8/lO1beJE92EV42aFjJ1CiKELJ2
XL7alftjgNntbDQPYxug9pF4QcbFmm2Gpke1fqXK1Rhw+bEE8XroDYNdPGRSCCz6XubH/HZjeuOF
ICDY7qgDM2QWxhUYujjfDe5E/sX/d9ah3+vLv2U2WXi1EAJwzR9aPcgV68RmRzyH0lhhft9ukJCe
73JO836yskRO+HMWSmKda5ToJX87epoxKwjPAZ13LBdrTklt8T8D9PIlSzLrlqqIGooWXZ0b/9OJ
UMUG1gh8cLav6nVZsg5Sg1g/ry88iFM7LaQ1+CRxas9J000+cwJmU45cJ1kQAlxYAofg2WB9mz1W
qrW8df7VmWREZs9rUMNPRB30usg4jq43PbYtkN627c5Las2yXOJJcgEACsAIn0J3eM8navij+G0J
1n59nwHoVldTMOkQvptyqbtB6hfW0hUHOaBj/mw7KQlUYcu4nkEoM5vtU4NAzL0QmtvHGO5rxaQC
3rX89E3SK06zgQMqwWJDJbuaqmyxTYZpmfvkIj9vKtr69mnSbRsZI8wq3RPxlLjQpf+6Vskx15kn
k2SYp0WbNCzNifZzKpuvT+X7qa3/55UKII5eY+9zLITTvARiUXO3o4GtOdq0hzJ1FvJFkg8Uu+Ga
TsYteZcdMt5LW9JMa/NbKmRaVxW1qag4/kXmkD9pV6y9saa/blSctCa9OseHP0yAmyBlZgKiyLax
lhl/tJR0M+8G8tRyrdwZApr6qBqcmZJI1UHDg2f7avao89/ktRQ3Q49OCbRm5vCwH65ikrD5M96j
E5PVxfTVLlryyd64qx8Cq1fjut9/Z39HcSVD3K7agVGgMoVgVgVhtlu+XF0jmYrY4bv/0BvZ01OM
pq5ze3bTvrq6Z9r1bunWhQHVOar9STH8YrLnE8jEZN5V9b9VWMoxJmjb9W7DEEcvyolJWe/3MejL
cfI5g1nJd8/19UbXjM2mB7mgF12c5skf7oaZ3569shCJBpclYynaiOYJjgeRpcdEjxH9QLPUdyjp
8tmi+YXaXD8wns9LSl8mt3QGsjbyST0DnxyaW/5OyIWyy11c+3F0pz7Myb9ABLzYVFPoLmTZJdFr
cVfdiueBN/kAqw87VCbETtiRG3poJt/bBOGRJxKU+cPn6mkRjdXeMTeXI19Rmmbat3wJQPAmjm4E
S4nSbS/V1Rf7zqZ92mKpgL7yBJaUA2BYRadhyWYKyC5BSJmLtCKkdoJKFRbHfdpo3/FMn/YdvHM1
Kylf0jKqkW+1GPS/MgzKVFxzLJRMxVAg+NHtehlTE0DAPPZnaWPCzlbfXGyPfkvXdVbKEv965gKT
NJq+odm1hSN/+CjTvzXOK2mCfzimd7g6JzK5DUZ5hxzsSw5WSnSGBnEzHljIPaNw3ypD9f3zGHL7
gYVEACMSNP3wjcf94i7hu2ex+omauVdqOA3huGWEJSiZf3VQQ6l9aWdQ4yKbaarq/tM+m7dpXmn6
JBGvklf6fKgKz/ZbefZPjROyR5k23DU8e9yAfQCJYDV4gkeAULxs68W52i3wLmDW4eJu1noJ9kSN
T/RJ/SdK0f8pDhB/TaMp/F0NOPCVJHtfKd7Ma3lEUe6XcTm6lEluohKbTlERx7bICjn1xDFZxf0U
aJcyZZWgAtyejeWTuYFgeKgGtspRCSo0rzOMObbbX9uWrvzWveeIOaPqroh3/FJ/7SoYkzQ7Nm1d
IM9FWfINO7O00pTaMYGaI4kjPoGBT+o222LiQo/uvFi9X5ukr5uX0O+UbshjhLu1SaTeIN5f8fFe
R1ASkLv5lTw/g9AlKG/9XcjWOedqBxVez7vs0TmyDY/h5GpYGuoSlK1jimidmRK0vjBOeQ0ZkiiO
EV5vDX7yhz1kdcGNzCv0WeiM78Mi4t9e0tdBSS8UaDqjgsW/kijP7mtkkBWhfjqVesbPdT1jSjaj
BvyEq6CgE5Iz8bqaBsX7/aSfvW5nADcRoHL/a6NBkPJVUlyx3qLhYQhLaBMhqZ4LIUvk8ANAElA+
vPtyKW2FzBg1dJTIsbeBFuHaIGlIN9m6STG1mn2QjDWywMZ0dXwohowYV12PvGd/gs56JsL//jXA
+iTx8ynugUzUpKggSmZi+kK9OW1lINqblnXNTQ5URkY7If0kcPwcXFd0RNzuUO8fdDqqHdvTaAh8
oOK99SmQfQIWvN7JO9dKip3gJ9aKSVbUkf0g14InsspfXZ33qt+51BO+z8ulY19VQdW8P0NfqB19
japGZUdM03oXWiEuKPH24Pj90i9YQy2Ge5wD8CTX4SahxyZwDeF5+/7yuDisG8Ikf4bBcHIcrRUQ
Dfu/a6Su9//ZLkYO06hQ8eUpZhScvn2Vqoxb2Pup+OK+q7tvmXQN9c+YG9Q2wOyLzJGwgmR4EUhq
eVDjIK2ea7SVigr87Yqa7xDJxk8VMM23IOD03pH5FmOblNJyHK73JBHhuAKGjWoP+CBd35z8j8y7
/O+qrW5/0dt+cerRpNYr/ScsFnI0So3RaelgSFqVoWkXPJm2aEZ0OkGZSPFV2XVM0dzrhf3wfHk0
AR+x8Ym0uFZTMhKwQWb1dC0zQzW9Z6QjKhTmhKNCzTvdqfDqfN1Ocl0J2PRn657r7Ha1jFlqqnBL
RA3/wV0RXzjY/6XzEzDOSHG8Vkv0/gyOcTVAjD5sTpwMTU5k/mGMTr5JqGRvhrhtQnWgwh5ZtITg
XeJ2yzJrzxkwC75Vr1ISzP/6fJh9fGHtplQzqL5oJOfwjUBI8Dqgw1oipdHW0xQwW0OGIth8c0zi
qXvFWLYfYNUdFLs0dSKAiuVQDcKmNzfh1B0bP5DUd9v1ACLCyt/Qkazuo/v/zTf3TK0nWbsbq2R/
1J56L0k/Z5fbUzCpACpmulU/XDXwLSKLDfZKNCkI9ca2NlyI8f8LaC6PB1relBYubQbMMgYb8RBb
o4IswMXzXhUEXhZH0PbbPcREgFv0QgJbL4cj/iJt89CAv9a7duBXPkR4up+L8unmdhgwzEqDXend
1kglgvKO6i9zyvR57MGhP3cH4GOUEQiOzxugmb493P4QijAckNlJrxBG7TFZWPTkztXUr/jG9Zzb
cZ3slc6Ag+S4ypYL7oYVVpfm7L+xhCdE8go1c2LD1+69g1ADaL++9hMmPyTw8gfymjvFd/+2hRqO
BDhQagYFWljl+RK7KeHfVEMHjNwaJF8LdSjt3t7HlFrnJIx2UFprjHDxhPkyXlVdwLQVxmrTZS/U
0oq4xH9NCDeHSSDAIx2Re5jJ0JLEJH1zfFsczzTWWHB48KV/qNn+wHRf2tdA2DT6LiLKBwEl0XcQ
sT8U9EG5ri4znFNTc71OBXT5ubaqzD1bE2QqMs4C+D5jM61NpkCpMNtCdpy/ZbDgWNkLp6jWXcui
KByJqAPH25qJUlnQ43l5xLVN/3Inlip14x9lN1U3t+WSN/fP0V8QpOtjFj1FV1vpLZRs7fA9VKAy
UqTq2Zl5uTqvi5kSuOdm29vLtgLfkNDFcw70fIcM6mNdV2WvS6dSod0jocPPJFtcqCKY0u1HJsw9
s2rVowD5wzPjTZ60dS0qu3Iq7gVXRRZmjSxR0sk3rqxJpaO+bKads2I5VUqSMyrXMJvB7Ea0JsAY
EDVFMGQMhMuidOtaafKv+tfwENV8dV9r06Wbat0vFt9l4FxcuCS2tpLvoKiBNOufw7qG3AoEw6y7
+6UgH6MLyjjTnQ0v4WT8ch5zAgLcctu9uBY0alrKxEBiIGRc2zpV9IhW2lDc4//TP8RZLSXA35bY
FOJivRTydRcQcc3bmSThTTxJe+c1UHau9p11oGOm8vpPD1YrPnPovfcCroyS5Z3/npfZm8IGOPEM
PLB4JIkgfZ7SFbTGJCuCq92QRpYbOtfqyRV4/HleVhCOGOPwtLv90070Qsb8SopBWfoiMnwjyHkO
txVGZaFEUkh1wLziMzCp2D1O6No7vRzI2xj551PhWY8bdg7G9IYVsVcDEfsAGsJRAZ6NtyYh8Qra
2lFALHgikQ5c13BL0BXSrjLEIpAQMjSaicg73rbLaSGd2ZWOID/kElZboBe/uek/3rxbY2NaNz+F
Sdo0lSTruWkmlpoqbn4SMKmFZsc9baw44tJ7zwRh2JC006B0SNMcMiZAv1SJRaIEoWeUlMCvcvbv
gMklpz1TtrsFER+Y4eEBWC76aEdBHlsMsq9jwP9lbmBaHj7QhwIQYOx7eEW5zzmtlbL0sdvvvxk2
ZJyGR0iUmgqAAOsPASG7//zFHw9WXD2Mws3T2KAhffknDhdGLbxYr2ke96EdKLnN/EYsapy53hRs
xXnRh/e/vR4PZ9v+WG5ip4JWFredEqYEn+XD+hk1eDk3p9EBeRdF8lPUymikH8qeL1dwExGDav9o
1pWJO4Z98W95Eb3iaIQVYvTQiqT6J0gCiLDaXAPXofP6t7A6Z6gQpDcg30FvVLVtApFLQ4ZUGwg2
q4Zqp9gmFrqvQDJSnlMZ9YlPJ2sKKWhzPNWGv9RAV1aLeg/d93CKHAEPaKVhAlYcfFtyzKtHgXlO
bi+wsgEDMiEQ64qL/2I/aTT8j3j9j4kmwC0rmdYiddDTgMDVFd+WufhLflGO65K9+j1jnCjTgg45
RdHwWqog7iWvxM0uC46ZEhAkfmHaI/+Si7Up3GaaiB3WLEYP5Tw7cV5wGdRt9PavZCNuYlZddmzL
EJwiKHr45sAC2Bv/7jxrLeFWbujqH314FyH6/M+vsVHamSrRPM+ScZBmkXTG5NEc8HmmA9g4HLd6
KzdyVJifvmtRitvO5/Mr7QUTL6vRjpz0YMgSUDvcqMYnCquUj0LAqq5qIJs6EXmXRWn/7J0LRAZ1
KWT179Pb/l6Qn/AZMWEaB4OYWYJrkMnlnnu+mcCqN8wCMhysUIbPOzJJFTbNHrte209Pbj4Klluy
+ldk5mbrpckaYAWbItV4TPuFwA/Pr9skOTNlnugse86Aq+rLgnyuyv8GaxiyGxrJhm/7o/zTcEbs
VI/c4QrK5DklwvLmtmTZmEV/IACHO4bcmpOCT5onaTSl5xn5txKeIvrNcxj/Hr2yrXgj5mdp1kK7
VJ01sg3U/Jwpkgfx6QF1DaLGvX88l9vV40ng1TgWyxhFH0i/kJpxn+ZasbhFY5fewW+iAE3h1N0b
G3ZlxkIxoMkXTRDYC/ztNA0DSBifX4iJe0PmHjo6BrGNYkiWpGj43PQssPYuoSuobHWYXgW/eRqC
h6z+SnRkMTcwflJTuQMepAMtx2uZEewXVtW5ITAUdCp/hD3Vn2M8uUrO47H+IXhrs9AXM60XMe/0
f1MtQSsCt9C3DdgVzKGiAw+T9yKy99myc0qqHUsQXn2VGvELIn/99usU+C8Acj+xxW7GccZ4Qt2g
P4abW5VQFamwy85i8vS9xzjPjwtKTGWefXlmOby9dIL1VwaQbwh0GGQ/QbWp7d/6epwARMOViTBR
/OrMSOUD6PYqqEpkKQJkSMjBdWrXq6qfmrOvW5n9QuqXVslFwgSUfM4ke6xLpTR52pY36buAn43q
XAIm/H0tbDDnVeoYFQzD5cgDm6MuU961HXgfj+TDpl4EcGqSgTUrB4UZqS4R5OGiSCBHwqVclDG3
yW3uP+8W65aOQ0Tym6JqThBaHViiYV9Nf/KePlXUSpPz5dTvEXLQNQRe+1GH6fHbGrmkSpN8Itb5
NlP1fB2DoeGP/rhurLTm18bHXLzdQDaAJ7/XW2lvv2OyvK1S3MzH4eHCeZJuVmQ6GWVDV5tL3kpe
5C2vu5InGgxTQSvBjrdaUsFweVd7FfcfsS4WxR5t/B4tdQGV1FJPSm6P5UrSGqmN8TQFEi8GRT9u
FYOwzbGkFOHeuhHiYUbfIJNJY0GO/c0H3vvrZX/3wfRFpsjEiTr0Gi9mU1PdR8nx7BkaWeiaYAVN
I5V2tPaoODevZ71VExH9pF3+KEIQebFSpCjKbYcbVSoylvb1GrX5EWYTvT/hCkhA2zTlUuujnQ5K
+aGfW6Ye0tcpJZZaOhZlA+3PoUQm1VhvkVYR6BihsUY0NOsR5Nlx3U3I2Qb95NKm58DGMQ56gOvR
UU3LpEJVhXxLVdCRqqKxXfjJ9woG5qkCMazPAprN3nfMUIJOMH4qc7gVg81kGbEaHQtcP0HzWhNg
Kgl26gz7c1PsEdc35TiVP7ZRHgl8vTrpGtz9hQ17RRTsuCN1a5Pc+oR074ffsUkVxr4MibboirUu
TAde9Pcb4SuUQf8aDjGTcn5EkE9alKZMr1IAMjmBwbL/IcwWYYEJRHVrMTDSefRjRg4kPX/CYDnH
vGyZA7GlZgCrPZWH797BeC+gQl3XEz7AvGL2TFe0+S7DQk5alYsfGoJ5PPgrv/yBY2hBXm2ZjDuS
01o41a712DizM3dy6B8TSxw+6wWIPHzAxRC4TuIgjdP95oqiyh2/U9cvZyyaLjzDzpT4YThUkgXt
ig7R5hq5IMVsVgSyBWmnfgohrI5eF+V5nUuynUsZOh/3jspAthGqghXJq27+Vf1/aE4vgaklLc83
i/A7gw2GWPoZ2worBm4jymNcSPzRS1ySAs3Yw3dlMdFGwJE53izJML4bBw0o3SkMsUA1QfTVDsEU
QS3aZz2vTmr9+riMhCVelE6+9s+mOX4AdQbo7V3mhNfDZWOuQNVA9eESvAY3nes1+0uA1VFzvbN4
OmENtMP4T9K3/QRwfUNHTR/g/ktbq38m5LFLTmf5CveshNGQH4PgKCEMZfbDlE/9Bic14209bxaI
m4a1VGzNZKRi2M/dv7xoY/80/YuJzYZdRcflN6HWEc07pj6JS3/MJIU36bVd1k32VfIshyxHkhCM
7lkaua8kxeSPWSWgHK4sU8vT6qeKupPtj9jxwu/e0SxvxvDXFSQeB1cM0nYsxi85Uono31RiIcx9
kQgi8iKZ1EmElM/89WEU43cBxoYglXYMQ5M+NhCWGOS5uzT/fXjc6WPAO7P6n4jgE4ViigTiEW/z
mY7LRYg347yk6xF7iwJUaf2obU3t21X+CmHVP1QFTcCj0R6LS96e5gqfwm4qOxh5WGnygEnV2utR
s77OXMfatZ1ZkyTjhu2fmU7MZvXjEDAbvm1uxTsAEAAf97qluXgC3yRZQnH+iZKeyo9qQAky0dXJ
gFXmk9J4x6N6N77l0Z71Fcr1mfEdchDpUpvHRk+bhM+vyzdA1at8ApSneB0432CY/gNfo4ve+imU
SsRxAHZA+Vve8OZqXifHMrXAughzLo90sm1oBIKyEL9jPcjInNK5P1b9hzVyQyn5FhRjLyU1jRM+
6qem/306L8RaMU99H664FNFPr3g6TM0DPmW2Rmchjmm0GPjcGIbP2w77zrjqOUd1iikjVX36GN26
dLDl7ijH0JW3JBt980jm66q274Qy+4OtwtyyMrCUoUkdRMbimi4ngzT3P6cSg/aZ305sykK49fyN
/QK7ObMtRoPzQCJuZghAl2CpEr/LywVX8e/VkX/kHbgAyRJ9RBhMIab2w1HX8Z0HJs/UigVP5Cc4
6pFe3yyqXhhhw2yIABEXh8+H4j1tapKtdj6H9RocyB3/51sNj+uKL7XYEdD4yl/jIdlqPkwq9ObC
T0cPa2kAgAxe/5UysTPVPdOM7iM89W3b+Gf6M5Ux1YMXqKztiM+lX4dvmE9iM8sq4NCqI1rxmWLo
AJ/LaGzEDrxkbmEnrgnPP0x3w8wSkL4Yp1Q2vP+E1UoiaKNuxv4CU2CKDkhh3mFD49poLUTZArlp
O7cbvyU2bSUTy3MU5pZ91G+DBqSe3tctz0nc3lPzC8BFmcVRaIofZV9SHR7xd/lxYC0aHB8tF0Ig
zW3XLNJRn7RBGu7pVfFQoItWq2FAsJAYruWXnIA8UITm6DZWizgQO+oiduCE8+a2TjstGyGhy+Qx
SjgrpbmMOY6SVHSVbhzmLTdbiLtK7aiyJwoFsxmkFpAb/eOfAAsohWyvLcLbImcdyVXsy4P3EGIV
jzzM/t7BOG2f5U0LspAKiPB2mgXlcDcJH+mKeSSj2rFlexHyFDeC5hNlpD211Dm8cTQWjonMv3Vt
dpK6mqAl2lzEhFbRgDOxgO9z41iwur9h90i98AqhiPl13oygDKEMhg+zRon4pcyIqeitOh5SB7Q9
5vNdceVxTJiIiaCsrXvUq4ZyFTPTrA++wGEhWitVkl9xoPu3hvY0pqUlHJ5DeWYpGnbruYbqyaQX
NwD/yWZvKjcPSV8i0hyUpzF5vGFeFIvUwpSc9phe0DXwaMuy2s/JVwsm+8g4JGjL8WxHHsS+svi5
dF9ecN4aEjn/+9Cjk6XNcjaPYBKYj8NT2YvxrNl4eULFYXskPFrn8SP/DTNZRMDaPgToFkl1mqKP
Xv67UckCrUCwEJwII2TcTxf4/rzJPNeCZFuhZ0n9/AxSrBZO36qctA800whHJ13JvwiaDqdnj9Ai
LZNibxq/jLSnVLOvpdWUVF0GfS2y+8TE7gVbDEbAKsjVZ5DUo8VaTQJsYpMJiR5nPFyrjpTqQlZ+
Nc8sf+J7JMqpfvCYvL1QBWrBF9du07oox/2ArE9IesWo+OlyiGmWQEZyrXXn+VzQTDVW8nK2DoTK
AEhe5XaFsBRpsDE+DQiE+YvrnOeplvfcXkKiN0IET5daCdVn6coAEBc1XXe5LkQbUfPqsbxuk82d
cVF/y6wHW7RuaIucTIKMkT8/mCA3NKhPVHAeIjmNzjEHDh/qzp3EqoYrAd0Qo7GpF4hpLSecndZK
XccqdHLGBj+iRVhZHxb6DhOz6i5+3RxM9mrbjdvp8pGQED3DnQjPifLFx+MqqTsJJG+9DM2Mdtx+
U9ErPfRzF3sHpMAUe7Gv58b9rIxv6nVhmAYk+JkqDkmfBfApimzrebTB+FJtxahSjr/soHPrX/Lh
rQMxvK6+Ml5k2HELs8ikqlpgMBRgwNN68L1KgtzUF/n8KqlTJfYq6y+a8eRIprp6eA9oQylnaySz
WTbP6kMDSSDU7+/WYtQiH5IPowDJU2g9KtpiJ6+GSwTBB5bxtr2rKKskcxZ8t42zJGCiz6hbnRwM
SufOAFH2SJG0Sv9S4iUEtsUyGAff4eYkGz2Yyfs13dyyzcnRhbyBoPQdCPyFbwL2WPNZ5BN0CYJO
HYBpjRV0ObOw9CUEpKL5az+wmbjJqv3qiRZa6IP+rSaJVIFAGnlk67IeZRNrZHj+7Dstk3LXnuly
yLso4Bm65pazqTf/wMDUPFl6ypys0I0ayBm7ZRvh5LfeLcXO7vIG9ZDPNVu5ZN1WVN34wOWBL2IA
qPheQ3JmIlouQNRZXdXu0bkXgtIhNiUGB8foMg8TvGT9Icx4Yz5vRpCzZFLAXTGkzjXaJHSDh+/4
rNlCrrTzdlsfm7FShCSlFBFwtnG4HSCz/qyoKV6TrkTE06hLHPVsMyono7phScCsVpkT5kFxnZIZ
rkJOTu696ze54yA7CPdWsUrZfRsNyuwHEeJTizVvvjwAHGRNgqmLpvPgIHSRQH5rKPwBMtaAbE7T
zcrPH0WikTqqUR7BvH4xuAw0Fi80Rxd0DH9r0iq+rqfd4tDW/CvhmjPFyaczbTsRX2fKFrUV6TXE
9O8JKb7v6j1hwK46KxXIaC6/vMBr0UWVdNLiMVNk0q7QEhxMUF42w+cPs8e9wf2HuH6U8UsUX7El
1yxIkziEOkSP9dO3xccUPsdcHHl/OjRU+VUDELDFZ8e2UvtY/CqCFA6RDEJKbQB1wIgA5FsAESOd
G2s2jVs9zr6Xl+Ly5p+zxzyhEIlvhK/PxNgYLV85BsuJ8kvJTy9+RV11i7fTAyTF5Od1QG5Yh0kg
CiRQMgts3Okyi8fexwWKNKA8qX6Hu2t12gTYjcz/LaR1tQeveiAKk/Etk55eCSN4TdHO2HPQm9F1
7LHL72hH7vu1JE9nQK/TLYPixkOj5xUb9PdEaM1ClIyT2ZY4Q5/8AjTMuKxe47Orl64BxDwnLmJ1
IbsIXwOKuQbJexhMPb52pqVcc+VsEmbgnM6WfXhAyxFTDQttLyyLYblwikk9aW2KrJnor3JufQzP
MtLsLaGgYyo2EbK6blsLNl4gefNORszy3QWjescGdlP7sD9admDnA7wc2UdT4ILc6kKF9h74F6We
i2RsrXY+HJUraDYMLe9DL2Solht73co35lpOfKKAImiNG2Hxa8R+UbnwG7JRmYMekz01/CKBefAt
KCbuHJ9pdl593qffCaUnN5eZX8HaIhd+u2lKKHE9RfsjK9Sq3FeG8osP8HwTXih8PkhJwbtG7uob
ab1gyERIaa7fX770ftzI/WMNVRM9pKTTGxhr+YheMOOr6J795LmC2awGLsgFi8boxwc7WkyUvFQi
KK6w9ytOYObH9rmYtzLMsdFgHFlpxf5T0rKaIxOkKSwixkdfH8K0KkKl2EyttBrcna+BP2g4LJI6
4rYYUbEbNDAOE7AbUq9dhWa1czrdrcFQtrzezugPZcvFqrVpXHTsOAnA0iI6Gq2eR5IFJ9jm/mp9
rFXVYu0CcXHCg105woHdLDq4HuusnlmtiXHtWQiven5+rpyWhlIpvCJfZCB+w9XgNv8HHOsHLYzY
zuRt1FEsquriTFJPtND1bsj3wzzA7xV8tC4jO8Tr3pCrMLRuzyuFmqiKUM9HMFAvkodObZdxr7gm
KP/u4oJ7b0G6XaP6mLw0mH2gYEEzUEGfX2EzdLuQuCcHT5lLQ5QPxmoYKa5cUCZmHLK7Hw2c2RIS
rzyCFLlBdfZvrl/3EI6QndsXLJl5rCbBJbQKgCsEXs+glM3UELWXP65GeDSEwY2UE55n/s4I9fYh
YlZXYUF+R0iWTrrDINi9B2aQFqTBsbps+QXrYqIs/JeKNkf2HrXansB7fHlWhO/7CrcZ9h3xna/m
yYM2Yuh9VgJZkrLCHexPEHMaw22pZzp7V+Q+9pOj32z4Lh+WOjUSDZXLnV1SQ603P1muDkNL9GK5
xOllbrGT2GyD0N7KacVjfTRdIP8CaO7nP1HUVhDMnb/hYWP8iWqwvSRtNaTWmEU68YTap3lEXRiK
kKLojK9P1fCZlenR8O95CYLrzCEcwScjXVw81RMqtIXtAm03FQ/6+qFCQNjDoI4l8QAB+u7jMb6f
FLZqQ3wZ1JnPLmEwJAtkVpA9fJF4j8H8AhMf4QKIGBxgMat5OQXOPTT0CuVWfzyvpz3p3NyaSWJf
+SfI3JaVNh1eTxwr5w2kdrHhdFkcez3HqRLS//1ie/AZhCptAgAsQo73FSfGIAYQrfghDuQyn3Tl
yM9ieZt2l+K5wZYwkD4ZX1d62eAjfEv6LuwP+VtHIdfPlTU6MFCXoy8J8a5Mi++jQNhUdxZE4A+4
rVF3CmCelLnpBuL/4ghplKek6O+rFkTMXDpnbnqotB3F+uGeFGMFf0cgg1duB4u7A7bRIgYpyiga
VSvlfM8hJm60EjEGVYE+17zuxiaCwxfKILk9GowOaI2WdBUBv1d0lnZ9ZlDm0UJxaVVNlchpxcaH
s5Z5A/E3dwhQ3oLHhmMvpnhS0OI1iVwn6GMChKLy2G09tDSr2Rct1pzI7XzVfiurTh2w9hBUdlzv
0Uep7Fnk7hI3TwEm9fmeevHUHfkiWA1ToE+N8vcyGAPDR40I/OD9e51fTPtuqHVkWsifKwkSOXlB
fTDKP91Hd/GR3xMvknatQcFR+PNTh5cutklkLQ3y5UQfk18iOQopsA1lgY+sAPKzwpijcUHZ8nvo
jTEaVwY/usQI+pgTGB42RDC+jOeq1E0OQ+w/JB9uImR4mX0aSKSb0sk5iKMo6ourEJhJzeAGTokt
yKWFp1h2ABMZG1BvMqtnrFlEoWDOpcRYV7gejbNtdOUw6OtcKEZM0B/y5ukLUvwd2PaPZJRMiF0J
AGleoNsdxpzGVJUOxcsAQFg/20kpx9PnyriyF4ozfsi6O21uWrJePSN4fz/REz36ePQdaYkmA1hr
ePIl91i2tu0crv6FuD3HtsnTMdn2UWQij81KPzG9ci7s6aeiiJy4sVZTHt73/hrlUGc209VkH8F2
vAMLD6Akv7blhpJMvGSPCFMEImcjH8itF126wO0TCVUmwbe3lSnd1iX1vNHcJ0p4qHY0NfyFauCZ
7vZolOyCr9pNHq6UIzwj3mpErsOkzEYJ7T25Nz/XcHkB6Ii2krWQJgfaNgqhgDvygQCvD42NuHNI
wMgzPDBMK2tMYlWCmdr3NhYYxcvIDj0L/xiO22NDZk8m0cCdZ7RIusVjW4A6zK17U0+ueAOZRbUO
Mz2QdMftNTn4VME5d7I2mEvUD/jll1+mdDMtuRNU6OTl5+fmQNeaZqeGq46KeDm0Uc+1Mj4RmJun
FJmU0wFqAbCYvHTzl9GNTw4Eo9q0CnBtP5fGcH2h2NVRykyfSnteIjh8YtatxTNBnLryQTVn9Y2T
kui+bWJQJxz9zT23FSMANg0gL3zySBDUKzLXdePH2nTvbIahYD2iH/mSD0Xc1MuHhrNdnjPmfU3G
fH9eJZJaK4na9N6PWxRkwOXjx/dC5CBGkkwoodS1AXNCAlhDiKkzvwUODy61tUfl2r35v5KtixrC
cisQQF0lXYDnPhNIXSTdLEnWHWG3WUx1AlFoEyQQP2i4VQX0thTXRtAJSSOvzDWlCU9k1dZtu/9N
RG+UKNmL4y7U7kf3K9eEJ9dybWpBX12yelE1aCKDUsYh/PzQyrGRnwNRu4LHp3qFAXStXjzVlsgv
Yeti++SIMoNwapp0bwsTcOCv95qaiPtR/YEfRBTLccqUgwLhZ6/ycm2+Iv00ApiW1x3v/eBPWaWr
Vo+76hpHRMq4La/ku2yKbI4F5U2Ez96kdFMbtdffPi4hAOVeH5vLBpNpB/ev+x4ZJ7XXu1WDT96s
ExL9Jd2mLKlljsCZgIrhIpv6lclx3/LcyRKYVc+ecP0B9alM6/vPp7bxMRVZLgcFuLemzn5Ywxoe
zJkgXxh6U9Uj/mPRTJ9HOwI3rhqpvsOQY15ly7nKOhbN7VmIJ09UKW8iQ0gMkl1QP+EgtZG/XzYH
ZCyMGdntUyxAz5RB5mzCcHkI0egLOBaOdfLUVD41e0EfvXo1UQeAp3kzEX+NJCe4sry4+H4zBCIT
FbSo5v9EaAwv3N+Qx/vqP7tyHX6e+aAnscG8waTSDLmyu9yl3rw7mV99JBtWw59PA4T/BaOMmx0d
h0ye6OcKingaw8b91a1QDokfynWaTVyylsC9I75PerU3ZE7C5OD1oDX1A8xtYWp+V6mfO2injujP
++c2/tg2KGiKATZDDOxXrwsZXm7AlNq9l7NYvjVH2OMtYq/T7otT7ONSQqLkXfVZQIOy7fmjMg2G
dCVObBCAK+uIzLAdW0ryTowHE/1yNdNpZW1pDpGbUiIc0gou3NY3O04fAx3qXu7/8gulw3QRMgUC
YBB34T1kZzelpbv+KmjvhBiQnJWGimH78aVuxf4O+Zf91UaCidghw6xdPaPTkgWxCMdD/nzbQg8k
roH8oC7/SP5sScNL/oFV/wkTdgsUuRXxrnavinVozGbzm/DdcWLRXigo3goZeH73RjRuC+OzAXCj
Trek39FMb/zEg07XKwzQNKYGTH9HPz1rWjIyOENuplE0mHp5WHeLey1urzvmbp5A0IP2RaQ/yVRf
SbCzB19RczBQYQfWb2hHvruTrJQb9+IF7xCHxS70i0IdxS9qi/ufPmHrn8NV7t0BAv/blBPyffPi
zGfl+B4UGpcp1oJGT5esrblF6nUdvuZP1MLSq7aFqEWgFZ28LAY6LE8KtlztZfK3FcKylZoRuC4k
cXHIufninTYTYriBWRve6p+fnJh8jRz8aR4neZP8OxsWRfj7LfzBuoGNotKJRlCHxP+AxaY/MUZ4
5bgNcp5nQCBorS3rqOOoQIMiY4JliX+h05vo1TVz0lVc9pmpxeofBpE21hcjMszRfaPnN9eK8PWi
VeNmc+lKIQHZnxNjwQQquVRZxdN5pQTWphi76OQXsH4G383CpB45KPW4q4grSVXbeE/NDYhF3JF+
aZ5JkzX7XRVTV9TqYbIWY/P+8gZj9yprTvuIn+0N0bD3Fv7Cjgp42caWnjZcyI/ap66hF+J8m8aU
Fn6f9gaNRF03wY9oCYTz0urrcsBJWqrTtczdtg0yfXzN7v2y6ISeI4+an/93bNzluZ0QVd2z/9Ok
GSA6CI3nB70jwmmXyr3W48iJCuzVBMF3nptE33kkOoj7WkynDJRYlfF0AzTnABUq2H0WKd9Q2vNQ
y4o7IsraN/Z2W6RR0e1dw5Y+K8gqoI5qJY1d0rvJNKtt2DfhMa8pnjiY3ceJctuPX66K5Bak4hf9
6PaDbLGvlIqKXFLoAWb8HiKfMTojidSWcZToOayL+Uh3ev+MWZt1rXN5bxO4s7arI3e3vX+G5uJF
7fB1XwZoj7VqKOnwqeR1Db6PMT4Zr6tBBrx/QBg83MlYgYxcPxtBCMJpnYYknBiPLOxBJeJT+mck
tT3n0CMMgyG3wDMKjpmi+WABQiHW8mMGtWUgCcdvpfVOQ94pAJGWvPC7tqXrXZgi5Npav7pQS7ul
zEIOfHFLrqeHwxdISD88o+C4pTKhphcNPjyG84+btmBRbJmqxt20TSAz7f0gmgE0QcbHq9MwjRNe
7AJnRF+IhXbUFM45EgobT7dcWgo2HG3XXl6tH+ADC6HRmp8ajPeIzMuNLyd6FDyjgbbC/Zwi0Yk1
VQEYGVYNUismG2GfmzRLYcHx9Y4nemqCq8FVAoVDD/VUApg5EZGXDzR9HXeKSE82O4ad2KLefRGd
//X9MrLxdFH4dE9gn48WLh4pyTz6SwgctZHfQXd1lwQFie0Oc1C+G3iYj2p5Xtvd9bTmMU6iAh4W
4EVTy1fRr4k5+jakMjpHcTO6YcfcYjyknGB17rWY1In8XhPA93MOyrPLZA2xG0uCU+gNw0JsHjm8
QisVtpadXYeM6OGe39dIwS4mlIKvCYRLM93wwoDsWtnYiP2EeBPBNLpMlEbyeahJfX2YNzRpDn05
XtZSj3sMu70BdhRYPQJ4gF1rhupawXxeIp5OHN9YMky5Rwp1yLc0djtwZXWMUzI7pL17WxfbN1bJ
He0MZx7pXAFuvoC6A9vUj5JPGLFGqFseFrqZHsxEXNo1VNtIPn92PUU3NmtPhRP3EGP/TgVyxZts
m5lQHKcC8ueMqNcNkfBNMzIZ9ATTaaDcZTgvuZgUgGqOpbIGtZuc1n7coIS5R07jtQRL28PRWH6W
gm31Foc1kS/0UuAOAm7SUkI8hLpF0THh0J7ohVQHt2xtAlB2Flv9DpxzY5AFOPj7XQZ1n6HtX3Un
0Z+P3w6+l7WokB+IR+lL5VbcSSOotcNJkmelGLyyCwXYR9JVq40B5vBPbBaLwsID9UUweo88P0iC
doIKMIfGfRT8Ifw5l8yYpHYhv6mz6EZjm1ubXHMUaqma2OhvRI2YtU+owXC2Ns4IJa8vfJsQck8C
M3HpoV0UBfS+T/MQ040eH8MvRFvXoMThKw1IQpeCB17ZUMkNKEN06BlvMGzIuzwjJBoTxSxKvOgW
SBMaN1LOlO7q6QJceemPouyTeO+L2DcXCXEPMejQtnVyfS2IvVgYfGIrlDan2ZMsIgTShFEGgMHy
1uKVr8LzYZ58xwUpX44y0BkhdK77ucLIQz7W5OoGzZ0uPz+BezJOyzQRIJgtQ0nwA+FPbbht7d+u
Y4BBdXyBO3W/Yx2ELs+uVweMy5RD0WARJwVNiYr1s3VH00DpYJgPWV4ywCMjQk0wJTfvSeAkVisR
+1NLM8JVDX6bb4Gw8kJFyW4DVW6nyRO6/iyyKmbw2t2/PnShtD4TxniqCQGlyDQG4jzaIT/T14JW
/KTAQ61F73ggC7JZnA3J0fiHif2Bf0IvHpHRx3koqGQKcaJvfL5lWg/IHqqilj8sjvyu3FKZFdry
owRwPumKrxaLQpJYb5qs/2lOtEG25+E2trkRCvA0oz+VDjDCHvFDCbRT0303jL6FUJzuxV96bvsA
9Xk3R9KABd5+g1vtle29hG8sl/5XuoKOHb1porn8+KOpwZWI3Y2FktUrQXFdNyamESDj6gucbzx+
bJpE4jsf0F/eYdNmNYh0Ws01CUpRBGSRb15vG4YOUW+U3ckGQzf8A74fdnkOIUGi3LLes8pPYZzt
ITZ7QTbGQNbn48glMxh65pVJ6bqJ4eeBdiikVvHymiW5z2o2ECKD/Tz8l5RZYhukrCj8BMGlbkpH
6po6DMlv+AwJygGIVyMFUUKLl5Fz7kpx6mh+0H/pyjt8ai1aqiLexrEXGEjjv/qQX7IyUF5JxBGO
1rRqmuGYr8o1sTOtdiANvWOv8muvzvJiUL8jwr3aIybQzncrzap/YAik41OZSdcWek9OlHo6KRfp
MHYmxaKHEYPexcLHoRAaGvD5FY2oivOCNe+IB2hBqvlH4rKA0LFLLj8w3wV1rl9F5ZC3MAl0SsN5
F74CxyqsqhgHt/F/qmG5Qy5qjqkhp0B/rqaLd4gCSL+6vEh4RuxqeSFb40BHrJqJrv+rqUnfAHrH
DE0N77IXutrjjdmIrBljnnNiRf9sH1kPF7VfW+SXu9WKzkXlp0+qCXWZF9sC0qKodwtwqlKF2PlA
NW66cp9y6aGl4Z/8FSfqwZqso5DCK0S+ze05WG7/KaVKXse6Mkc/HYivx0NCpswinuVUKv+5v5uY
OzfJtUNDuvOb3Ai0bOCKWkwYali2oVjz5YSVzBUxsBYDnW/99RCPpAB0QcNnjgnEapBcdmloCfp2
hUPl1c2se+xVqxvLVexYiWaRxQu/+arxTVUDmkJD/HviYuaw5ZZlIH6fgjzeoYa3kIFG5TWiAmM/
AuOmHKPgWZciuyJ6ewjGXtF/8P+JP1z2U/NGd+A6c+XF3BI2bXj8xvI4262VvYW4C0c4J3NRXh0m
NJagLnidGsklsrpqe4Ckfngj44M/Fsn+OiLh2501f8HnxiZ35/DZZ7rv6G5MIA5YFSI0j0o5HWhE
s6JklTiBvQgpRt0QkwT7qR5BaCExVW4ktOSgWKJjpMWu4NR49Iv4W+xApumCWeZDgamU/xgFgiL5
gXsNd9G4kl8BLiI76cZRVeTrfg9C55qFbX8AdFv346tbU9P7eYicRtvuAGmXFtFTROZ+LlWYmq/f
LfOlLmM5jrImnz8vfbefaqlp2jYAbt8Tk5No376WfNTZhT2HztnnX1W40MbsOBwNVmtvtsKiPVML
ehZFMM0skrc7xL8aN5Ohr2XcENqhMW0wKpKVXiRWrnO0lEGBVh+U7zdK8NH7eEFpXuayhlkigSpm
pvKy3C5J3hSKR3hRLwgOjW7gZMTjGdaaIJrweSLyWyhNug9bGegWLwSbcYfpDkqdfW4SSTEJAhNe
7OsvijkM1h86SOsUtoVzsAJqFlg+n/7y/N70K3Kt4LF1V3t01rtGhXtNtNWoal882EbHYEF6g5pU
v/w/NPm2CQThkGx3LMXHQKCkJKyi79828pdHsH1tXGP5H9NpkgSDuA14lIXLbbd6GAxg2eu++es3
ZZF17Q3OZB3i+dDND/Y5RL93jl8/gq8Ug87pDncav+4mHhimNfFDbeE6WI2RdkGookwuthJ7BaSY
yxr8pCI1f4XIqNmI2hQwsyQmoWl8t0qf1FbOq9SzdCkppbgqnuPdvuYuG/z/jd1bWqcqRfZoB/PI
4ogXULJp3wlna5MRzavUvqL+fz5BtIyWiyX7w18U/lAa6sDClCYTMZgcPYLspKJRiTjy3ixed6vl
p9JwSSL4hePpcQZ0wj6oEu8DnMUN/TYz+lhx03mcMy0Hol5aoQUpYdDzPEbS/KmaA+u5RoJbHrNg
fJiIYuB3ELqUtgR1k6iXfoyovzQr8ab8bdKmIyF8aUdnDEpCCHCfsfUlllSti0vz2yF6v6bZomaK
e8wHaS5+OJn1UiUqypTMv5W4x/NiTd3MzotYI/iqkSpgtlQ54hujID+uKcAtyVORZoGtUlQih01T
k3yzSksX8NibNv2pWWVxCLnQ5lN5fN4ZfG+hjJERKIR1U0YvbJ6gMJD1aqe7MEcCqL1/73C2spkp
xUKWLZb2FSvLDCbPRW8t5cs4eXcg9QQxfx6Z2NHCrwjKwETk34lHLOxhjjiChov8KCDYp6cIhVoN
RNJ9rVPJ28qc9ad4fPfQ3VpGxAAX8wJuEa/scLxwKcUhvztgOcjq1yHz8EghatxrY5yY5vm210Kz
fFaNQEGUKFLlg4Ezdgy8reRdaDN5ACgU61XIs+4Lj4Eveq7JXg5BFAKvDxsp4m1uMgy3aZiirlGt
FeLw8/3FbdpxvLiUkoLoxSfvJrJzxF795aNtDfgbLU55si5IPuiJ1OrJ+Dla2c53mzrxc3POoiGz
kC6EhnPNg8X7PCDPdXwJlfR8YAUZSvWKxH7EhbyPs2VdF/4+36sZPouoM0lS1E9zyguWklY+oYlG
CKJ2vkwSQoi+gzv5iMBi+VWJS9CwuxoO7d2RQZY+aGGFdZ/brT2aUuy+ArWY42hI+ty1N0kCin3a
8V8wiid+jUo2Ap74qQ9si7Q8m9pjS9k/4y6KBMHMu0FbavIxdIJZz5OWr2owsNAf4DV+9E+WydOr
Y8xBIqbM0b3FRwYFbddKjRFw/Vf/GXvY6ys1SxYIHSGg96BYGcCjwoCep1M8l9mR1hxVuehuGde7
aiF/TYjVpp7qt3cqEV9tgRJ7WUWA9mp6YQDxPm9m5ZkjmySt2uMEvdqyz5O91o+QD0cNE2WoCpeK
EyBoEvW4CtNgwt8LvSXZ49iPDUwocF+MysMhAd3tYaDdjerb+6rOUYKratpkXhyi4zjslfm8SkA9
ej1Zi60b5F/TTSba5eESbLnbFyfggq/fhfFb/HqTV6l8bG1gJMo+THCu+mat1lc/junFyDo76bJ6
b6iKAxCs/Mb92u9tJpNr6oKzWesfL+5hDsUFa8yyLEw9BYgQl5VUsUqKkgUT4XDAj7GnALsLMQhc
rBpt9J+6LtdZCa4LCsvVAiXwlMQmlCZzUUj41cxTYOy3qG0E0bqhpvHnxGYKOIxb3vHSeyJTzuDq
JsJBjfLQAAN+xcw/+AHdhiJ973ZC6kjIWeYbscq4zWli5+eQDywnwC1ygnzLtSoat71ab9xaEIQo
r9OMGYaht+bNY1uob9GgTplwGhd8Q59gFa/4lgt87PhM1zUYPYp3QzmA0ztyXX93PB9UiwKiwd2G
uR8HH5PTqA0JfHeiawluTnCBQysEnMw2j6bOCYaU/0XmTp8LRdZvLXEYphRA7yDFLiav4H68UYfV
y6ckB+GIuFALGkTIFYarFEd/8U7EnXjq5UpLQhF7vvqZjN1BLxQ64ol19RIDm2sBJ6flcO2v3lWB
V1xapeFfoZbG1zlJKisu3mvLYnUDhoVwkKjOlaC4w1DYLJhCla1uVdUiSaAJ/aqDSGbmRYaULeQg
3m3ya8rIBXetOcmayaf1MwBOsxWCSvGLp8Y83eehMOCwt/8JMBEWUMekknJrRrxW1OXWvHOWVdzF
S1cOPzrAbB/uS+qwEctEffuZ0smgAJANrsWaUvNjhS9RzQ0OdWaJd0f+LMMZqMvdbDNO7p/BGPy4
NBeGpQrlKYVvAgneM6u0FWROQw7jVcrmw9tFTv02D+yxi7reBYPNzDa5d8i4IfHE7GU0VsMHgU//
Vin1M1/0YM5JEXr9vAdAB+Q/E3Z2VDzsJAJlu1YjM/t6xk8fF8ugx6lMGV4yqeZJNM/0ySDjGGNs
E2pO0gL2KAOMQGGiNh/phSML7Y5KYWcfJh3QQm6mqdgcQI3+FBkDy9oEdW0bLEMbzi0AB5eGr82q
0SkO1NWhJX5PR+HS51JHRvw+rpqme8LZZVpntN7xdv3C+fbf2Sh+ZvJm/zVDn05VCBw4CBZM2Lh7
CjKSX574SbczLP5uKiQXIbGsjm2hKjeNzWkIqwqAHymUNma02Z99BWUBEn9U7v+4iTPC6lOg643A
uL3LCiGg7fB8ih9KK0Tp4NyVUfosaIqHCulSuMx6rezfzLx/d1X0MGhmtYK8vSQ0HmjysyXH7vxK
TOLtsoUXmgh7S8qwYZFA3fAVkFWS1sJrPR/NIPzkrocw2ddrivCkWbXYChl6DIZ+O7RY/Mu3DyVk
v1DswQtA/iutTTsjV2pfrR9GjtayIvga9j96FE1zgfqGBrlAcpPGJ/QpKrvd4HT+0YKrWzxspwJp
tj4emSq2Uq82HwgDlTl12t/Ya3RyY/ldnlZEYi1yOS65fty4C0GqgD0TWc4N97YxKC++hz48N0Bk
bzbH0bUrXFRZ53Dout1pv+C53fvSPlDalwOl7ntDabUaEJ0mV8g1aSZNe15GfjbVBAspgP/Du0GQ
CaQcefG+RL1IKb9TjhLR3JFWUMZ+jOex4riaIIWLSHaTAQpgDq2aaGINelUAXyEGTRw0E7x2fPuU
yx158BNxmrDyFY/f2kRAMoNHnzGlJYRpk4u1O8PR+E/XgprU+3itKJvXmsQ8P4cUdDev8+Hi6Hlq
TnApKSiCeBVll4Y35o4kLm1CsLxHLjOhd7VX9ZUPWoXFFK1Lq7IlKT6Ub5mdmaB5ULdtAqtkbAzJ
DWis+KMlG8YDGIpcO18XheWR9qvaKzbNKsnNS1YxLdHXG0DSrkFVMA/gSbTJRbc6Hq5FMTINa/RV
vKjgeTxgNWNcsQ5HJ18JpdKKyPnO41U2N9jr9kWrppTNmwvqLMRZdzhM/btA3ZHk1Vfs1Dbyu1Rv
P4Zaj/7LurdeB+OxEgVbfVhAnOdCyFKInHOgznKPFWW7kvCUVcmftlRN8Qjy1ioQ9Fhll2mA7CTm
/MguUF1FMiPRySQE8LRmJF5Vhi/0L58ZOHm/mC+9RX/aIfC9EctK6prdbJI8Zd6nHmBUH4mwbELp
mAYUxOOwJ54ZnfOM+8V+CQa5sy++9n1CaO1fG48RbtcsOs5z00Ai4IE2pGTuBqyNCZyaeUd+CBHM
H+IE51SmzYnOV4WTe+VA2SmY5CTrhgjPpzoQHDgM4jDLenEVYR2CXYZkxbmPOuyCoUb2kJnwsfcG
LZ+0DSMGd3OzyyN3jDZnsJenGc81Cffzko6LqYALDryU7NGuF6alqMmAgqdY5YNaKiq1DKSQ1zDA
pmzJ5GyJcTeZ4+qcQXGPwOswflMmKxR5Hss8fwDjAbZ9M/JhdSzTo9wI5KUJSOL6dSnhV1qmc+hs
Mt2/mLI2ePSnSYtX87i783A3e3clQ4mN8Ae5kgSGF/vp4DB+DRtJcycUuPHCJueYLp5gefGla4gH
pWxIm3YpGmiUp/UX7OiSXpO615hx/M48TKVSKaI+uRkpfWUsV98p5uS3FU7Qke3Y+cJVqFJaCUSP
GTIJWHYIqTCtyiZrBIRbT+zftYkcYXKffEzUBIZvlMJcLYYV09godKLiIFPJszA4PaViqzsxdNoZ
WEacp/B9cGRAceXnKREQ6/pqiL0oYDEuPdT4ALUjdUKIUaKoJsf5JElSH4qukgDVEykxztvgw2QU
9iUMsw4CVVUwcqOSYYv5jgep/9urxGB3xXL225RTQ0jQgL5dUDEUhmKUj6+MsZAfO86FLDH5xW4a
vaWv+FDmEuyKlJ2EUz0cE2FeOBSkg0muwxpyscM8UgcnG14rL0NSZUS88GF7ya6t3YI9FkELCurV
RbqvAzt7Iar3ZiwPjI5I/WHZrrg6CYXkz7lFRXLC7lB2BPlf78WY2/EB1yhxqNbp1pT2HE1fzE18
dEL34JaT1Tc8h4cvBVOfzw8yvV2UQmrVmhU7BLAnrWuiW4qLPmLU97YX41V999GOdGBk5oKmtA1y
8VPTaKePqBdIWYCgyOJlT5fQNYeC1rO4rWBVYw1kkK724J2q9Lfopt2+cuZdOscHgapGzYb6TeCe
Ov1oe9PaXeq6KbqFtGmAw5wEpxbo8Uv58jMqY8rheYNRbnviEvzmSUunVV9LhvB6ujar4oq97ksF
n9DJ6IA2BX3pU4LtVGIgQ40s7ErKWVXNDYs/L6pCB+UNeKiRRjmDLmDlDyeWCzo5jC9T9B5iwBF1
B6JO1977blF2CKtpr0BrXOusJCp51nhqihwokMCDvYB8sZvJvEdEvCIraspLwUmvYcus21xrcsU6
Igh4uSf2gf0MQIehKdYCjeEsiaG2bHMdUdCougp0MDM2uxM7Rh95ynOoemNapWCQ1Dj7fK5BsReY
C0z+AukMcrjA8z2RSJuk36lk8VkjZRITAnNsmiiT/xOB+JAAlqEPb7c/PQxH75/8lkL1IM3OQy+o
m4El/IhPQeR8VFEmd9UxehhYd1an22eyUKFUU79uOt6V9oImcjvnwi0FoLyEkZg12LDyjuE7tPUY
0uEdWbONMrZXidKpbTRyEnqwEtE926gQsdKZteNCV9RSPzbxfA2IeNMKVlU/W9sCIHcuNk01PiOU
sd1aM4Lcv0PLED5jP3dkyiEXSugB9hdiEmtP5dY/mtGJmQS4MamwlCEGWYwnftQ6S8djeLcNxlB+
j+JERBRGbz2P1lRsUrdJgMl7/Zm0vbuh8TO4qrhVPd1Hnw9DUdNcYkbDVWPc4P6GDAD6BdgUhNzn
12545E4D+qBrX80Q/jwMBX/3M72CZgsQ3D5NuqiGTkCzINihw4q01+3capSjkRtlJUQ1IMdP+1gl
ZWf5Bm1EvqWdiXxQFRQvp8y18B9wS6OpTiWUmV4w0gtw+/eoV8znOjHfnc5GN6fR8tuvYJtuL35o
dUt6ybofx2l8DzmWfbapXIGlUPk6pO2eBVXkjL2HuiHWuLGa1vr+5OmTrZ63XBWJ1XRl6zbE+/KK
pOILeJ50bSxxtr+T/ULiRlxoQf1e19OncxKePiYN1UN0sGMTLncfVAkRUyKoUC3+UtpVdus9rvwI
nhe8vjgZbGOnIIATLD8IeorVit20Jgfx0owmw2lWdjIWaN1S4gYuCnH03jxOmWm5SM8LiUGgMCIs
nTTn0+UJYPqOxxXr/c2EEfo9Xs+Y5fnBmXByr7KYxInwNybIWqf7aTgpJt0uo3R8fawol/eLKFAF
qZ7Osss2EpORNPe7g8tyye29GYiqZ591q6ybP4Vb7oRK1l64AVykcxszlZC9JeO9VdO1RQ+QJKnw
akXiQ+K6haknPGiogybXx3n24CtuXn0U9ZmGduHWd2bG1+2uKGudNcKvNT2fbXMVJ/reBF+vsHoE
jVQMDN53vv7OBTndwCG8wZWhEkA8Ksupqu7ywPCpXm56ee8WgKIbvGGTneZMbeoOQ6gshCGQx7us
W0LYXHx04mcF1hGCpQTvNXkCREK4mwxjoDIWrvUlWAb9G6ikJ9vrBc1aznHgJF4lnm2cETK/sjNZ
HtnChvQdpkeNJgCBdqdFWlGVMD1KlHjBcQbmA4DatUToz3elfBY4D3q4NHaYitFM3h8ccUX9gwLe
tDrEwkf203GtSVhL4rnCqfSbaCuyqeJKSXnIME5DywHQMvrPKmVCKNIpfmt3N1yenErLjRjLozr/
MIseUDINR6q5l7e7SipP5V1sl3AVUbq4bxL5SZjXR3Xsi1I8Ynmt/VELclkwlhS9PPoG/c55neMG
5NhGnAxgVjQbRuTYzeoBLmZEyowVicPx5oH0LIPQJtYT637dZdFakAz5FvxIQNIzf2btl2ao0jRM
B/KqGzB8LO2vF1UyQA1sScKlMOJKl4afAkd3vsNhV7aHHfqeeELSAHZmfrglNkSrN4Gb1n8JnKOJ
xvNtD8p07/Ehea+grGPKuTX71i4vNIIq3fqMGHLrsSL2mzKEI+8dBKySNC1jKs+j4gQ3N5/e/11t
9YYPxSyOgF5r+kqFYcapddBHYsW5eQsolTusvDPew9TeqOg2sTyzWfZ4narqtewJ+kQpvXxoJ+Pw
JQbyxMk7jjXXJRnbnbosa1DOiusGBTp7Oorw8p1/vFvO0bpAgIwg+1ku/ZwUD7vNMwJ+6ImBnxkf
ZA0UvIbaJWnnNWuHDJajdjoFfCqwTY3raZY62RJSjgiMKx2RFja5jwNdvjDb5vTY+Bmme/eqZ4+Z
gs78ECk7YTYGvTLvVsDUIl6k8bz/kaPe2sMeqmEuz7X79/K2hHAIqeKHr9quGJXyQB6zkePP64XZ
TXHeC7xxth0LtHn9z+qF+ZwisPnxMjHMx1K9I3PYudidoscSt2MCpzq4k5MTK4LXhavUueK9HMi7
d4A+cnLtF3MflafW5zSB4avcVxbL9JIfU7/D3GjrHLECB8H8tT0miRFHzKC9iCc0JjgIFhAkEX7V
9LLyLpYtXVJto4gkxojNYMffS7aBzhyLKHpV5ny/Yn7Jb4L4CGGtfvoiPK6x6k+qpIKNExo/CC6K
qi3s5afzwtKoBJu+gs2zsGErHND/dVpvo+25pc96rKyYIkrEJAjwRuPGtGirQVurULnE0vtHCidP
G9FZNDlQ6W9thCzIPhgmSSL9tR3t++k/+fDkOHbE8pLD0bn9rupAWiYSTrEhpr2SPAd2MucXO9Ue
5jUP3302CtDgSFVLe3Rqb+/9DAZmJ9iZZWiT5bEFQ2zUGz/WqHgDVCon+Cz22o6BrGU+q/U5+bEe
9C40QI3jYJW5+yLBpldoAvlkRtEwUFkTVr7ZX3tKYN0bzC24OrlatmeOqK/23mizvz+CaebTqUmc
nkzYNKInlUOw+LiIXx1cppK0mLBpPORC2vPpguImc9lD//kVzs2TagbVDJgZaBLBXB+0pGVwniYV
6QLY/JrbL0S+PEmH5TbZoLql59JcPMzj/s1B0jfKTDTyi80a8zV6JaNBNrDxKDjpieWZ6ftDxzDO
QmDOrU5Sf4oKrtqtNAA2YwOqoARHa50Talh5Pu/XQnjWt3YRX2QWda6rPII7lPrEwFxA2LhNeLGB
DD7qJ/MzqJlEHo7FZS8+egdkTjQ54qahc1IOc4C6pKP0B76G6L68fUQ+lnjzOzoxb0C6btWcDhfp
mPpnlJ7jFK1sGWERi6Sh8UV7ntokzAgKdjUALbaV3C9vGtogtEFeawR00DntmZNx8yK18NqRqfZt
NY+5oj1oBAoX0wQZSXZazZbKjT05OdxUrv/rV7tZJIJU3YeSa53nHTx8tqsiA3W/XrN/bTv4X0J/
dT06M/sxIegrxd6wWNFF8ksu1Jz8EdCL3kA+rrIsKnc9SImElnaXFkyjIo7iNxusxv9o/D6yCcRa
lnVT+ewYHRKLnsaic+yUGbAo6ZsD2UHd04TkGcG9c8I4eB9sxPXJrLmqfH2bD6J7aZZdvSxwY/V+
/WzuwuznyjD5dCJWQDcCu5z60S+Vh7icR7hf+j6kIvMuU1rtLxkGp9sribA+gaFK34cVPfA54dK9
RHt7e0HNh1CS2pQaky6EPUz1Y4cfdfI9d6mUm+GopJ866H6eO7UMVVbNe89TVpldzfXk832iQSwo
mHYk1pA5DiZowqFLo5jOqN4t2lFHRd7sw395DeSabqGWfprZW1nnFRh5ofKRKXnZ+2y/yWHOkEOa
LIfcSiFdr/T3JTxZoHBjqe9wbXnWeCELRrjeig0JjCgGdKuRgN9j/9gpVYlA9IHanCLw9W+vn4ge
NtexsMRQlKclmK8xbr5XPM9Dks8CNqbTBsHFF7pDJMte1ywxYF6B1Z6FufWeFl/CofOmehw9wQQp
Eh9jCJg4YSclrs2578ba+bFGja2fK4Hjozf0PrXZCC2x+XzNaA+Dng9JSQsq2UhO20QGju+5kodU
CK58Gj0fyvmZ60EXWNU0ZD0BNqH5MRK/hzw9Jz6/LnnWWN0DkSFt2wEkaTeo2ijgcJCLmmVNvjHc
jw6LFSIb6MQ1nTKjdjm9qJgaKthU6FXUIMm57wEvB+1NMXuBjzIozirtnyYiNV4MwvkTGT0KVXjB
3dy/nNLr07e74yQSzfiou9X8s7rZotjKcBWlTS89jS/3NLHH53RRBVBI7yaqIIvss5oXq3ZxPETY
e6ukOtlfL6wDt4lnJ3xTvgFoaJdptqnKWblAVVIWJrngjzUaqXqgSlxfx4xLNIqHncH5GBNbNRsL
s30djaups+Q4sqnnDlq+7xbRBm6kGtPUtpJuNuZsT/D3klBcKBfUpFsNyBO0DtQTeRCCbJHc+Ygg
uIS5A5OAv49nQ6dPXeAR/y6iFScQEtAqn2VEpt8hqpHkaMtxo2kyBYv3k/cIu5PmQFHnAiqKhVsj
39B+2D+9AdqZOwcHdUaN5SuejswQgFjtkOlpzPDm2+sCwPBHGTHhhR/kj/Cxl7EfX9eEcTmvmraY
k9/XcGZN3fUBbapfU5ujT2HnrGh7Jsq8BOgm6NvWmUxvpQ+j+Hz54eNLk3UdNpOowWBoUIVOoCEN
Qzz/alqReVn033eWLjv0uYILbZnXOjNlrR781nSa/4CbV/MIrxhPldtcMmjSkMGOOpb6zZw/EUGD
JjU/pYuCuUlLG8MIB73JAW+jPCP9EhUHySXXyR6zfNvzCAcxx1ZHzjE5/krd9XgXba4gNFhV8oqW
6oDNyl107G2DQThmj1PKareWGNeKciHA9nJcuWFD0AwsGuvjdcjlvNCBVefEXyAlxtNXkHZfG7xB
oALN6x+5o/UwU3106qMS0Z3XHDgfH9GoBoaToK8/uSE91gUD8z95jnCVnkmPNqqNnVRobkqFReYX
phb1DMT0lzSRqqFyDF7wnTwZwGhl/WFeJnNB3U0QZJStJ+i4IpWgjmPC5xdlR4KIuapLY0LNtG3d
RoJffynVYWL6CfMKTgwe7GM0NjmUfVf++gHvlpjZ6M65rDuJ2Kp9zkBeiin/pIvxijuWvioIMCRd
ZoFYMe8efh0tohoT5CvAqyvj1J9G3ImfqySiNxbNgQ8kikERVjii0PXtS4zLVylAl2k9mx8mfUAO
Hktf32S6Jspj1ApgXBpESqYmH3Ruihb2FvN0tppgN52pOoG3gVorsJUh5OgmdWq3i9UMsxNOP/UW
/vwrFM+hlUayu/dWY76JPr/lhxDW+wlaosW+iHd/iDDK+mJPLLiwhW5WpKMV5FC6mzymtMS2zOHN
haPyfY7vfbvVnbtxJaIgFBMWzGVBVWy6/aebLO+Vxs+8nN/L8vSxaGAwsRaN5D4gQKpEWMgWSz7E
kvcTWtxRIoZNOfl7W/Rt05T1TvwRMAx+CNrO137hqxjIPkrppCYYBmXJHcO6uNAqHrBk37w3n3rz
ywNGkc3N80wPTFepx6Mpe86bs57vPWwIr1QMq0ERvMTjNKEY8p8rZ26mCjUHd9iZt82N5jeU8sfF
fQv+sXwlFGEYkSBzLxQiJf3sJHO0zJ3Gj2Zot4n0WL8d1vUjG6bQ4PNqk+yPGg36Qk4mUDTX/OVp
kBOcnS/Eo4bBL7BveD6E7fTbuYnmYwYl7Ymzn7sTEF6tXtSAiXc0X69Nl8+mINuCmgLOYmVAyVX0
6prInS5WBmQ96K8y3wSq8XCGiH8jLPIPcXLXiedy1KiuKuHe3s0J2lEBvg0OgFUcPAqZ/ykzmto+
Jf52qrEdaa75/drjsJvWhv1i1g6hIFDkPKGdTMIHHpIX4UmLq4aGLTqXRzEWLOz3nFkKpAiKfBC9
hNc5wKMVfzZPZatl1szzVAQQm0wQAxvXHsXGqdxZ0p0ZjpRj0xbfzbaPNll2AwaxJxLWL8DlGmOL
4oSNw7yE0Z21gyM8gMIJwoi7jJozPGigqjwmN8kB60AKbgGp0Pw3s0XPN7GzEd/hjtgN+Ohqi8Uh
6Ih90zr32ZwD4Vn17Ej5+Gh1agtV+VkH/r/zSNTds95BWjunY9JN3+km8t6kurrH0I8M+yYOCJOw
wFJoGsWnNA6oc04VqFwe5IeDeOefnpWDjF1Q1JqSWCRLKx4gnXjViqcU/x37c2t/DJrAygrQqhle
0ahhRkg1ZBz5nr1is+Kai4lUW8UmTbEBlGjNPis6Z5snaIcUbJPHqbRiQLZOzTGBRPouPnqE5HZl
EF9gzvaUnyPy/RUhgYqe+BLKZD01AJp9XREBzeji9IypUohV5diVxL9xvCniAHtqFYqYMccsPqCo
QEM3Fi8n2HffGN9+H2+aiAKyb3OmZ4z7XCZH11HC+YNtfJIv9pd2J9Er1dCzdaV41RkYcuZOLRXL
aUgTEypY9RfYQdHPfmgH+ttVU1Z93QdecjP2OIXyyArX0K14WfxV/llj2uw0oXeq7W/Xp4mquIjt
v/2q4UuB5PEwrhdeQL4ramms8RBKIGEgB/lxMH6unoDkOmjYXl7INVfeWrlKJsgtXNVlfk2xeG8k
HIj30gCTQ6Z5nagWxzi1F6FANM2e4mnRxe4bNj+erLA/aiHrE2Tyzj4kZhc7AsBX3i4PHuPnhOel
/UV4E5aI9A8CpEVfvSVURlrO0S7ulQr1Kck7uHbgiAA2CYlaqq/LHxlR4tx5QFWXUwoHSomnd14j
kd9MB/7hqL6m6oeYM4dk4GKClpOEiYkrjf6IHAw5H/h4PLb2S0pGp+SNoH+sdj37cG0mv/SmjqFF
H0D5FLWTgak8xnqWTJ0IM8fmZ1pzwSZJQYpiAkodi4PMDDGa4OEhJ4d+zt7DEHA0O37Q1IVqPzjM
4FnUi40JfX3qvBiTr+RufbKPCAPi8dZz2pBiHV3kWzA+rgUEsZyqHkXMmz/2cfGkZPDdTKdeBj/4
rPIBSPPxvlqHix6J9paQ/pJ0YkVo7+YGKuyINLmJgOD7bjFe3DWsr/syOuQltrJx8R55PitqxHtG
geCpIkKo6o54x+wZLTyyzb9SsyQHamqO5p66oDEPUaAucdtUpWTjau1o6tewiu4ipMGc0fKtOTHL
ici3TYEqe0AZ4p8wJWPLRZjI9BjBnSIqoPqIlLk3f/tdy1IzqnxFqki+mE19RjiSUF1qCQCZHaUL
/uffgEMuKAGex+PK/1goRp4DZlrFsG44CIryF2vmJd29HsfAtNFR+ibNN+9LeaHAyiIr7iCs0mHv
4N0TFDjJPnV4/PcFhJ3puuUSr6V9Uc6nqRT/dhdBKg7X5IILGXLmVnqccTwwPWu/34mOxOCQtaVY
aWzOFZinsJeYvvumZXcRTM5pniSBT0wCk49/FdETWypK6dwozBDQDF/VFhzX5mNcw0ZZDP1zbBq6
VfFg7pi04WsKxJi8967x85eoCdsq2jArqUGga5KSdZs9oPnlc2VgrRnlZM7ij9Vb61aq4p5lpizl
76y/oM+TsisU08VnNAayq/d7SF/vITol0dYV/c67HmZrbdQY1RE5VdIPpDR2ww0Z8xQR/unrytmw
xrbgPyS2PzahjkUdjWIHW4DU07RGUcZLWTeUrXAHwc+OhCLtPdBFskxn/4K7EbuYzI/OZuqp4hns
v/vF1dVdDxXV7FV877p4aNZBQxp+RSQfQdbJU38Y7STB0uashkdRu2/NCDw4i/WzBffMBiCibIlA
1Md2/Gthv0GTW8V3kT+1oGvCPR3Czqw8AL3r0MFuks8EwzDJPVVRJ/zIONpnkQsuJuVWRnWORGm4
nGho+oR1uC2OGvo+hTBQlPbjDrAYQzKk+GlM8KuSRsuIvPqF2RmNw3wvpTRAhxA/vVwxtNQSqN4l
33P9QPS64b6Ab2u4II8GhCH0vfq/LUinvXqJKsKf8u4ethq5ttQq8sNmrJ/zzYppsCQZW1EccTrH
V6TvXauHBv70DdprAaX/HQYIkVReJQ7bWGVV7At1mWsfb11XhOhepsTNcuNb2bVO0RzG1uw681yB
IEzOVgndWuKKdh1Z6Z4cuF+ZAw5xUX7DeYNKKKx6yB8QRyYTfm45hXjtCQq977bSwaJcFW8Z4+Tk
VrpxPc31gnCcJ7GoPHpTOYfK2338spUDKkSvLYD4m0SDCPO8TV/hMUEreJoiHDItx66m4vTkbvN1
apVyBhocYJ5tbkfXrNMfP/HJGm5NnTK3matDGwJPzWmjtwF4igzspN3jNOrczgZI0P510bz1XN9U
+dmSVxUMa49JTymb+PqF39/DphqKgBMX+bAwJqGTcWvX71vPxEHnphFdBuN8SLc09N1B944PyLvg
7QJHb6dAKXPqf5m29zCREsncXmKb65gmslzHbDeZUChg1r95HELu+5mVpO9lrI0bVHjndivaS7sC
Mn/oubWHdDma6YaKmvWjt8wK4AYYEBdnm8c+zIGcITfO2F9YD/YaEzo0Ll1jyldhn3X5uTIk7nNb
wE+zGwvBALbg3d8d7HDdSKnSpqmi03txreRufOYhs7djJXGHP6wEs7KRkcszVi3N/CX2V78H/0nB
UXxyPpItUT65TVwiWPoGcP0sRS+HD/EuhbYChQpetOgn/Ysof9sSGGtz0RGaCxg6omRerFNdb+UR
2jkykEQe4KTenEHwMKVefdnp7e/TPMYw70N4SYWnNO1sCpbcQQqMcsd3jqjeO/1d/dJyJY6OrmwM
dKYWgbM6tjle5KEBonUSHjKmw6nT4yNMt3Hs1cFEe8RKRTPR/oWzLPgKIc3ItcpuXNpeblwIffSA
+V7mm6n+ygj6+ouJRzVa6G6/Yh9tGOJYkIgfKRN0FlkbcbeRH5fwD8HOYpv2+uKNKLcteTue6YdD
sd/Ab8zppND2n+7HkUgQGAfIfJ+WAohbkY82y8UAhYH6rw+XctFhJmA7YL365n16xebzh+9hkMhJ
SmH6zFcUfQ22QCGhuaOFY3RxH0a397cnr1xGZsS/JRmc0VW1WBaxyWiAJGc+XcYoU39BvBeF8U4G
gpdX2kR/nPmRcOQ4PSX0FVhV9ylNg3ZFfRLHRzi6KbOjYM/IAW1xxFJjVB/2jJXUwpLd0Qg7duxz
uF+c3wcbisTWx0V8tyJx7lU/HyfASDj2Yk6gbluTdCd+0taqeV1yvz+Jx4kqSFSadACEMqvWQBqv
AAn6ohZRfaY5Mof3gJOtKcevtOUDiyJgxw+Dp/vy3sXwx+7jYFpKk5SgKe3yssg+CgBKY5ZVOMSH
+ZsJ2aCvBsu5BHnhnxqYbEWLiOpi9wDXQKig/VU3mffjmggIJRYEFEtCOhbwpYX4B6mJtZrQIClZ
eQbU18wwPNoT8AgoCndpfLBdp+9lymolNMnxnpHF45fbVxAc2yQenuOgitlop7+8TBwsNQd1hia7
g09muC98UwL3M238l/0NC4yKsj9PepWUX08OkY0AIzuzDs9GREslJRJALPQiff7FAbgogMaag4o+
3ivmRhblRdgkEjqrnzkIK1Hi6VXqxV0LxaMpw9AwE9AQPWGzolz+N86mT23+AbpY7vEmEvqtPov3
3OyOFH0L+X/FVHoCMsHIFoenRYQ7WYyr5VfCakOrMHYud1Rbj8+HctU6I4l5sanVw3xPnNjM+buT
I8Iy3QzN3t2FCdx1F/PxTsOz2r8rLW245BF3fgxDksaWhqe+FhSVAGqs52i+WMg0TxYJxQHSm3Zk
LE/EXjLQJYdc2L5KiS3dpux9yHxK7e+ur0JlkZofcJ313DAErd9x2/6CFTySDBQ0BmHIEE9m5mDQ
Nec7UQTuWoCzGc1vzGKAww4xwH24Dax/fsofj3ceXe9DjeYrcEpv5hIFyGAUQzteL+qq0jnixgkB
KmrcTqn/Y6rNGZ2djq+/UVGrBATQDnMo5hqj06Bu80YIdGqNULlwV1HK4qTpalMaOHnou6pFoRS+
NPGGOm7aNSgfNEH47lUfWbiVDaLm1lYMopOwwKqmVbtXQqCcGc1D88v+WGQDaYOoeT2AlLk3w3Gy
C+ZYhYjCc49yU1uCyovkDkAAyNnVS+n0Bf39m5R6htHMyfcELuI2seUCTvMYsafVL5v7au2ubUa2
AaU0vMKQEIBC83HSnh5XvcwkHDPjdv0IjiQ8G9eGYAOtuXkSv2hmvWLqDQkfufB+6Ox0sZ7Cejt6
Csl+IVIttgMji3IEm/T1XPViSSoG99hCyy4g7HWKQbrRez8yNJo+8ZhR+N14NLY9MFX1W96lMD7c
7K2NVuAOE15KHO8up3nynvyy0zV3+rE6NjhKUJX5JbsMFasMtF8cfm3bMm0oKSj+C4f/sWwMmUSO
d+gB4AV3/Ynw/mcygAndjYzjlrhukFnxuu8PWjMszy2hWU9FRjwEdtCRIWQADaCKaZDOmPP4zANl
pPXuZ46p6Kwe1XW2R9xZMYXYxiw/GAzXdOCY0JipPSVZvQXCyIAbGhFqNk6RQHuNIjitfntcZTnH
/Gyq0DCDAB9QKZKOHqpg0v8al1G59ucu5lNIwuDNNAV5s15Epb4uEN3ZRPQcfeCLRpooLzYCxwf2
DwqVmkdOJXW6TjKQ0eBowqP84cds0YItRJsEIE/KobGgxhhzMF5Va/T7LH2mGK/pjGBIQTP6JZcK
R3PeI9cBh8jAOdBPU6p04+qKyK7CktMl4a7uhGYysPTko+JE7/ZfQeimQ4/nMKd7udUPm5tDxX6+
dbJjiYxNyntCbcwFNFf45h0JFYQx70d4RNLJwOhQi34DfoW+3b5KzKyDYoZyiC81ZbLoaAAKCidT
tzbMfew2WToPV05Q2UGO2YBPY2TThy0xA8s0aZqANyqXjyJJR2N+CSfprp8CrOtObiHf1WmPM+TV
C6wK3+GriLCNya15r67OggukqYTzUzQYcMUO+mYCm8daMvEfOkZ/tCYQtKTyD4Tn11I9FuZ2IfV9
ZBf9SjDbv0MJrjiPOEX/NdScrWwz6ugkO5oBm3bLPFbmoC3QliXASlipBWuEgKJilfXY4ncXc2MP
s7MAeOZJHFClbn1mHihF+N8dYiKgVwN4nbqDmzV7gwCrFcTN/zHpNksQDLIOJiK8MG5KZxBwBbar
8jzHMM7mOZV6YP4OyceR+zAfOemoFOxCIvjqFvS1FcM6DERL4bp52aG6Chqeizd7QFgDTrMY0WiG
tV2mGeqOrjc+Biexs6BimvMnOHMx8xLaQC8IVHwRXelxmCOEmAW8IMXkoVjZnvrCGWoc9T/s1ReU
JuW62gEvSjrOYfAvHVlpnUG6pitl+QmiEDKvd3XAYhY4jnCqZmHaEQPYTmBGlb9aVckgxM7GLqFY
13JjZiLRWD+XPZ51TtAyDEPly6YGnSH0D9HwSp5wRgjMZJ7HF95oBo0GkAxw5KlhOY246CdMzvJ9
Cp1fj4lTqyJxg8jtwRBdbpiT0c+TafTdcvbpRmBBUkX3Pm1n0wrJ/tFCVECHzIr9nrx8LuY0ZJke
u2w/CjVmS24MOaoqdLmca9cEuRo7A+bGnygBOZqqAMGVsE7j0pTpcrUiwJTjJh9MOxcVBXEwoGCz
0Zxns9fX8pQxMSjlzri9K1paBTzxCmY5uy9VPVZBU3ZErL9Pg9pKIyqJ6g49LBF02kpgwe2+m7tU
Bx7ycuPsEqp/Ah1RWZ/PApPsjGAsTMp2mrq1tOq7uURJFxWTiUkAWH8YANgnv6PMk+988QSAwi2M
oxcR2rIgec4zE3KAJKJZghDAvu0MF+Z1SQ8DuWykbW22kHAcauexk17vwBaV/cr1QJU3xuC/iNBN
H571td/rAPCfbIR8LGfsKOgad2CsT6BLskxoayeSE5bwxgNcshF6q9J5Iw6WM0KvgrkkGthduZax
xL/K0P51FMIW/r1NkCnaKTFWLB+lEZZ8NdzMXoWBra4gVaDtJ52uOf7ccx+W0RcP0DmtMy10Ppju
ORctWnQmAYoYyuaX99ZuJTbS3XGn5aiOYc8xpFVjWYFXzNVdfuCyt0UUvraZLeubGzVrDKN1i+Wx
iciTpLLjGs1Z01rGQ0aNVluoiGFUCCUKqkARILNCl6Wvu9jCoiyd1RCBMGzuau9esfp1jlYX++BG
2EVP65nhEU0tlVTkQ2+m69StgZvNqDLMhIwnHhdWut+DDajTdBnkhMVxFSG7SHjYeV9l+OYWvwp6
BrkkrRuy59PkDlIXxUxR8JK0J5IDEsFK9IWKRESW8Ywa6gtaqM63B2KjWkUepaAM4hOYM2TinkK4
liStWFGPx8Fiq3HNQ57clLcgwvFIzXSX9Oj001BOkSXCggCtrxlfHbcmeChYZIjOPMhytkLXDhPM
jZcaapw+/vRrU1h+0ONBEt2nkxO/IhWyMR8PYgLdd7DNC29laZ4ix/O2R3sXjMW+W/+ULk4vWIPI
Yh05GTy/wpyGr/hrjXfam6aep7FPYMqCGtWupRAWK73Yx1rmZGSd196DWHhZCxju4MRDWH4opod0
75qTYHo/P3ijWZyEDiP9EUB//ElBIO49rLCMdbhPFV6wVYUkCoRIak/emfGOz+Cci2cLKvIqjMYz
EjsCWmkLMiEu4mGJuzi9wH4PFPs4fdm2sO+nlyn2ParV+rHy03xK4/8RAE4frhSG9y8ej0+RZk37
LHPW25kZ35w3FwiTXXrRVXiHUuIue3h7k57NjlKGd9Jhj6t85eND8RlW99MVCsEFcLfwTBzLH6iM
wvOlmheHAV6isy5yDTqs0XBKEOvlNDvpGB5Wly5S+OT7GX9ajVU/LGR95EF+58KyoKg7d3wpG4IA
JWnqIMKrTEqPeH/mnPQ3AQHJM1CrUGFDdMFt8Ennc/nqaNkVewfEq/zbT3MotFjV+3plb1Coxmo6
XpvPFu2kaB6nh7KL8zTNQhYwZA+5nOnoBGUS10rprfT8rEawfz/TrsBa+rsYPLXCfg2Oy0+X9gVf
SDVBJXbAKBtaChQkYZekQG0BY/r3P8jZrQIJH9DIpoRGYJtw4+ZT9F++v5wrKMx5hem3OzWraDLR
B+Hgya9oR5bCPV+5njiPjrvjY/M2ybyu18dgKiucIEzOdpkS+CnvuHbgXmJHdus1MefwGXFETjwN
Pz5/iqJNbZrJKWC5eGzakd6vT0ulJubQ1eM8V9qNigZLlAdaG8iiWPZikdjM3z0unP175teQbVUt
khnLveGjow6iJuDfci4Akq4BPkmEkg4NZQxJ8S7W2SYe4uymv+HMOt4yFEvlHI6Sy9/fdcQXGcBS
48Sx4iUnBj9QyDZoMTblFur5ED0OiyICyK6poL7ipnwTag0nP2/AM2KVYe/0WTrFh8K4QZan6hca
KuzaMn5ny2sPPOS20PkR3cwz0yddc7h88gyZ03CnOFsRyJA4kcJFuyirpkgRDaiUU6l9WpdZkGH1
DetU0hoXlZtTKXFutdEdaZz4v1+KziIiRIhG1nP945RKEcSgXHwauVf0Wkb9ZeTsgEyyO4Syklw0
VmZ3piNMTFjO04Rm+hj2bkNSJETB7Pb9F7vlCqmsLIq5h8I+3QkNaPUWzAtXmHZonCAE9tW+3/YJ
oqQUV8X7QGSuIpkIaulHJPQm7oKV/f07GHP1kjzoXzyuB8OaHtOhBgXtDhCaHVqWU5It7bIM8JWM
pwA/bvYEWEF6cD+rtTrS7j9rPxSfWmwx6qlKyww6jSrFbKU45+YW+rMQ5NT3w02/+PRNHxKbnBLW
fzG8LhlSdgJAzlLr15ZUT0YD2XtoMwToJkXQQt/tAKsfh/yjSGiJLGeoH+YwkpARG6k8rbYLQ08a
DY6BsHSsDJR5w4rgKh5yq1hqS10WKGHC+WhWiHgxgiNla0EEJUIPXkUchPZiNvXw0fbwxIDYwQhm
hNviKmYvAMAMOF3URcUiqmdl2Vf/bOXHAZMaLfo9+HZteSpOmy0I6dsNoNQO2BoBxcsKkuRroAuR
zjhUNBl/09WgC7Ij2S55wgBnCZJHzcaiki9BtORLOF7f5+lFPuL2fq9QGGLnw7Ec71JKnn1wKVGA
Ac3LGrp+/uazmQGDOHu8843im0sv4A4xygfMu6bcxJKUlwWusNgLQlaQOSoboCMSA2a0mIlYbFFj
hZpLBZq8Oqe5vnGy20MlK4DZg/uBMOnbeCCCL25S26u94ajnPuSd0VtkEtWNBpRemey/2BoXd6RZ
jKCdIkGBJzIDGDVj7Dz7Q/9YleGSDygSG92eNMHV9EnV8WJsi+DpLB3QJaBkuqcfkrXohdo3CXfi
3vstExpwsQA7buE4pn67jEPDXJEEqGhHfUppMgTgw6Va4hmo0BkisvWwJhTLxlVAO7uoKmfATaUR
jbTl9IDPkkGKC+nj9kT67ZOMmC7DMKbtVMNhnV2BMKra99In4BHmCdBhEz0GRbn2ridRyogP3NFS
D7de+UgGcn7yVJ7TMBaNvqi2c1+YIixiJ4oN2QmZzSXpLtI++hMjiWcFo/Q1/pXR0Re852RJKuQT
Ru5hHM+RpfOmx0H2fWUixvlkAlLQfHccyGpTvD6ISZbOR2MjDKMIq3HXwPOI3JsnhX5NrnDuJP6x
DJ2jVsgzpNlwvgYLnoR9xaNG4Cp9I8M26nyrM0XoR3VGfPl1UdsgnqyGiYpaM8YrDnky7q81PyTD
VdCCMlxuauCGNfXSUB4f3+hzIXtuDZ0j9W9/kjNnFvtxJURluoU3eMY2i38K3vxwxRa+7ofpC+f+
Z8KlTj7eAXEWe57u+YAE2w9gXtvmH27NLYjLEy1EVToMXqmqi6I2oeFPlv9pOM7JYAxpeCFts2+T
JkEKG9XDyL4r6CpoVqVZoFRCKyvtaKV6oU8XzN8OTHVff9IAuOnrb6pXatjC2/bKFnidJr+dJdYK
bfKSi9myiZqUZU5sJbez/NG5cx+4SPP+/d+hqjt8t0fMDhedjqPGUFRSh5tJaRtUDF4wu+9+03aK
B4Y5tkF63JBPhgLfCXAnn07A+fNzuNboFRYhXvk//BEv4lCZiAD7AUnL9a+Iqo6RxAd/RWucyowy
0X+I/UAdwPK4kGjOPYoDBkQJJQG0WkRh3mQadqDnuXiPGernN8UiT83iR1loO0FS4jKEsfWM8qBq
zrQogWP/Te3HnAcBgwdmrELjmmqDY6TMgnRK1EQ7wO8CBpTf5w8MpIRkkKIKVQQK8Yo8e85aFV2I
tsemkqWhWk5yF7SAqMsbPaUn/7jL+UaK16lGGqbTXC3bt3ja+srDnAyyb8ocFt9E2aOjIfHAsR4U
zA4CGO37/BnTsp1FwN5ZfssE87232642ZK9MRyPyzAQYhJJJuRuc4ATfsi25bSzvQrFHL6Vso2hb
70/N1g8KiMfC+j+nm1NmWPNQ9ZR3N0Y5CWo8f46u8E8F3IIfBMclxVFOHzSpn3gt4oy+siKN/M0k
QAa+a2tThkXTqHf4GrxvKQQEO6AMR4lPJAbNfEfHEKNdDgQ8l8mhIgRZE8eUj4FQYvhk/H4I5R7E
Mm6MPLxQX/BE/L3z3s22PZov37txaNeo0+uJD7QG+k4dpEXuf8RTg3Q3ny1ZaqEporIxUTySQXaw
GofM8Hzqkk2d/tstr/cuVn9o3Jbm7Mp3vPvqsdB3HnmALqvJf4b/T470N2exgTH8sg9jIVe1k9rY
q0xoAiIYwSRHsSNR4LhsvqXxBqdpUCVkAydwOQd5nzeZENS1nZuItzsq1haqvck8NylbLHi9JW1v
/lKirth41gm0fxxFWJVrGdA3HKWW4jm8BCwZd0DOYE/9LQrBwqf2+tmG3FaVgi48BxVfn7lX3wJt
QkbJLbRBSi5PIn/fqP3RWNqwTkccDYrtn9awC/hDQl6WALk4GcEdu7sRWdEi8eqGWntpcddDGsm+
s56ZrgE+mynq0SikGbi2Q7Af7Sm2CJvV5gpjFYcQZJHwwXMukFXmiYvBq+YW9sGdv16Qjsl4Q3BI
jtZVzOuw+egBPA/HNZSwUN3sgy5tVZsSi/XTyR97+MGjEE0/Wj6fureMY22PNyBjxdj1g2cHC3md
d2zwnwmae3V4sY7TEaz1WGtg843wyivbwbDqiFd4m5s+NrS9NyxDzlatDatRbx4GjJuTPvGGXIRr
8nEVsbvuyvqTsLTU+jFXm8NRLGDTsEHryh1lMSnr2ElIzcVrw7/PNRADKm1pcDr5OlUrjB9Ky5Y1
/9GuwAdErkg/NEm5CYNMB5go1oArnnVSwHCboBEAcCZF07WT0xkjl2+nrd4oLNDFicTgI2UVLl+J
Rx+2eWeuDfgOkiARkoIrkl0FTyTnUNqRPFhDawVDluzpWO0BtN6jzgqHYFDKp7y23lt68ypS9Vuo
F+tnOyw/V+JHpfdjRL49HnSUIYTFtya9cO/Hng64aPWKVbkqREWv5XI9LR6+8YlQ+7VUf+44B9Fo
gIIQLigdunDshQQIJtNeeE6fX9M9+1zU4UkZ2j4FrDuduC+MygrezY4UA9kzI2yffhJu+mvnCrFI
WdsrpWpnau9Q6E+N6AqhtNiKT2xfVnmnFzDL2iaqwGSURouF5YX1sBCVBOAuiAgRjpIVNOvC4wKO
efuAYJHo8oHAOgLnJZu3TqjTJinJFhWY1xfpK2rFJNReh8pR/K7CS3aVvStw6WudSZgUlilQx5Pl
EGpOx9teIltb1i631NSwnWc9kX9fYa2hs0xVaV2yBzZzxN1wW47MizbxJT0XMGFnbLda/kQNEoTc
DNnsP0bvNOrd7z0C9JvlkG2iRxBt7LjKxvTp9dQKumbd1PRgfAsAHDepNrShvReEY+0bEhWxyrl/
n7i4R0VimjUhMwax6rivc/G2+tD02z/rd13cKoaqCMRC60AuGNuUzgZ3jTYsU/BPAYiIh2kNAyb7
az3KyvrrlqN1thrSF9kfKhzFGpkv7+025R6SGdgKGw+V6jVr44j9xkV1I2PQQU5U+OjTE9yLp2IL
jFtgwsnoliGjg6M3mX6juOYEqZaueIfbkcGEEa8t2GmudB7IGqVIOAQPrv31yYryM9YTz3JeaQUy
X+6KOjdiSqR21tDSkV9wcr31g64JEqbIDsYBtMlZPV3gmUufbkHZpUmcreyIvtoWG9uuFhgFdVeN
w2DyyA4j6QZpBlHNWlSay9ZC3AIcPgTGQrwunllbJJptQvxhzIxul42GdmV1yIgR5zMBfNrB80HB
uIapvvqTiDBTUyL2zgE5QUEXTJ37AwhoNhu6Z+bZPqRfQWfXL+3vowDrU/QrpFNuAWXFVOKxMnun
HFcLhxERXhsNOShLuA7pf1hPU9WjjXWEj8Jh9NXx2+ELgX6zeTKhYUz1thIa4uN0efpk7p6+0hEY
50xJARNfpP+iQRPQU2M5x/prIu+Rc+ilG+X9v8vehcEHDdXExyxEq/Dfv9EVHyaG76o184Voxy2p
aFNER0sq/fYIfZTCMB65OHLan/Lu54DY+CI8aAvpVwCiXsANT8tqD4y6I+VXsJkLWd+tzSx8Vos1
TRYMQXSeaZ1TsoaDNX0yzFpG1vBuucU7MBxomFqpp/UlSiBmDLIpIORVDp0ihjSyiVAkJBXHPupP
v5FO4LcSGPQbCYGOu+8zA+qeix89miSngF3RyBofz76iyHgyq/8FCuHUus1bgoQUjXHha/t3F7CU
ClZpuSrFG8ZGgEmpHHXDzhaZ4grZsx/GGEzQkbnYu4wXrcXuYpkyf13WYv8byVetU8JfcaSuX2cJ
1DKMg3pu5JXOFubWd9ONmln7xYuiR9gQN0gUNJBJJsG8nwmhIDdS1tR1VDkWgwNSZJQaUkWq6iRP
D5Obfi/Nh4EiDNmQnt1NpYNwpDwBsKtyC98OVwLbcAdX4EY2U7FmPIL1CPk5cpRLQx73tx+7i91a
qGLZRBxYxcFsEFZjvEB+j18cFtJN8OfsDbuxxXXUasVvcsklpgfB79nkgWbjh2mQIKMJDTEU5q1q
UnXtoyQG3YoABt8EfAyRKZMRLTp1j7fRE6IWBmJ1WHlqgPdMPpXrL5BAOGQ3UdKeEtX+tglmuatw
xD8dIn6IcKul1/jGx8o+4Wc7QVNb38jFMWCJcMEH/l9kP2b+Bb1mgBNkksllhHqjtTi1naOoXrZr
W94m2JzEOH9Zy87MCYKx14CAMcWeytYekUjs4UG8d7uKj7dcHjPNPcNWKMXc5p8a58WYEftwXJku
RExM8X5Ad0+Rb5ayzoMlNAjgf7BvufXXMuADrKsmjW8RF42sL/O8huUMOSrzbJG64AZL8C7t1Z0C
vUyLaowyNMBzY10ku5t/Lx6p1fajTgkXrJ5TxkUopawZXmBlzqS/2FANNUjIltZCQ5VKwJ5CHpc5
rWAZETIZiZigv9YuuhCS2Z3S5FlXjSLxfaENsKedUyz0jv9HCZweop+AjjOQoFgdO/8acEk1SPmd
GSmFsEwEN4G1v26YfyLjyD42Nas2KvT/j9QDpSoR18INUC/ghW0NSuz5qPR/7ZN/5OX6ZqxvpCkv
tzD+47JfGaaJyFXJje6dNWa6q7ggrVmba3PZyf88Gk/UoIK+VNfEknUG0KQBn9qLinNf/WPJwyDX
dK+StDW/qNVaPCN+SIAFr5TzAmjQHbOMkmFyTvabNCYDRjoUCAbdQNLt2jC51GBxkqDEQ4RIQJvT
/9I1k77HiBoQi9JQPnyk9nM4/frfhmo1OHeSAHWlXSCf3GfS3gzehw3qR8BgluVHtgNuPn+ESFUn
3Xlr5C1lt3WrtV8C7ro31Q20TGeu/nW9UxzFNjNOqdAj5yN8TJMgmJXCT3cm9dpVvtgSU1v0KVPz
ZjtbMVyA+OmYt8moGfpJByifvasn3LQB7wsKBPuwmvJ+lQthfRI8D4O3mqqKdPjganhqFK4Y/3cb
D9WTsNgnfnMFLJltwkodzhPYiYGiarRm00DGjxnN1/5g1eLwlEmqtXhLgfPLjlcU8k2VO1OpdDeV
uM4SF+1slr/O0ONNL1NRT5H0n4WxQslq+qDFk55jrjNEPQN67UJmoCivFHlWlqrElMPAInXc+Ga2
8/zv2GBM71ZIO21BExxp519tq/iIXk3R7JYSRfXQmoetSZUVythlNd8intnlUfWOSP8pJhTqVrUM
KZaTPW8+vyi7oIKYFTBVCpHGtRj5Vr2iq6vxOUruDEzv+6F3uje37ifxI5qKVtKz0YA/hDYJG8Ei
yFJBVeWJBWRS/NPBdIUnsyPFpT9frFZOySq1Eo/EKl79UupixWLtd6sVJ1cbJ5qN8knf7Aj5nRH2
IY8law5JcHRx6B6zTdxAfxjZLdRQZ70+6xIs7UvHxqlKVnCXWJ94DVguw/DWrTjq6Ov82m3rLDCV
SaJLG1pwPdouTxdnHBq97XvDZvVbyaR195qHO95d1CAg9rljipicPeKW4MHNYB9iAbietBT1oH3J
J+vCT2Ndw/7CYqs5W2AVlOG18JkjwivhKKty3T416oN3XamrzDvC+DS/yLfQuutuaDPRincNowOz
dUq0BzYviC0kq1tnad1OiW1HqAGLhwh0EOXCvhUv9uS3TAwN59bN6+2iaeYpr9mzPQctPif9A+YI
gJMAC8ag2d+9gJuITIxF+Ng0rDv11NDwNh50FLD/5q7gY3Um1JeJZ7uqENlgSRhx6HmyV4aqLCDf
CdKKOYfV8wZyz8+WFQR82CcLbZbERJmC5Dz819jhyNamTK3U7kIhjX3UbDlms2C2hU6mrTH4bA6I
I4cjyP20XrZlrt0YJvujGx81b6Uz3xWeoQ/RgM4gu8dOCnx6vXk6EuJXX4FTxEvRSTr2tCrh4eY9
rJ2tU3DXitH51sttGynzlSNmoBRHbAkC1Gwxw09T+6TSe0cXViNvx9igrHeC4IJae/uZvv5OoUqJ
0xkWJ1dRVSADXwRVNrt7+ay2bAQLSTIls76XvykHqC5deeOGloOeWdf08nme5Cw5aRzpwmFs8U2o
9omnC159ECKjkbZEEy6T8bYfTsVP74fh8ScxO1n7xdvKls0PQx60RUdV1sGzGBbMQgAYNRf7cNk3
6j5yDCRZ2gYx1pliBtuZQeBZiUuZrIIB7gsAoLKIWHgh/T7PjABKqMdZKHmz1hkz2U7atOaw3EI5
l2dc9AFvoPfqK0ZkPft2x8+gdRAnm757noR9Na4cywgG0F9D9srl+ZUGYTqTXmCZBKVPbPKRqPVm
75lbfVnCseNqTGu2lRa2BWZTekE8W1MKmJaiIIZf5nVBwOTvTB4pWVWg4j0CoC1Y3gxGWxBaGRDP
5seYuM4XI6I2q5MyPbdVbfZTlnIYJjI6ARXhywUf6CDz8jHY6mpKKaPL3dJuRNpkgTMNFO2CDN/L
pj5xmiZMg/xx+FimAD11N25IofPt/omWjsNjitqVw7VIBVHnlgB9H5/xVzqf4iK/q7sdYFS5oLnF
SWym+vnPiofxBB+YQ+Eep+E6pA7ZhRqBu+DZT5Hv1X/WGy2sB9K/0Mt+8RvgXaW4uqh7XBptOQMk
y+tZ10yKhKdlwAAXBp3/5l/6OuZTz+gNrXipGlvBj5NuoRKX0/Jafr5TJCn77W2kF/Wjxs2do8Re
ndYgpQx4Cl5k1WfwoulFm02EilQbtoGArr7YhhKWdewg186RJW3cbH48L5tia2fAoh9vJeCKztRR
x2IWGZXJhKajFlKvwTxfEMh9ifFEy0RQ9o3jtRe9LdfJ0en00fSGoQ/1bPx3T9Tp+cxOKToPJ9xA
R+WGXIBLcqRqa2wlJ/qzCq8zURjI44sajlVrtfNcldzfcmVUA3pRoCjl5N6dvyB+cQyPofAz4wx9
RQaCmZRO9CyCxEii/n5HvlSZu1nGVYyMkc8MO0rhL0wSLaYBD51ea/82z0eSWfbkiXnXi4f79F/a
j3RG3ulyFtmyiDmJwqlu9XFpORUlZbl6siee2MS2Cj2z2YSFgorp8OrzIVwqKvJ7pZmrFuSLswUW
P0xVu+tjSLyiwwPlKqCMw5puM0qS6Qmzpml1pKkBcccJx57RLp7CRqwsevgdPY6U7gIPM6NLCWB+
vwgMgRsmyXwZjGAIGASWYNc2iZn0ZQA0rIMVy5VZ/OgAnl/GA/D2p+aISozeBHNU1OYKzJYIM7FO
BwQnwpuf+2Tvx9/a7b52o6B6fHi6Tm2KzQbiFbYmxB99N0zCz8cdDPCUjSa1hynafBN8VTAmmAL/
yP9fC3f/PAXAlh8sjL7sMKufGK1FyaFhMQjGmAkN1S8Yq3tAfxxbbeJ9HxHId/sffPTOF/m8RMkL
cMV7vBrbVPJax/cZSF/hb8GaDxhaeSKL9oNSFi0dUtUrgwYjKC2h2LQz463yGOiaJsWK3f4Nf8Tv
XWn9nCEo2IY++vuwgYKuaEpNQWwSAvLqVcMN5b8KjJY+39ww2ZhuCDEljM3/uShmHbeFN7Tm/oJ9
73n8cWStcFg+t3PFLw51fi39t2aenh2FTCtprmpXUYoVIy1P8LkGbjpnWGsUd7ikOVVdx+PAMYrx
RZ68L0rX66+wlm1P8SGPy9kDewgM0DfMJEGJ+BLzrcUnQCCvBh9DV8/qe0f3HvQ6CgLJRRRU0n5v
cdqJiSjcKT7MnxjfH11V4l0iUWCS5ds0ELAhzakabZM8If7OYApjDaCs9JiZItxtMqcyhqfykW+F
ff5KChdoXh6ykIQIZDNpluN9/el4PyAii0IQART1dryJEMSkeWddZ08FVVF2UjWZa8X+jCA7jiUp
sDVc2D7VwcxlS1fh19ZSLG8K/FYxT+7hMxpZzjH+FmTewPR8VZjd2SN/hn1P4/FjgwxPJKNmAm80
FsbBSU1uWdGqHHLDUJsFqJt+pklNUqWHAboCnBlLdYoo3ei5LIfiMFIWi1iaSConaeAW4YHy8C9D
q41nurH+UwTzHcEiL8Ik/fOlZkf7bPYHwsALzomtXCBHWvlOzQ/qQ+muHcEY1FKDATXiIZs8nlGO
rYSKQb3sBNLyHFrk0XJkTLQuNhbxdDxnnzbuM8TQtyPJaK7bFfTMSmASr/DWov+cXJpjM2xEu3CR
1KOXSOAR1G7el4PGmcgkvy5eH4ByIwsGy2+CJg6MXoQcy+4UcAV7QLsYo0FrLxYFAlbTZ6N1w6zG
ArjiTTP+i07EkgxyCW4+vnfU6m7TgLDpypgSAt0JZngV79fDfeHMVydPcvNm5DorYe8LTIEy2YyT
UndC0veRG8gKY3Q5/xFDhRmHe/DrjlXOvWgQydFF6LwL0hZiJV4799Qdsr2iFXPyCFqaEB9LQKdh
ygBu6BzKLlvSOspZFhUKTnRM8E11bEfIEoZ6aMsKTjR/DoNBtnQtq1+hmpcU6ZoDfxF1p69yCFVg
03oLnv8nifcxmYSxEsNYfFWGwoyYp74pD/4J1Ik9mt0xAAaJ8y4xQCGLkR5pcSFeaIQ8JoWPkS0t
/2Gn8hpiFgMRWgDpP1xXLyY8o06P3f6L3AuTB3xQ3o0uUYD8g6m+eANb8d9Ebdwj18ZDOLOlr0nP
haIqhPcVKZCi0lhYtwwwfk9NhA7JsITEoPW/DLEDZs28qlXXUFMlbfbX8rqmnDaI99ckFkVLdQOz
RP/bsh/yK6Ts1FosvHerXX+h18zLsg9fOnGAtWOU4iiENuFvhDMR3mJ00V54fDkeShCZQy+GKZDv
g7I265C+mKpzZv1lEw75m/bLwjYJEp1qrt02f6uj4vZCINtfqeHTHqDFmtPQeGVCE95/guNpHBWn
d7M/cdJ1FEsMssjKVnTPluZ6DPiOI7BeP4XsrNleEEL2/Isq8AOHTPbOirCgnDcmfekF0r3AKWwd
M4/Mjto2i7b3gCGzR32lzVPPsc8qxH0X5QZtATy++o4x+1wEMjfMi/L7/CebUtPwwWDy07QGPlDi
lx6Rtb/cFqGZ7ecv74j5GVIYhCwAESGEdkTQOCnmi6WNQ4wxgVYjTGd6grzTOAMHI6c/yyS6N00s
oI+S6O8Fmw2nNag0V+AiK4uHf37zgK7KNy5HKeC+x6VHdhnEnB8gdpdB1c7elAi1Gb/aqqApGL7t
h/gstek5NqGU8Rkl+qtrW/rPxCvaX2zcM0wBMWLJCucwITXUnkD7bmj00jlR4YkKYJLXVJC/eQ3G
gGXXarJiBK1NdjQ59QRkhkZN7f6HAojwRj0puiaDSFEOG2y1fB/FhLTwOjI/cGCfT7FuNhDfZ05h
NpW+RBgPyc6m0WAUpEXwyMDzXYGgHvUdtTXKqRzAc7CnKz6uFkDoQq0C9sGBR5heJxCAtj+G3W22
bXj2cX6NMuCuuEvFTPyeE7QJ/B5LXFyX59cF0DRKo84ik+TQGKSdBhnRdBo59XtBfq/01mYoDuKb
Bq5Znnse3b47ERQu10XKyh1Bh7GRYmMntwdSeFenaFpWbdd2MMxW13UoYYVH6kXQAY7G47aQ8o4X
1GpoX/VcU0ENiUN3yzkg9fezaEVyLkj2uxM7jqdDQXnx4/KhuLLxbM15+41rCjxTuqr70VT/bbV9
D90UxW0u2TgpnvVW/0XnXnjAoGn+UFcTZOVB/puKfT9NdYFTCD3Gf+DYOhhRvyD1evkmzS2HeHIa
U3W2JIuj1/hi8m0BS+3nPH5U7o1YEw4xvzqCzVO3jCRcet+o/ugHg30hCysu9iiFTAcCQbp6l42f
AE27RtBuBHK2JPwp0Iqp26DtLOgE6+KTKW+UZiFXIxetRVcml1zTtD03W8ALqJa3l6m/Gusybs99
yrjrPb1vMTb8PK7PwknJxiJLWx+Cl7Q8QYisW9R5MhHEEK3TYgI4UDmqbYW+AmphR4cPcWJN8cOk
MlvdsDUs+Fw+/oFgA62SKSqZd+zwYlcsKbyk9V4xoLxG4etc0FkANJaOxukq/lvHg2ohxCBU4jvB
fVbDfraPqS91zWeknhTt5DxBqJWhLibPVTKUYdFcw9zlqzFSxUx+Pv8cEt1E8tWBs5dgxTH2HH+h
yWfD+Jmh8ooh/sAn3lQRvQcUbreTjkZQNtnIOWm3qFr+MbEz2w1J+ybz/7ytIh7Ee8PTK5xHTol9
9nmNb1IoYxGJJfB4d+Rn9aj13CpSzPz6Wyr2lZ6w6ZZT7DcleNc6Mi8dXnMs0bbFzMPshqBJnikU
RtZWkADUcMWsD5yosOhFQDktEwNT9gBAJd8qiIVm0S5pqYtJpLWyUvX84NS7Pyd8vXBw49XZJq9A
RZGrkPOG/61WpjbzyUG+8ozNWcGUSaxxhbUiB5Nw2D0IgVnAPTZnFDtCSv1n0gA3fuM/FxmR1HEH
Y6YYVvD2kzQkA3DsxZoBwAAsaWKmDYUzT2i/iLvEbWwwnBcWu7BW5ldS53VnsAH9NyOs1cAZLWT2
07wrHJa3bpNoPGH+39ZJ4uHf6n+2FYlh6LW+2dkNTZrPrl1mfoi86VTXj9KEjP/Bp4ABZpz7Z5tw
TK/FZAagSAUVDcIpxL4Ro6jKPXlqyG6Tl61GFeiOEtmcZkpf7oN+HAMG8e03XMvPupaF9WY5gw4i
cI7a0NN8Rxf9+B7u8afUS4FllwMcY2eapEIUtPyzN/YGfmLDB7Gw+f9mgNeFBvTkfZ76YxmrrrJD
fRU4aGNWWbjsGautjm9ZB5CRt7WKs8fjXZJHeJnMairFRF610B5i2VV9BJEMHIBvv2FDVhjBjzcL
1NS9tamKYXWjlybRIl/nOayjO+Elz+i5ZSX3ijvy3rjlK3DJaee1bZwlmcUGk0rgkvhMgsVJaoB1
E9hmv8m9V1+tduw/E4wrsCdKj+BG+rV7bRNYbg7mlcu5/NBK0zEDRJg8MTxTKv1LqOV9Ij+Mrw1b
rXcsoFagB/lrRIhrho5TZs8fARaMNb+/m5Z+zTAwaokJqufzsO/AWVDea91e4Kaf9lQv+63YCZ7g
optmeMA0aqnVbZoZYkEQoP2Ndul/vjQYnEq5d543oW0AHRDJRfhf+FbSMDt+uJ2yFXCtqwTGAKLU
2rzRn+pLZbVTTagWhYg91NWuo15ylVbWJYqgzxlwiwz04v4mnritB6Au6Fg/Shdba94rQPtaVXvN
rHvXlaWOTTL9CTHdhUUP6qEAhYPFuElKxMrA9C6qeDncZm6a0LQAtAs5zn5kaAnftBwp2q2rJEx/
Zk9CRZRPV/xndC4aN4SqTdBAwYgTSMxyEaTP2cIO/skOl1LPGKuJWBnGcnvgf9X+6WAwRPSBiLS7
HrocQLQSaPFuGVdgzmdBj5jv1LbV0s1XbGkJlFMZiVLl9olTcXb73HcUnGG5VFGvnBb/9jf11ziM
4C7dvm+rsgSeAKAHrR0ccxdEWUba5jhy4WGS35iWg4jdTOGouhwEvejgx629gJrERycWQVRTPL2N
SujAd23Xl+U3hK5xV6FO5SUxMS4n/iNCkyokoRdJxmp/AJuAkeahMzV8Icnb05M1ZcGlexiFVNUO
ShJiBkKGJEP2OyR8yGIkbt+5CvUqF8HhSzSppn1DzCsx4r5seLdBOXM/X61RRgMqrWbYn6hLLK3r
NCFGX6QnB44WgwWkkyV3otVwaW5aPzDbEK78n0CWCgXWM8G+qqAbs6ou3hsxRetTBzqyDZPnNXt0
yBr3erFgAwNjFQbV+Qn6H8vUyEA+01lYxjKrnqlB4m5PhkrUfYljQnwKzXWFhLI6JMg7PZ3pzgwo
qeWjRUs6Tst4u2RWHkHI4M786z1qYgUSU9282FHB9Bq0YFrxEe7QI2wv0wxar7ZFSUbetHJ2/VAZ
pMWO35sg0Tgmpl60FAxRz4zayM/o9vG3ckO8ROynKOWfPGzxVdcriWiJADhdiINR3HsFmxCG/Alv
W2fTsAVIw5O0DG66170vBkMozbst5tJIAXelUAYecQ8jremmOI+/YKsvcEkkW42uaO2uCvyhh9pP
YSoR7l6O6muy6seSlgidBrb7xnZ/IcI95QI9rxuR1O4eusyrU39IZoC8a/LlagTmiuK7ruMkTsk1
Vgy9l1I7CIORNKvXVqdtp7YTLnpagJqxnH949LzWBzj4OHloWdIy3wIZS/ztW6fNu+Pz9NvsyCsd
QA9jrMh1jTK42FoFi+SkU40vI4it2LCWr2S0106o8uXph30ONRuCOiGWJHVIn7ZXqqHwCuYYgBrm
hFPAlt7w7I6prPJLLlWatcmf4cD7lKg3q72woETZmPfZaTzFcBJQSp3WCHXJGs9nJmMGY5VKjSe+
gZmK5dHaXj5XfJNVIxCUExdo+2NoAWVViy/8PwZTuvKXYDN2WHeDdnDSdjZP5j66wNUXzLExNCfa
GFscVZ28GSKPq6/9ho8dhtjmIkKbhvbjZi13YoNUTXZrJ+IlUmgOQCC4F3N47/xewEsyBh4FrHkH
vRzzdb3n8SoPeVyvS25X/kcL3qB8i2qvUdfE9pWCJDXtswrpW7iADXggETMgxNkBOa23ZvO8+0wr
ZiFBVPOcaeMVqz5ctRtCoUN5ngWNdK2LZWqA5XIJ5kkpxEPyHnJPtE9KhUlBPWJnN/C4RO9ax3N1
8OUuy1BY/jINQxQ0OWJ6kKn8Qd3XaI8KGZ80QfbDlbY/64HaL5qQkLURbiUFTxbN2NWu3WK4994F
zUlltyBLQsFAVQKel/RnM2ezCpo9vXVF4+8K06oaZGhHZ6gHlKwoNW/ThXOdmzMb/Zd6yfqjFQ+h
O7+Pfe+j9drWQnf6BPynmXhP6YAjzKpEOAnsaTmbNTpbDQ4s03u7RuP8dDu03TVTyWLLOW12dj0q
Q3tPrLG2NKOB/JQHEsCCyZNATXgIsLbT7DGmxvcnVkjmoX8eDlrnQ7Bco3NthJh0UB78w6Tn0mjj
8k5aQyvC7c5VYAchQe6/axtRsZ3Px7umB72Nj25NUjZ0MCj6WFgUJ2n3cfEzx3dxyONMaDrA47Hc
DWtXzmj7ASXacmYu2jL4DXUdi0yx2J+mjS513xHt0RN7CWBFzgIKXIthMoJj0CdkB5nOptC8xCRX
sK+ydjB1cV96L6BtxnOVsDA9ycDUjdxelq4kDSg4LXXxv/zGOPaj0bV+NmT78QgpCrKvNVxZ81+Q
ZF8QexkNKb2KBqwqUtgIhN3068mR+PNeVMLG8Z33zYjenBcHSVxwxVAnqLMhFQ+NjVLbHD8sTSEd
zvQmzsfzPuDYu8andcje/cky5A4Zo7npkHnLgbdPlLlxJoT0grGB676zdmgnwbMUvMgrGYY4TlqZ
v0LFptijI2xFCeJI4mgA/lHqyEZZW1BvQr5AnUZdtt5FSCHQSgEzkuDf/GeWe3kbpJBh7qt9eU8/
wv2dIuDnmkAi9uUMhQ5juQJ9YvI6pHQzQuiJceGoC/dF7Nhg8ndU0D9Vv/co8EP8bMScrnLAIjqs
BeOK4Nk5hN5TYvDXR2G7CosuZPI+yjBDTNOiU99m4UX7PVaHERB+AN8U1tYFed0eMb6hLChkjKt0
a95biRXKRaZMx4mRCs8sWqi0/Y1Zh8bAFabfoomLsdmB/eXi35d4H0ij88yRrzq9jfcc0HjlRKPH
JKN0jnBqwb5+CB7Ea+9StVeR4TFW4jkTYv1neRWfOHHGbTKeWo0xoRvjwFKHbBo95qmlZJ/JMba1
ofu3MtsJx6KI3BOQmvnLnBHi6+e4tdFNu/bGS+wSUgq5vM128dzp+TRRDM8hYeE2bzIKQRfbRcQR
yZXiKPNb1pjenHCBqhaPyRBLDzXj9LkMFYMaY9uicS49P/CqMX+gycbW8Lv8x6Sk+C2OT7XrcGM0
3M2IBMPwHefu7PApjOcs8Bt/bsODpbgDaQb3gDXYJ7uuoEqrNOERmJ1NVASnQLPH8h8BtEdQXkqx
NyxBAiZpStYJt8hAPX+jgakaSsQucxZVMI5hkPygbv7y1tQ7zfEW+Mcl5EiID2cp69ra/1Vd0svJ
h5MPd0Iaocwr46uhEFgMis46mrL6bkiVonKhqq63gYkRR1rfJ4vE82yVlnHHw25tsCzgNiECpZ69
ayVyjh0p6yvTUn8iLJOFQN2+ejdNl4H794dJbPjHV2+euc3sBmd67qUUcZ+5agbj2hZfIG2Fiuf4
jMO16o2RclSJmbYT3M523JXhBqh5oklk0CWj5Y7BozvEHx1OCxDkew5l6n5HW8YlvDQns9onETG1
fCBVu3AC2acf9lGFOFm0oxFY7YAFNVcHDX/97mARhvkWgaqr5KKbX/O4v0Dom47bIEnjKWU98eE6
rjN/s381cLzjb8PHzKmluozJzShgqsAFFr0jmyxP/kPfYe36aBeOLxpVyrGO7mIohn4dPnUMm9mX
9NwZ2muhA+qG8YI6O+foVBP4jIPbPu2AcVXUWmhB1NP1xQSxy6IR1epleciAyPQPrzAYnrsD9ntn
1vpAWv2HcywKwVZ0SpKUwOQLUnFBz1fiiVasAFRG1cS82lUFYwQRXldYXFT+BHMwbWUDxRav7t8k
PMzRc4EVBxPy9NujFfSd9EdrDdnQ0/ZgTH1cyTVmZv3Ls4/POZcz2IBWIvRjEAHVHdSt67gF81xa
4g13r8uCViQJ0Tn7eNMRf35gh57kac6+Ekg7M+QHl2uFWWFlVv6v4AapGH+jXFun1sP+m2lLC2wp
dpJmsBxxUufoXFFFHoILpQuyO5fAF3Mf/rRdOK2Yc69EvjBaoomngT5lnwTQhFN4gsPm67GadkSz
379CL/DIwtAk1VlYTs5mQiAlxeKULaJhOr6XbPWHsZZScu6Rwt6QMaUh/gTRdQMnXwEQuc3UBXN5
c0QcFYmmdd1qOOXqNxePZoeDm9HTBOWlxUAtQ1HsN0zSfxsXP98Nuch1tckYQHI1EBrTFiucYb3r
9UKu3nydhGCpJb9s5LjV4XEMkw2UN4JtVU90wbR/jwQHJwBG0kwZkO5ivz+ltFrIHtEEVFRlg7cK
uPkjxXvYdv7aI0lJS/U94Hck8P9NYPs3uy2hVEOxAgZT5mPWmGtJwi6eKW6W7XnAIgPRL6l2HgGR
Upazi6Ry69YLXwU503t+6D36jmkH4NSVPC/iSOXG+OSJgNt6utT5LJ57u8WM7Pj5/Df4XfSRiPw3
uD4ZPpNBoaLACbY06V4XZS0AiyloX1P/Ugu+9uS9zO1e9f1zrjznUVr8Jv9gHvhfiviLlcJFVyzQ
TkthP1WH1tyaeGSY9blWztWsm5Kpw9KqcIlNNq2CMPhbmTbNo+q1YG9OU32jEeadWkO91xBzqsdu
z5VUzJgImsG0BIggdNEdx3D/p4GQBJyenJ6NjCeMvACmwW1HMhsRxMwvmXIlL758uamc2HANqFQf
CiBbxbuYtNZLxnlDb7T4gq6AioUsSNoffCapQizKALmvG58tWjpwuMj9oC+VYGndmMe2qZUXvr/S
RDXQrt9Fa9W1KeazfGOMjtCUV1BpXEZMd+fdJz5l9anGhKvKmhx4UHi1GVohzaCdsDSrCMA6Q8ni
eorMir+w33aPB6GXSrx8co0cZfE9ltFgCEKFt96/kXCOrHLX/QdQyrM8VNnT9njFxoe6mwIimXlK
OckCNS3dnTAP/2/7Ylh4sYC9FZwQv169HCyVrJQUPNz5v/fjbweVNCxsadXGO86R5k9mlTGYDyuW
YSKNeSDtcoH7UPK0ndU1P3Rdgii7hz2/ZpFPuXUJUuNq3/cHrQXiFVQU7vySJdJ8Cvh/fNe5Trjo
MtYWNeclUo7ErjUBmrLVMK7L3TIOYdkxddAYazHBGWcqbdnzQsIE46XMunM+nMl4oCvr7AJyPOja
zAO8Vx3KZwmO7wjzSXTdcmqeDHdA8lTlCf+xOWm6lzT/tujpWDEO7ymAb+o1NLdi1aiNdBWL8g7T
URdvFgNVK06sMnv8OBXeyIHOTk0B3Lwq7EgDiUiLb89RQoUG0EBmXFu5jCnixg+7xInWoP56EvaS
1ZzVrNMnNC9QKI+A6V6a5+D7uEvXg8v+iXFfoKI7X34FvcdIaMDsKviwnRgBO2VLmXTnAv6cV2Jw
2GsT4ROKswDv2QWNZjKIhFdu9kCPUyd3jwvFttXE5in1lBTicFQb22NWZJRzKdMN0D9/ascFhxJh
U+VGKN2ceQs2HnVZk5Fd0CgLUlTU+DCLHs9j4buKQsOg5P6yj8eFY8pr4w1EZjtV7C1maYX5ZKWd
k8JiLAuYGsTIG4n5zSs0H8rDHcnX1tlhzyaj7qPw5DSD2DS6iouJ3F8WFM9VVVuFse/CRhBqy9IN
ZKQy4yZANG4FS4c/wgQRemBTmIWjnEemipWSBMry9m6cbG31EJ/An7+vKx7CaS8TryN/cby+CWn7
ZiCZbxtyPE9ad5NDsGxOwXJ9gRxpmceSvTXnpvJKOnsICq9vk2x/oPcm1cMgyRBls08y3Hwagq+k
jfp2mSr8W6aiss5Za4hHRID/pvYOLds+/X4ZAkYdhiuBiayh9fbVlQZbLdH66mfkh1JWbqc2MVGH
XYOjroyyvNiwpnPrePlQ1R0503G2AQ/g5ve5SCYMBGYTImP/RnQ05nkZJGCHVkhRfPEE5zcsrduz
KseFvYyIlXxCjauBich58CrZFWvKNpWgr0esqPTsZ+CdqyCUunmGsqmm59OLmDlBY5Cd7vCUru15
4PjOkb1NfYJrdiSSPXmVld3jdBnGM5B5MayDKBW+dvwBnST+bIrw3AZvOZR558fzJa4afCEHex7M
x83iMQ4IjDD3yi8QU1APOq7D7DjsTaxFCRbCYzxs7kHpX13A6Ce1iCN0NOAvDsL0QlVy2mBiG5du
vZHlDZwedCPNeWN1dYV/dF3/7c9SO2JU0oU+XLI1CY2+t3WHtd5zMYuE9alLV3yy1OHp6TxK4IJj
15FPfIt6LaWOVRY7VUfX2HqLZO9wZVyJ8cgSwsB/TBIPu01WfMoPQJ2VtT+PvZBgiSmBb8u+W4SB
8lc6CcE5uQ46aiasxz9C/pNoEylcmzdVHQBOC1j1+QEnzP+c4vmVHUxB5eIHl+2NsXAmu0IIefyD
OUcB9g5hSXBCEBXiL+DO8pdOOHtp3RjcMXKdUhwXNXZtz5HAFgt3pfCvLKs7CNIsyAz9a+bVDOG5
Wq6fIFATan6ETKlFSraG8l1P/a/TtXItDcerr5B6m25hGE1C4Hd/vz7rPKYs+iz09/24KdlJsuxQ
i9RlBnLn3nlLhFCI2A0cAzRV+LKIySOevuXc2I9U4EurSHLxwLXyaFwjP2CxlT68IGZn3HwP7N10
WNTx+XeIfvx30qFoGXEHRpeRMfwCslzVUv3PLCBA2fm5r2sTGOD4W0tK39z9ygvdlftO4T/+TfYL
mXuxRmdmmyZGVbnBYYhub8o1ZFMCKy82GerW+QsvT9ZnQmrBATyWiqzqHHxCTI2fkJPB7FKajh5T
FHvvFCtEesKmUXj6cPANsCkbnVh9Uff9dQz+0QGJzFoKk4ycliNchw6ybKROwHtpWnL429AO5GyW
IWsunATEuOGBF2DTMUBPFFSwSSCyXB4TKr7chWdQU34jBwAUSEkl9qnXwFWtanHxkNzzy4IBboJP
ehlCkyRZJVFO1D1+QJXi1YyI1rZxCN+wPhFdac2RPGfvT07AEZh32Asl1K/lKanYaCIoAT5XKydi
L7zBT2cgwQnPDbdnbmI8D9g2n+NuOj3gEbnNCn4xoFJ/oKdkxW0a9qP+SgpkC/rCGvW0WFdXwsJA
j6g4t+4Rdf6LDhoSM15NkT7tENlBGRX66ZdWDwnKd3bwH0mfHVDVWWWlANCRCPCtxcgpjnpFrlUZ
DcOgA1Mdh9FCTJfzjIgI0u/cVlC5c++6XC1QIQNrxb83gFBMxrJ1R/3S64aPjcG839Pw4trX1Vlk
Hpi2NP7LDTDd4opCobxRRalTPTvxihoCMvJb4nYS3vr+IwMA1v6WgX15LfHfYX9CkO4nxX2afjLL
AErq4uoAp8mYgYSJj+8ciFEmBOBH7DktGD8OTIG8m+lEsDaQjZssZasQW+Ma8i/ffz/id5cdBHyX
Mu+SzwYW2ee24ZP5iIDvIWfn6ok2I7f70Pepfrv35OP/tdc0UfMBSTxn0E3R3YzUzmrX9drpGzwk
kgV106Lh7YwMbeWATqZnGwhNsVuw+wb/J7T6DChEE4xElQligCfR1UvsR/rHDZ+es+dN1IPVOnGn
UcAyajUuEfrS6ijnmSQ6egYLOzE5X37ZyrXJCNQ7zJk6nwkLIE8GlkOscStEkhXCDMTAxLtKp1y2
s275xNaZ2dCXQIVaRssGbtABbcSCkO2d7SLhAGvvG8jawF+pitO+DHl8PbejFebY5SB3i3ly4fHy
49ah8s3mnLbvS5QfvXL0TR8EI7LiQN81MSG2tyz/fmlfxXimi5mn4qCmqV1O9pab23iYumh1QWcb
5z7MBwNT0Yel4tJZEssM+Dppx2kHOMfY6qdAcXTOse6UHiUZDu6vM0b8LIGvRZhwkhgYHZoqB7uX
hZfZTPqlccm6rcMnMLqXtg6++0YNSLjlX9GtBQwpkJO0SRvHXlyv0VZ2rZz2lxG8VmwlVswdpjpI
r1PJJkTbduyRijqu0mjzDagFgZPowi1hrimc6jsNvglAf4xINg2vthqWaVe6wcyxH36TuAsJqkL8
Bzs24UMxSAwbXsXcU5ERqAnTifVgNLpnPViauzOFiNZTmXFHTW8poq4rHjJUcF0zxJ8a32KUPExO
di4p+m3SQ5z1QobJYsv/ghoFcDi3r+MMdbvUUW4lKkTZMZ6sStCbP8O7fM0tfnfngLM4HKQQGa4m
ou+gPaLfPGop6enWBPIUnHkEds4ESaU6Y5cz60Gdvgbp83hYl7SvUvKNFplYU2ZizMCymnrv0RbJ
Mhh7jBnUgXMAPeFVwml7TWdATAA2YvpKIbaGKZq9UoVZAUcp+S35bdHrjABtyxK1/sWCjlvvUnbC
T4tc0Wa/lUr/MTsvZlAPCl29L8olhgUiS1hGlztDrgzCXkahgIsIo06As7K7TxtC21Pr4WxgLep/
0d2BChm3Nmfyhvo9wiHwPQLLDCkNjRVciUG/sUYdfM0g5QHobUSy3+P4IIerV1Y3JUfmLsMawEQu
RE4qsvL7UPug2gUSfoezThIq4vMCarQjjO9A0DNcbjM4WkVUhlt8o7TqmS2ArqkHKmyD73S6vjco
emrC8Nhl9ukj83U0i7WJ4qqoKxenFtwhCxSwmuhYOuzmMjqcnKtuIlt29cIkOhjPgeXY4hh+Pe0u
CZfW6bpw8sBiWolWGC+rDblBxnCMshMv3kshrLKpa/QpxaZQQEoanIJ22zF/Wfuf4ECXGI+cv89u
TxA2RkgpMYbLU+c/8DMLmc/HC681vwIeJ0ZT4OkwPlPCtT/rDWRixUfLzpPQR/wpfhgfdXjez9Rn
5fq/rbURPlOCkh3SZnkqd/0ZRxFtqSILkfq5M7sVwtgSExv8pgmadjAtKmaV8d0JWRXZ+Gxg221r
sqN6hyyR6AiV18USmwWeX62EtMPFKduim2hAOjKFYKj2hwk0wmLoe+cQ6P8Ew+8KosS+6iqqpanc
Vm7+xUbZkwWDzEJAGsKSEZ39IZz573Aof/E8O1pp0UdyqyiIC2hRXsAUXSE/f1+rVIDdUd41+wZj
sM2YxsT15r7m71IuCusppgLaDB6vyRTPNBK06s8fZCJFJQqlq5/TiZ4hZP01aiEsi3T/3IW64QHA
0p1fa7IqIcpaPyvcn1v46Cu5vpREpe87SAb/mNBDIR2kwcbNsHk3e1nv7uv0/7eZA3tD/One/uxX
2nIW2aMdh0OhdDi4CEh2pjPkX5lu7h07H2njyeIE4MAr/KL57hsyjESV4KydB5TBipYliliF4KjB
WQV6xVY870KG4IZF35vLFopNVuUq/6mKjjzfiDkdZhV4dCiOx77H9/MLYMYvzVufTqQEOo4ZT+WG
DfPc9BCTi4iNohCrJLqxCuueFoz8efDk+qMEhV8CncfcfMmFAX0oan48jGZONhOY2doU5ylN2yzR
oV8O0T1lFQrwBiaHG25N55WlwM1SEl7bqp5s+FQgSsGv8osZLyWl5nxKwrHouvIIOeWl2r3AWGmQ
0o2XDmtKKUdafhDOtojqZXeMxLkd8stqbeTyJ3jBqxn3omsRUZaHI6IGwcp+r3ZMUJjZeKKOkoda
jH/9UWOsCoE64RA6MM9614GRWpPnNyxZOFWmd9ZXMdSn2lOqkKInF3RmrVKrBNhywxJ+guhTgVY0
3JWnYPV2iJWc4uDSdLcegpMbZbASKOlTNKCr7jM1uH35f6O5UIq8UeZOCox7DLsEdDawxezVttJU
5D/0wI6XTtOXb9lJPUArSBF79CnmOtUuE4I5eK+d4lCmfR4C3EmcYh+cT0VM/kvIuNBDh/Vw/0OA
RiomQzaIRCc4SUSvmziv3S4ZCRWDlgXb4iLUGqaL5cRO8PlcPYkMmYB4mu5mbqCwqUm6aaMZ6Wk3
d2Cbdif7wMJZwmwBkAOjY0Idjwfbgm/Xs49+csyE48/bQ9vDZW//TISozRLy3BImrUb0TYC6Mq9V
aVwab9vPEqdyLSB6IbbLEA5BeCldGCHeYNKtXtY1ZUnmWFn38ISLIQTWkdOiFFK0qcxau0JyjdTz
iMSWyACHiCK0soXyyNDWXoKm+/kinacUyy93b15gBFF74PAH8eMCpX+tb1LSuk2rocbujHH0PTeZ
vi0iicCi7qOf9sYVA++uIHxsdiqz2SxZ8vE073LhTcEDWfgDGJqxqA42o6o1GH/E1Qsx0cqpAnlh
sxukemR64xcOvfwWU9LrwH8r1AWUokLpYeAnzmDgDw+NkhrBm3TPGHOrLpKQ4+TwTSwLz18ya2m7
QqvZW45T10Kj3mEl2lZlQADzazQyXuHG3TES+KCT0pEE2SI9xmRYW6AJcUyKBO5re5y+ppQEZbqr
EzMWhnNzvicmDz9mNSzcC/vjMEJdJ+a/4kbooLVyG4IQlvZyc8Nguub3z8cxZf4x4hhxFvqAwSL+
W/o+ZbvQ6evNtGbEPKVfYNygv0pnRiK/tpF+8ZMXzuOY6rq1TgBoBQE6rOH8qrgDeWbWTVaqHrpG
7lXfXh+HcHg6h7bdDAP6JL6rM49Z10uqINfsHk6mQDB9aEgcOPfK05Uv7AwzHumNt7PxVPsRLTHh
MaRPfKadmSpUHeV5+OCCUcxyz5h4mCfaesAZdZuQLjUPQKssE1dll1484DFgO4PQit5Jhuu9lfsH
TRZ88XAfNVScp3BkvFL24ul3D0jJL6mUZB0B2kWg8uWqps/evbEAhn1ljXhxikfooX/iytsDrKnV
6y+H4onwCQ3Gq2IlzzH1vUgq0uzzoMl2l7/j4qqqBQR7PRYiTF0HuqhB+LMMShrS9Tqu2CzZ2K+n
DAmf073Wp8T9PGJcqLuPWi/HTW+BYUSNpY9eMrbskWpEHC32UuYsK96BDxDJV94C32CAe73+hBSU
TICAf+FssS2Uv1jAUS4lcmMNcXHo7c94XMkmotG3Xtm3/bJZslDfA+urG9v4Jj4rz6LGPcP4c8/v
eAaZyhM5DJR4J7QkJhgyJp3ZtEGKcv6AOrKPy6+avboseUSZ6ArvkOeHWAuw5szgwnWtRQ3rOZ72
t4KZFA8ST9WMx3Zohlu3+l1MqCRpf5PfRomden097HRBxsn/WJDeTzau6gxe+Mz3iaAjZNkOvb+j
zgn4eJTkOSiHUTaz02fXOG2dDHCadUCGeebtS4Ijpd2UFYv5iioZaoqYk19IE1+JHcxHMD355BBI
E8kv8lLf461HupuUn0DojtHe42D18k8b5eUwvi8kXxlqsxfYW7shbWi/y69DEWbwKQND8fjTr1YT
v93ZueZ/131kPqg3Fffxm+Nqg69EaNW/GNEIXazGWmSqGNd+YQyg9NDYJMVeyiQ0slSdj2JDlX75
r7bqpVG6sYqQeCBNSd/zpkBks+rDEFgDo+E81UzowbcbsiNtCmQjoFm2qWQwtSFPI0nTe7NlD5LR
IxcXBiyCc7u/42NymCJeb/XyzoQHykAnNXbRQVYXaw2uITPvIgX2trx2G1a9W/xCgXdw1E4WQ6XX
LqGixPHnKYhWWIy/FdaaDAP9tNFM55w0b8uokwL8RcS5NDiMOucaPm4pXc+HIKTmNnw4YyYPB1cG
8uyy/MmDhYmVkehXmwWrnq6IfWf4PXpil6c9DFjnihrKE0I/uzBsvdmX5H5dPLXpVXLoaFmKC7/q
EbK7g93V93fE4buoeALRM8n5vxxR6iJkrH+zyheZHsFREWAhD2bwXuMIkB6ITc3XiPGZ++n8VL/A
3Ef9PS6Y4+tRcF8y49u4E46EhUJRmDXuulONpt2Mf6kgZ2o3t/KCQdddldxh7a5q+/A3Ef5HKoO7
DVmGzQrXYqKv8vwNYrSbuXCFniLI5UqLb8paHxtNJm3Vq8DNRfLGTpJKvGDuoTpYqw62QVSi2L2/
lSiNTAy1cgCG1EcMR8533TU0qsCWlL/kDQBQKDrZEMcVOS9ApywCismrb/sJREvaD3Pb5YgIdS50
OZ2p9ND0X1JQfbjPAvQrIZdC8fw72XFErAwOjBT71KpEjLZi/rJPXKvI62YrtO8qhUF14w//DP+D
yNXWxV5xOKAMhuOhNgLRm+PugijatVRTKXa9eJNUmNkmuPYNGhQyWIsQ0iODdAdTViIi1VBrycit
gxW5YKYG13sQlFaDhfXJBsnDlQH2yvDGQ+086b2sYvyygQtIQI+SNFVEmtSG0pxyK2/3iryRLcvI
hNT1W3zTUn/b/Fqq6JS1u3ZCeocsI30Qd3iSDEz8TAjst+njlkEG0sEEH7KmNdNi3RsvuOk1Wu0+
K80/+ppkHulRC1eEnutIUYjphFcgUYqyuUyjtHTLF68DAXmVupFMK338uMQDbEwQ9/r7i4b/l3+S
Zq4v1Fek+rdAoOos5PgA+J0aKt4SM1w9zRNFNrv2bVwgm+iBlHZZimSh7HghKeqaXLJW3ViB6nMQ
hyT3L+5VQLAkBbjrDmJyd7mO/2tWbk9FXfvxmYYjuECaLBXaonEv0O/Y03DE8xizWiSk9iIUepV9
HnYpYf6a6Bq9dAWjK5lvgeSpqQxgGYk2UfLBXQqAvkSwjFv6aJyMBeMskU1cPL5hNBcGbIV/tvzo
Gr9NUNlaP7+XiugiOUvqqVt6yt7dHKtVqMAVF29YeG2VwqIfNWPxL2igxD8CSwlL45xdYd7/nV00
4EHgy/PikhRDQj805qA3oa2BTLBzYGCxqZ766H6WkSO3kHh58nGIj/d9U1DVzvOCIwfDB9YGctB4
vv+Siu1Geje0X8cevaWquOMr9xDguPQ4Ll7olRpnN58CUaptKwz1pkLAVcVQgIX7L3HGMfc1YdmE
F7qR49mSTWdvWbrH20TH42oqqoZ0sgo5yOtPirLzm3thV6rXWdJQakwQ3x50PJ339c1L6Fz7j+ho
U6mzjrc3P/e8Th3MnTr4cfbYkeYhwMYF2RQm0eLfp8sAyknSgeKovc6QuE02t2yHOU5ld8EA6RQd
mCA8QuITWMl80jG44myK5y9YLpooxC11d9sbw/x+UOsqQc85tA7/tyCAv1vFw6MtNB6IbBEXdSh9
mEmXzMeEPpYRU1F1DMhHCuGTCV+gZyYTEmZOdkicli1tJ7a0FMK/zkLkZ/G5Pda6p+7cmP2g2e25
JlgIJNr/qlEdGHG3vTzVJWtqaM43NZZnugBv8569Dh4WsV6/QJhl1bvaT2wxLrJUNjOuH1pq7I7u
eQm+uN+9W9MVjfUXLG6XFZhe1b5ww7PbKNvWXW3QiyYLm70OrZz8y0vxMEXXRH92flcjPw6eBPwf
vTTdr/LXCOGD/8ss4hnZRuqmCtkQjt/kZNfT89voxNfIch9iGMeWs8Tk4aQVrr1WCUj58xghTnhO
E64C71LqgoC6wCmf1QPcJHJBCiSX5WY+POmFgyvVsDxx4Ts8vzBowhtrDANHb4QJHpOzRzemxb2g
hkr/ZhyGlEByycK/sAkBiekHlky2AQu3z8+YBPPQda9FwIHT3GbkttC0HDTFjNwYmUlvmqvhJKHz
9URDMz396G8ZGvDE1Ak/YVkoEzwKELw/Asr1hWJDOTIPum3MtirrNju+yua2nXVhAj1hQhDi3xGc
af3RAVzuzlwsMIDuCtilEKJLdwLd8I9JpVNcDfkYCgPIdD1SQHvFdiNJ8kc+pFssubsQYkkAzQIe
DSFiu2/tIsxH+8V+GqS4gx3Y0BOUBS/00qifat/Mdzx3wjRYXU5z7x+3wrlrvvcpFK1AH7Clhm7O
ZHCtOpbHyHNzaZ2MT+zW+Qm6Y5ywf6Tx8IvqLwEUN4B6J2VVPws7H6xpSX7uC/QUMBlIYK3qVnTy
oPKV+ve32RokYpGBPItAGTyQXCqPsjrOtpSO4IAao7uml79PLfYjd27f38vNrRhQq0R4CJVRhPMn
jjJWtqtP79sS+eSSR83t/8NlibAuvfwo5lstun3nUWG3Zc355Dj3TEZxEoJThCYZvzAt4qGB+Q7y
r7O4NZiV4tK8rIJLR15Ndt8yic/hLPjPmeo6LzISJxc/jIZPt7dkxGGRUhkSHR8gxbn+BBIaQIg3
q4uE2IuHp03aRY8aAWh7w92mNlR1ebV/8yfnfFyPjUcEMOmxsMQONGfamCL4qVim5WKF9JGFf3+n
liLejyHV5/J/ZnK30zauNRglI78HCCmdxjLLCbYcRNSNhQ+Jr7fNXNTSRy+KWOpFpt9nukF7urSh
wVbqXW91tZR2YPpI8/RDENM0XTcimlhQAD/7smGswIcKb561PjVLJRGrT48749WNLPocHTPZkz7R
MdVaRtIWOEIj93CVi3DYeogXklLGEn0OXl4yWP6cIq7dXub9dW1WE0QPT6vUyo1rB/77Nm8mNnU3
FGXCMPfSO1RwrW2tT60f7U/BUEyucOQFRIOnS/a/hS5buJ/mj8xmKieeFgk9fB7eQe/S8GuhAa7D
jWdfpJYo8HLAu99g0xCsgXXPc7poMPpUZb7aMPDWt/WOFQB3sAvu/5Lx9glIwro4cW8KVBjWUKRI
33DILnMQOvMp6iDoGo/EKCO/TZc79dj9n5y/eoELFSIvqWzJ75EydYRYA7+XjJTPgmKR8JUZxrRi
qaeT+rbxh3wLvPPt4s19oG6CrbJj5fqyY7d0GOM3qegfT9pTXGFEzpC1lL3E89AhJhx1TVoYrOh4
WDhaSVnshJrVcAJOWx7T8pT6KiIDDcxFunXwpoOcS0zaKpCI0sx0XJM+VlpehAgZC8cFsxwgPldB
/HWxrfjxepmgc11f12UYDEOkg8SmeYy9wQPVUbQiAH3YdgWMfpgxiMyFnZWSCslt139H1kaLzoVD
szaAuRouIzlI0/Mm7DfVPoQs2W7gVWiIpeBji2mw/9Oq+sGh6kECXiaJSQ3cxwncNyLsw/lXiMTA
mR6y78VpTmY27vSldHFKwtzjCzvQ+Miyo16q/C58UNHa9qAN3TYv9IJPPwWsbKHNLY7YIZVMc4m+
NnGW+hRb/ZLKeprwu2wpmpRUZ59aUGn6wC9MgfLw0gCthdUjwZTOcFXJLptednAfcmFzVOL6Mp51
C6oj+GgykbOPt0aCMEjRRVtjx1a02ZLm/KAmoiDPB3Ca0v1nv3/7repJJ4NtECeErydpgtdP0rWj
TRaZ0idggoninx8LbkxlzO+9J7/X44jjhPLz6iKXz4dGRih3ZbKPLeswpKqW0CpyD7dNavpOouPC
im4fIfjhqI4KZxAIXL5T6IeWIiFxLbQmCAF17O5pGGqMkSW9j0zlxWn3bmshly6shcA25YEV03sS
HOIIXybEm1vQHOTVdCegooKyP6mINFzplLtqrvr15Jq6kI8odlAiAyt6RX+H4ExCzs6dYrh5lat1
7fRHyc5RCAO3/6UnhxwaR1akVC305G3InKLxjI01n2q25LkBEDv2igReM958CjYYaRudaZwKrsiY
Vxy01ZZZU0DHwhsO77lmoTKGP4/yt86k+q2HSLPtHRvjPAf3RqKhmYcSqiKv3tf/5UmPXaxc/E7B
hBKVVqbDxtVp6vcxTxaV/8vqL971TpxgAfaKqMWNleHyhtfPxWsJKSxGwPhQk4WlPZ3qcIpQH7B/
Fxv7oKz+WAQohnGNa8+FpeNtSKf8/rOkmsfRNAkVd/ctWlnY0sX3V0vYued6rFn5UZO7YHtvPxVv
M/GIdT2gtOL5mU/g/U1vyAYYBs7ikKX0kDGSvbwe5YzX+242ThibFUYEOg3MxaBtc4tEgHEvivtG
nA1usqYjPwMtieNFYnW1O+lUCu6Ye9CvFzqghi51DkMt7eZIW7HXpLL2GOeKet7Ky57j3Wu9kQTs
1a5cvxAma09L+xiMOrGIqMSeePfAATrV+n8hT592VB1SPW4qnRrQQ3f6VPIn4EXhxDygYA4GXRMf
5Qj3Anz6vzVhcjke+8jWXEilorkJPkHkIYVpPW6kjRnTOG1PCIyWeDhfGA+twzxnmO+tzWAhgcwu
Gu7ni4D7lnqHL4y9m+J9UX0YLMdo1emKwj5sVVRyQfM5EZMBX/PSS/lB8EAo6nx+doh28A48nvyU
MTsT4OBQc1HulpYjAViB6r3DsjIStKvEbpaTSDbGcM35jdX8ZkU52BsiirUXwr4b+FFZy36Paf35
jpTrdTukS4LmZaGWlEx16R5y7nRj0s8nGJlTPwo3H26EtdM3D3XILy0n3y84Y8QN3mz74TP/F7l4
ZuuLfba3nAr558/znP5wgdwe/5PHO56yfYjbhbb61ZxVBZ7NeJ5VGs9ZkTPKfFSzKXyk0RlOoWqJ
ZT5lfnZpipNGdFSkTnJyjjL9s2rull3TFv8DDxYueuZfFm/jCoeqeA6TIxj9tnPSkPGEC4RVx/me
T6K+nnl7U4u0x6ZfAbkm5jfTqlibflPz81dff8hbTaJtUe3+QuQlqCJ0/y1aPSWz/ReubO6kvYJ6
iu4n6xJbwzf7n/Zm4RJEqLhdYU2NEWw45zu2w6e8Pq6MIACJ8xssP0B47UIZZaFB14uhqbBdt5Dz
ovKmdUPq5AINAlVhbWCEXbFF3TaRam96YqiB5Xp3VHcHmLwejqxQwrhkVLsnN0rNyhIV1sFJl+Rk
tPsbdVC5+MmqkqJx6CDAWFq8LEUPsaNXO6uX9l+zrwiCofynUVT13e/yc1aUnY07IaO7NogNwzj3
xg+aHBtEFUbXuqfPfKdp1IQAfQBL+tCiztLQH4Z/5TZTuj4WBZWdfSXfbzZVROBoQPTm9wceuxGH
MYj5ZStew9j8pnKuy6A+WmNep83paJhbEoYXst9PXMxTFzR0zodaKHjw4pL1r5qtVnLSvtKcxgJd
XEi6lK5h2GcQJl3w3qFOHwC9mosOsRHsW6HQb/Ll2EY0CXkIcsIJBNyX05K9/7HiR9gl8RTH/L2U
5sGz8Z+XnE1MqgE6xnJWFDlWd7GuxfWCIEG3Nm8x0mEyTIlr1OwkgSKpJlPXv7y5TkFkII7r9leg
q5/C/W/KTnqpRKrHJc8bVIIeEdQvF8nZWLVfrxT7ieIfRSBfskN5VvJh7LFXvVEv+rl9D66+eJdq
sZJ1UEFNr2B9rqu5mhdNxwN+re8y0Znx9GFUc19OAtOCEXKRd6SWQppAGwfAiWkqC2dKTnn+hHpZ
exyl0PBCM8EJ69jHIRRYNo8S4C8p9HqFRbI2lLjAIUNhZHQ8Jxm4aYnjq4h9uEMVZRJinXHwiJtP
20q3kMFLK+QrtKJojjtNavMwSwqs+X/Luyo9DLwDysW4QQaoFzoB0pqZsMjZ9ML+3qB9+OF1hoG/
OVEdI+YVbpjD/3wjoHtfOfbHZm7X5oMibZP79ldWct9mzqB0pM5KxBfLmlKIWpeva46rmjsXveh9
X8JSKzpOqixP7sA6vHi38QNKnM44t/y7t7SX24ZVXFuKZlpqZTaG/BU9kFJDVSsQJyUdpC031bG7
Jp/iWlC2/HjTWjj/y7eONqvbcRgGFaLr5cO16MuuCnBJvuPPQgT/Tn8bMOq26GgZwO5+ucush3ZM
kl01Y3K0RDZbZ9eFfVqtY8+7QqmPhifESc3S2c9vo8iSLRlF7QrSxBZ91E2hWxuowpyqFCdy4QuL
r8LyBdnLp8bur/8fbCXHFQ2jNAT+1CJAvVIG3C4yTvLTZaVkXu3SW2u47YRgPtW4te8P87i2mMmA
wjLkLT4OcZF3t0EJ6EYQTM8trFMo5ZLZaZW+S3BlipxTMz4gOz42rbwfVyRwIMSgKeCUTbdU3hLP
kf8EvpEoTheLM5ZKwhgo5h1JeaT9pudq51E3YOVnduApodu9SegSLFn/eEIbMjv2ORT/PHhzll1g
2q5+OaviEvfwoCzIWQtkFtRv3UNX5mgC2PIoSVzHp3pbywlQf2MJREzvY3D9hXcqVRid6j+8FJ88
qeaZXlEXbZVpXUS8XjXMFbmCB4jalkLMO7s0U8rabbd7JMosB30WlOnoB9LB6s7/L5uwD6Y4xA2p
FXVD61Ty6vQx6huBHp6LpSZNy6QxV7nDFYIrlwRkIVY0+MlhXvwQ5Q8j+yQBgXqlBvXCulIxV4iy
6tqUVxMOEPCkBHmsLZAhMz+l8qAegRT0QR+Q/Qi3G8Kmtiy+U5Y5nwuZS8U6QEB2p0D+BYnLgnuT
3tHSRkWuuKCkFdV/Oh40DPbpLBbPsB7BYIRC3ephW5Q1VQHCypHKInTlLbdvDpI1wxL3Cm/q84gJ
JP+gZN/I7gitGLJOXloY/rpyNFZxrVERe3FKnmyv9+6IxLc1ml6fBAz8BxsJvWBkR2KvEup/KcLc
OW+bd9qDEJaDkx00hOl60wV+U9tQNzNmC3e+2buMbJU2Z2jf41rWmyhupkMu7br7+Jy/7KHEQqkg
1kH+AVFVklpjDeSyJ4Hxvgs5rq0xk5NbXl/2bQYl00ruPZYU2Y7ngwB9YUF3UFlbHOw1L5rlIepn
ayQ/C6PHQ7Gv9vSTyKmzo9m7+6YbEjzKetezpOQJ8MuTUEZzJ6x2juTm3clIf47/N6vktg0IIuw3
qpwzm7Nu18TU7nSJdjYsRvefiM5kchSWS9y3IGp7/QOCqJfhxZOdX6M3fubhQBDmQuBWhQS2vSOv
PxFoMVnXWquPuj0kPQzb8cS0ypp4UW5tUChErbQxo71u1gP7KVXrmrzf7fLGihPU2nbZ2euK+3/1
yxicoDrQAb1/sSvHlkzbbPLlV6fhKta4wRFEfS+2gVVmNcj/h0iEPseA3jo/okQ6iPPZHsv6OPZ8
l2sGwUnDmgGkWvdeGiaKlLqJef9ZAMaXNaziuKVovA0+W4ZM+cxSSYnqfFhh1F6rtFQSl+We1Hvq
gu6RWMb7Z527/EEeULGDl5elHIsuhXOCGASVBqpowIWc3gjec7EGB2okJazcWEXdKDermgfKRohm
6zMpsoZE3TlitU7Ke61FvVGWqPyG4x3ut/VAdGq7jgf9Z0hK+u+L1CApbaeIm4/o6cxZycyy6OWA
PL7pTb+EwydOZg5kdlr8Foth5Y+EbAW3mOOu4iWBbq0+9NdJTS2S5jqjTssb8F+q7lCk1Oq5K97H
p/D2wVdfp1q2sFeDIhJGM7fBwajQWyescHVRVTEa7q84gU5VuPnLYJdMsFJr2QuMUofWSc+FPR2J
dss6TzADnkT4uYETWz5QYEXOvTmzSzXUfGh9xyHKxLWDYZej8deK1z+nNQKOWRqsyQpHuYkjHiPY
A7OpAmyzSiQxYVLACztzhdh1dl2luaz5QMCdV9poj6cUPu5ol6Tir6xTYyZw3fhRpAJ0C07t0gX2
wy61PKR4fYUqcH3biEuWkLmBFEzqnb8P+Hj0kNBFEFbRtVOhPkp4tApcId59grQ+ZVCcGMyKCQ9p
0XdQA+5gTgYrqm+JOZlNcLn2UHgSpoZfYtTE0gH6Dbh2nh4HMSx019iuIGpW2uE4SEm37DIcdiFJ
/PislDGULwFi12dSmXbs54+tIaj4X3pxoOjD42rplmeWQuYmvurjCLTND5B9T/fn93EPpeG1zqKX
aNVEr4ydjlFAbuCKWDoYQTegUajGvZsWxSvshzNQQm4Xl0Ahr6Q4OBzDiCHKluuc8d1fsXw/9jaA
DpLGWqPSHJEDjtaR0zPvCW0q7kh2Y2yQZ8jZDshoti94ZckLfTQ4zTwLWlGARgzzpY6l8X8/a/Vx
zMHPyNAgdvBFGSDM+VBWxaQyq7gSUmZQkNy7xPCnr5ci6b++2NwvlJN2eQ5ci1qYCmqmAcaxq5Bc
Ggc2I3mF+bzEhpZY2FKf8DFR5zV/j5f2tuOIHtCAvUQY+zmBTyX+VZA9OIId8AgyWMhCnggJPzpP
Mxdj0zcXXcbAOFSkbjzohkuUGl7s+8e7QA3EcRLStOtFPFgpesuuP+qHMqxpKMUziUzJK58KjO+g
trHTAYm1MM38y76fNWCiHeCcufB0Rpep1kEAhuF8WxOW7IereQp0cURt6lGPHJ631JPnXYvh86Nz
fIVlL4/5FEIKk5SKcyozKR9BAfhSCe5R3YkBDtLeWrwxQgUhXyKg9HHkFFvNH0e5vD8dSZUOvcsj
pQ9VqK202TwUe+e/ABA5mmqi6A536epKXWlqwwUYkDW4K4IuFGCiGvUWLqUNN5hXhw4a4N+5TdIr
/MOdTjZx6dwC6IhaQzrLTLBjQxjs65V1ADDBfnCLOBrbapveU+slvsoGS1yi+ABWbvREA063Fjo2
tDua5Lq4sJsAQyKXR57rhTcugTETx/6boz0FrtcKZdgrR47vwgJhC1A9FZc/Y9UWG2vyZOLMQ3xc
oQMpqt4X8RyJrlWhge438nBW70ezJI+awbMoNgLRpvCemIqaagobaQHOuB7EhM4WXjAD9ep+YveP
juH5mh7IaiNfRAo54RdyukEfuGaqQsTaDnNq9N0SHV58B6V2AgxOrZgLKjDuRHwvJi5xfZ2Cl/vD
4O7hxvi2Ts7ewxIhaSLST/fScb7fHB63wx1qKqrDoGgbvPvb6nY0K8/8hvnon8qbAx+MNdu/46B8
XPx6anvQLVB+rKl8htP532Y2nihhrU2RsnSWskSoC5Hyq4qPyDx385PFIMNxNAQDghU41GC8xaE9
ewRUaDTH4XFHs0gFekbBYyGbwrKFg7pDy+s/y6OXSXi2GVVutzQOyYMUfu4nolbu9+UYEdeuQ/Ns
juxyyIRiriqBfklUb+k7K8HJOqLJSBYY8UjBDzrqmKn2iAvErFz9hBcDhXhn+ppoQcJeSULjRREy
I+trL7uzQyeTjEEx2X9MWJkz7W0iWDiFvFjI2shX6KHBvA6RMSgAQuf5ZiNiWYowwRhGKiQzSvCZ
uV/vE5+3j4dYnTVspWoj1/fIrTFvIqI2qLCt+9us8hub6G0bGEaTtBMC57sblcw7aUG/f03+J9jW
Rh+jOdC7HO7yDlmhiDskNw7lvNg+Gu1SxQurNcPR5+zXONFOU7xHlGCXBm20Y5k+h+N7bi0aV4QB
VWEvYcNiVU95E8eXTNEEMczUO4Cc0V9d35QvrjNplyARm8ev0UQKGOkrnuHsnvaWOug3oNPZ4MhA
DBWqWC866JTsRvAmfmQdXtqPn9KaFo4fxZ9TFF8K6N8PMrk7tscgiv3SCIyH8/oXnLiIJEpvkVBs
ejxK4rdSdAelQTvmEsbHDpEN4YFXSaBPf2hkslU700jzF0vfZyWBzncxa96luCW008Yo3Ly5trsW
Yz/Vz7nIiWAknMyBV9xpLXtMy0BlA5A1iX9Eiy9K89zHVwbJF4prmZlhtRUgKU+xfQLJ2OdFcNya
72oB2QWb7v9Jfp3ZVrxg0WWm5OSFOHLxSvR0c3Kd4AKLMGRGoUbf7TLs4doUHgejSmnOWY+vSs8Y
wsTDwEwRcRiIaQxsvaAHM67YzeY6TNDHhD6siDG+um5oVMC06BL+EnH3TVCZAOlFtW77SobyWgB4
lsdg+pEfU4Npi+sOinfygIYNXHacbKajEMKMZLT/3IfpxqgjGTXq2fG/6p/HOV5mAyw4cxHgK5wk
Z+tzGVDwwg/iPW7OrVrhjH2nCw+2b4DbUfurq5W37qUilkftXLI4c8ilzVjqn7dW8KeUYNO6GgfX
YW5RPL699hwbnvwUpXIvWz/XTZH+6D7p69cAsFDhx4Nc7M0j8m+shva/rey/8w0s1OmiuvqlMVBT
xQjHpM4OQ1eDR0+31YNmA5asirhFUGXW8aaJfhCQBjlfs/jz4QuP4axQBE1ePOShXFUd1tsZcN9u
2FmUT5KhfRxEpRCbHbEbt8xjNdlX8UwDMd4NKrJUA7hmIu0XD99JlaUMbgZ7DurgFKr13nbFPqge
cdfKPWyWdujSR57iTtQQPEJCSH1wCArvmWvrD3yp0xGaqtwlkXRUplNxSQsOK+lzSDmeziPFQpSv
4Pt1GSiNAqnQHe6UCzRYvhw2eY0zikhf6UCO+miAEEPwxqHhjD5xdfb5Fz9ytSphEe5FhW+ksKai
HZXc2/DFvk3aX5ho7Lrha1XlXjesyux5H0Lb8TnKOhr64W6yeCVzVi6JL4xcJgOgsZ1NWKyH2MOb
uJKflWZI6+6VCZlyRcCUpzJCibcZOQ2c2EdYb1P+53OKQK/8FEgMf7R8miZQ18ev5Yby26H6J4r3
Gjf2coqxAM4813AyGaxcRYqbMEMOUHG4dNQjteZFYXFFqkbkSMb+yMSzhsDo+Ut9ntugbUS4B5BF
yq5fBR+Y4xoU4xUIOWCmR8NTe/JF/4mMXGaMw6icrJXIO7N9CyS2zGfRp4qS2EEDTK6Ly2QeAluJ
pDBTa+p7mh1hqKqVndHGId0Y3mbmVE8ZaH8/xQpcehngrCgKY8VdSrXFk92rsQchpHEjAiEb1kcC
9PvF1wRmXwTen+3NxG1owsNUjN4QsnzNHal8530OziFtCmCFKWiNC9FV7IACnQy3Ai4EZiTaqI9D
7o0pyv0vVkUFEYsgw4/sRypblbDSQjRBo9/BdsmLAO0Oyjyb4ErDeev5MXIyrNm/qVulFdCT9SAv
Y6ZJgUAqyIoMtoyR2RFrn9sU9bqKTjlzYk0YKpKQVex9BqeAHdZd6C65i477Xs8Ns3i6tVkrS4mz
csLbswr9oXOvDbbXxvNtH0F331ZuUGtuKpo+kddFL/ZR4SbED1UX+H7ETm2psRkKR87Md45Ylxgv
/srReI6EFt2RIjfab7CU+x3efv8eEX5Dq9Ss8xtyOjPMgZPHolk7s3MhaEnIEZfnHm2iTYDnQ/AK
/uy01Ei2AzcPRdpgzzZKrk+BdnBfvSnHud79RUcI7nwNo77XOdeI+ndThjA7JN3EeDDFLTR0K57o
CJN7LzcI5Wo6C5GcP6lqlmtwQ9pd0E+6ej1i7LKepd5QSOEVO8lg0gRLRG/7kgGDOClZFtRQyPrM
BLvCcdq1SocuUDirEnWRC4ItJjWcNs+KJR0BAC7EIejn8x95lY2HYjRxOgglq9j+Ajnf5QjWCJ6O
0OHzUZag6RigjYP7s1SFWKSuViS56EDRlrta2EF+ozL+ijN34SbKiS467gOOkvbWqRNgttl0NySM
prWNazr1nCogom4ZOE0yMue/mT9cwWaIBpExPsUE/u9y4m61vlyxRzD3tCLlQOGVQriRDdTVRL86
fZgRWrJ3dlak/WrST7a/toGx9TJkXiQAdWK4X+fPeDP6UR6HFvdFSfwKSu/nw9AFDLihF4evfa29
kHztiX6iPFcCfqbF+bG9noYJgZLlscT7ILWzWdNJPtwgTrRY0m5YixKM+yGlce/U9OJooV3kMFBO
2OGPgWOxkLuquKxIszPLLxLcBo+0P2SQM5BlbU6RHfE/25w10gtARu+J96HfqYMy26/ZJ2hC8dNP
rRRynxO5RJYWHvAd1Pon5sW0ShcN+tG7zag1spZyXGg7Kv8QXMIbNu7CWHxRffQqhYyc+IJ9McBo
u6H3B5evHTXTXHXq/6LIrExoi5cCGS01PYmDsB9/QxL1QMaYjDStG8YUJYeQInTK5QXfRyOODNr7
45/Ol+HmH59HSiX2tx+LitIhKVSVvHAvivv9QynmPzdo+076B/+WYIC7KunAweG98kJ+xhU6OG72
V67ne1wrnuAdGJJMbK5DCSx4quMO10KEVcaSlg5S+DIQ0rTuiUiovYtL027JEgMz6v3fKf+SmvLF
h3CFvq0t+BN0VLfvHpmu7sZN4DKlnhdmu8mB4C1siUqoCVwMfRAsB4H6LsUUMZsRL/IAx6ZGTdKi
twJGzgpvW9DP28QuTcYJDukgQ/i176JpgX4OanMhHkxVCWxuY8nHaLyKTidkNxUiimr8Eig1xPNy
orpMWVzLenJYwnxxJkOA+UEslj/RZLSskkB4YsquGeDi69exFY7uyAYNGuRTVBcZ0UCZYdM+8ls0
Zqs89Ow0G+2Gqgt/sWEu0kYsHMz9P52bczutsavtE4ayQu1JghR2gvIT08VoZCWJrr2rc+1HjZXY
+OsUarXn0yi9+K6XoWpaPi2uckuIMA2WyiHnj7Ht84z7Q52dF14b5LhxzoRQTrF9Pgd1yV2imoMJ
UwXTCr8SASTXpNm+6XXtAC5c4qrQMH7XPxZegTcpGSDZ2zN7+hHBGpebnaDE7wWxnOEH8TS6YrGw
3gcfgHunaqYuYP1K90l65Yu/OaJVReGrXiNlZEreImDEXjpHRcr59HyCfgQJ9D8nwVL1BRD9n1kv
Db4tsRinysCjIM5sRUIh3/qXDt2XxGqHn0nz+wxrQ9C75zbDxRRKlMMf9d0fJtK9/vva3k4bGrP8
JgfVDXx+IH1UUeUPiXZViVPY9534FS+g2LvfsSVwpMdlouuHQ/bfJJ/8sciEbWIC0kz4AXG0n7hR
pP57qiDOk8hUpNl174QlIhoupi2PXHRoiuH1bqM2SqLYQtmycpojbJ8CLLIKJevgRdKu7X7YmroX
HOyBvZUx1xNIemzSp6JUcbW5PeMLQK2dxkUIoCY35LocLozikT1yxpvOQByp6ENKvEu3yyJwsXkx
oep/23Sp4H79o+KKBexFLXgeMyO7IUo/HwHP97DSk578CzsM5C//uXKPk15Qk969mLfSAh3E4A0N
/t5Ke0UWoGlvbtk8qkE5iAWWiHS069fNObzO3VCJIAFx8c0nV5okcW8UOOPkgkaMOSxY4HZT8mI3
MtgRdc0jo7nuYM2HvZrsrw52qlw0Z7+e45roSUBDuEwJOii6rfviHPVOB/HD6Z6XbKnq8VSTHHhv
yKEV10bpEW6Rr/HaFUOdjuDWCQofY3VaLXXBiMX2qKsLEcdZmyFebSESrkq4RLa/PcE/mEryZ8BK
kBcHe8Q0Uk+8/jnAKAKPHLkP8AT2nS5Lhl+KmNln6CW6ojbzL0CMbYh6qcubC43+m6RdPDeVBObj
bhtEb8f8V6brfJzjO+4MLL3yH2MvZ+Mz/XzlDWB9DiVfyDUpdjIeEWBonGfsjcWUzGq+dzqllwxF
1U3tcBzdngutJNQufTVisk5vcDKCBeBwU3/sYrcweSL8YUyfqevngvbcqENG0eawZ2y+ofodArsS
HiddOeMoZ+/SKmj25YOizFpWdDWjFwM5vYT/E58Ff/yf8VBDl8jLhJUtkdKHduLfusjpH5PU5Hek
IQP/OC3nNxeDHPHs2FZjiFFG+jklcbPH73e6g7+ythypvgeMoIUK3BcmgjzJmprnTn/pcXNshtHK
CX5+m+S/Jo2ccy+NzjJAAk6bKZ337ZYxPkyjOkMn9Zw2tIEeclyFkwjSQkff8a5Y5akAzXjw6Sf/
qGUFp8SE6aPZ3uF/t8LoazLQXLCzDg8+oHvxDOKS/PPFWe3usNIdCr97Q+hx/Gx4j7jOmVBqfbqA
HKjk9gkXAho++BRGIgN83ko68a1+oA5Bc2lYcmOSljyhSTQ6jxu+8PS+OaJ3bmv68v3F9x76hj/u
TuVEzsL+gYyaTmI1RvZajWvxyhl/SnRjlgcip292DzHt5wCHfESMf9IeRGSK6FXe8cXcpWPBMaT/
H746mzsjISZrvcCuGe44ky5DQ/5M7L41MBToHxM/kvZYWRyN6Tfk90Ahb5MFLx1zwqpmlMSQ3IHL
7cGIh08gDYsqIIc78vZTmd7oU9sNazbQ6zfMWuRHDt9IOBnBG6dTjbVCR/NM1UPAjC1f6EAkIaK+
SGwkWoEauHyiJMMhJfddqPdsn43EiEpLJHoHQtACzM+65GoNOncNtu4GPg+aywW1fUC+6fSGZFKi
2zhq8SmQx0VJWbHdQPVMW3KVLrTxbvkew7a7N2DWHpDiagPOf7ZbARL63yeJYqWw+YcAjFPosQTg
hQUkbysk9BZdRT0elJOyB2EY+RNhrt3N3jVE8atnrikfXgqlz5TJfLDCRXtSb+ygN/9O98ScPaTA
A4y/Yjgg/V7perWs3YMXW4mCn5sAbJ0P0C+AWwpq/DYsAXAeuJkCV4OSC7uZ1kIIl7KXBozDo8C4
QjQTnSN1jiAcGHGVMSQ5vke+HfazBqC4/ZJPBATcMjWYwslt3EiHE9fMukU9br7FYgFB8jfX6n8l
MfP0oLNYMyaDdvHO+EvkdS2EzBAXEUZMizjCrWBovgw13BIhx4eXFIQf+srvCBVaiw7QQZEiyCm1
1IOyf+c3LBbOYiqur2Q4W18E+ww+9H4cYJjF7IxADWs3cBl6VYeWq8CDceICv4bsKl/3aVdXfWvZ
SgQmGcdCQGLQ1OohpSeC576YrzpDdCJVZhuRvAj4VS9wjeq3vz9DN5yjJokPxoivWWCY4NCvbVVg
prJ3RKCRdpxqYAtCwzb/yYajoTODrtJ8lfnnWYLAEmWzwPX4ncQQMs8pbHU2NdnoB316yh2Iu2us
ak1FjscM/DiMQduHN42j5QVjRcPIIIzVEER1aNVxAF2TK6NsFYdTDclm7DyPHQGB1qhesk4xW8s/
AQqt4Ib4ii9XekQ3Vs26PaZZ5Y3jKY+XDMWjAX+VdV7FOMnXzIqz2XuD8BI/gUBAuTiLYUq6AFy4
kUuyNX/q6xcPasB64rCJ114/GdHam8gbHFYYjLBF6PWofDe6gIdNoUqsWjf5nrzo1ieECBv4ojrg
OlB9z3AIKUSr0dKnjEBEn6ZiH7SR5LkBRjspC8jE/fZL5Q97r1i20Rv0CxVFJPHP84/ABxSS+0pd
DkNn5rqXbWLm+aXxc0TN7O49WSiJN3nnCjerhpNpzlTeTBj0BL4CRRolC/uGh/aWR+84kq5xJVFM
sfNYRlT00seKL75PrY0BsI/GEKkAlVxiky5UgvHmffxjbRnJ4gnQ/ZrT1KomPV8exBcEmjYI4lvx
taCkNPmJJUwU0EdGY1j44GZVH0sfUQuOR1bbmupXApKcC5M5w58RTVREbS3fsZeHISvNDI+AgSwZ
GUNPihGjAjGLVNTElyDKHlL68pNx+3VX3b0HZZ2+NdsLbXnqR+GS+sYT8FNL902NmZRrIGtMkiBo
cWbHce9967WtPbCVUZgWnpKg7kYW6afqMcx90e54O+d4vuDlJ1RdYXFmKmlsvDY5YNJrzqGs4Gfk
ZwWyfxPFd0lX+gxDsjLMulXPXfw/aovu+zis/6ak6cqy7kwEdBXHRlzrZP5SURYICITOq+hj1GJx
FFhkLXGhUvrjYcpwiEI/j1p2D9Ooq3tkhmqgo3Bfu1w95i8jonjKlvRDbD3UQg9irZyqxkEo78aM
d02BTxJqQSEQst4ax3m2RQ4k4kINB9CtO7wXMOlRmSjfZB3xHN3T+7lzZCrkXYE1rdo/5o5w2eco
xhptYtKiR6D3PhmiNwYB3FI7f2waQ6OBLGTwehcqKYmLzjNDzKXkEepNWxfxTlrBXtGBDVaFBbbJ
ldF5WIUS0yIKVvKw2JauhxopOchVmucx7vS2NAOu+ukj3OzbzCAatQvKyL78xCWRLp51I/oXb2lI
cL5QZY/dRXNM5jLgyJQaDBGxS0v0TiMNL7tP6M6o/jntv3i8Y7v7uesfENWgm4Si7AaYOCE+giJx
wMKd6E/m55LG1Da/H0cNnj5hBG+HCdICQE5vZZ0LHSojGIwL4bmzpCuwD7hkkrxl9Jm+e3Ahcir+
mny/FW3xrTaq+atVS7m6K2DX4GlFkSPv5lnzcZcOQwUbQhA/6/TlCAsO1WoLw//f4lKwXvd5QLsw
vl0TdZMR0TxHAoruw92Yq7ysUg952zLPopUkAu+cz4yzgSsMxLbU0IwuDdpYUAnNIT/1h7gytliL
23dcBZ48g1C5PCOZeTG0LZIcMsSridl10qSF2zHffPmRk7mnraJYIMQn7aNw7emdvCHjKRZuGN7X
QmJuYYdG42SArfxO3XAZBp3RI0OjgUcsmumRDcNbjHOqHP9TmRD3VMAjZbl6S2CHmk8U5heC9Elw
dF9EMt4+EhM8a7Jch0itoj1sjeOQMr0DXPLVhDpSy3URozgyGQPch1uOqOR6QwdMuoyQxqeQ1DTr
3fJ10+bZjMrrm4fGx2SuMc4bTdvChAxSrKGjeS7k+HSdBSDwSeclmSwlYwT580JDFBCcigl2RVEk
JMDHmm/ZAhuWwduxmB0gou5cVFPZynTb34VxmA1QxfmFkUmcDVZnkESGjLjNVRIdKP+jQCT1X5ct
skWFeERMH3O3Ko6eMBqQjIZXT7rJ/q2RguSRe4w7mRSLvtjKqPXO8iqj2gu0sEeyV/B4AzaWqcRH
3AHvl9qq9gNH3GIxB25iuYSmmax9I0BmsyQVfdYz22JcalFfRXhlJYFAs2PuALXMPbvZ6Si9P9DE
jHPVBDjUwIhxqZ4IPcdh/qynU5pqQNlm/Br4I8CEAm1nZcYlpCofOGJaMXlWgsLf1VUvRQU4i+qQ
88fZcuOI5RwRJjcSaKtYvHh3BYqWtTsKeff9viQYZJOGDoD898B0eW0eOaw2zTD0nJQ7lPdOjyaH
/G4Y3+aYMIB1c56nUDEPMkVZaSZDm5/+fpBj7mUiQCd9pdjuIiq1uWXJMi3GLus+T6zP2bgURtB8
6EFBqJ7p4KIN9nizaBp/GkwHSeFBN7mfzFvVY4VYSUYJwPNRckOL8/iEAkA1x0VhmeoTG8APWc4l
LIMegS5lZnJiwQX50Y8AU0JB+m0RhyzQWJlh1j44huDgpVxTeFKQQoa0HM+a5Lmm7P+hN00O0m7P
oT5atfZKzTp7PMBzGK0jJ8Z5nL54od0EUCGADZorLd7XOtq5WB6fm6qwyaQE7cY2DPPc/W+gtc9b
rZcDiqKDp+FwU3dVwGyFurTi+Y7f9nflO/yK/DgMcQ4eogEbuopkY0/b8pcvI+BQwG4mz3atAV1R
Q/dj4RkYTkT8WTLn1cQcwafEaIRPSICmzYBdzGUmfHPiyR63WdoJdrvYB/QDO02q5b1yZY1jjaPw
1wdEWjlTQ5NIHF6z+8uK7o9XVuzTmZxmtwkapxDCNORMIcEguJU20PIFIsZDTTH3Pn3j4XBNu8E9
RWsWoA8PS82kC7vOT5RjVlcnmcO6aTzBeaonhjoHMCiKWvrnP90amd1eQbTcH2G4+WQvTwbeRd4F
IYS4aUhqhMwxZRyCyGpRzGY9XlRNWd80qvJzvucoZxi9ONt/8Hs7V+5zDxsu/8fZLd8vHGSuAwWX
kPfDjGnwOgpi9wdp+RCEd72Kd5WStKmG2/IEkLz/PcZZp6vqiz+2DIIXtjajr2P22OrDhjm6ttaZ
pQXZgIlmlvvj5iYKYT15Jpc6zTIgjvLz6FcIyBK5oeN89UIEEEY0ox2dl3KZgWXuAE1b9LYgoPQe
6I4ijjDR52KIDZqSuQmdFSxuH/xhZNDsMofEtfiVaVOcBn07rhFs7ch7SXQ8WylELZSZrK+Ce64r
vkhb+1pQrHE5nqXI28sRl8S3+InrJImTj6W0UaYoZPsGCuWFzBsV37epBNCjgsbHcXf1upApZUhC
Ig/Pnh6Xdo5m/OOLCiRII0y5Pm2INNsrE734qfQrgclDtpsT5MxCurshEWgiB8Wtjc3Y7ZOMHcmG
Nr9+4/Vb3xn4qHQ6iL7FaBD0Ltyp4GtVJ1E6aKoHnblbFxeLn/EW3aakRvAGZzr9OxYwUYABmDrw
ldOdwv5qaJepEJHPyoA2mPpPa0FZ5+41Vgev67e8LREYDfGTpHdag6VSAhARk0kmvbfDH7S4raFs
r4z9I1B7a69aRUCoJ9vItbPiQi+TX/vbmpTpRQBkerNwl70m6IlIP3cHjnaMD95FZrBv6GR+ilAq
SXmMhCTd1aJpCECmUadT3p7BM5WbuRKK2OXtU003GkxMxOXL8SeCn88By4hqfR95AaBZzAw5I8lG
DfUiWIs8tMuhXIow/FesPVJ0PaR13ckkHKTShH1hJzx1787AErV9Y6PtVoHlpfdb35uPVPbDWGty
xwZcD+RMcETH54bur9PbV5IbzOgyJmuMAPLovRTCE3cGJcrk2MnKD6Ls4kbT9wWukz6QjNJuzFj/
XBLt5iSFeF4CgpmhYBV8KmqHpJsc/qp2X+SZAJNANL5Ied3kX/XX7P7dfVGmqSpBgfyLyIpU3bJ7
r6wXghCGJ6C2dgi2wP6wb73CaRhfkhIWFrmQNKnMBoeSIQYAVzG30Zw+wSCoOHQgCqpu/XAhanLw
DCCjcUoXzIrrP5cjDv0Kpyl3gqEK5O++BAkm4Fvha8PtAJPcGanj7tV9f3fGJvEqgRGEjHhKsQpm
fsNCHOwOTdR3sl3B6I5dMJH1Ij6vBfzyrfyA5FmSvPAWG+7kvpcX8CZC6sBGyaG/boLK3mu7hYO7
00jy/smtu6k3asLj20+leHI1Gv3ze8oT5l+P3lG4ecXZyeTCWvt+FtoDdU2JXLEbPB2T9Dj5Rgi1
vbGu9F0y7KGtPZl3gexNVoRjMF6WRfGrGHJFDyR0uJrtA6qEpRhsd+1d3ae9Pyph3UxZ6DBB8D9Y
VaJz/xNTxdWWwLdWidj1fuINv7AZePuouuE1BwGubOatAKpLYAtq3G2ZiCsmqVbN+gYz3LJOvYNU
YQ2xJQeRAkLIGMal8uk+9nrhG9OYwg3K2jS7C8owF8THREmdd1EMexak6OMEVhp74ioYq0LgH57T
6rStZ48y9Jq6sZh17Bxg4CVS1cmt58JV2uOr+JtFsn5QZhPw0VMbGVEJ0TY7pHYoLC6BcOrbQQEs
8TKW1TrFAsOjUJscCNErzyM+HqGi1Bk8QbyLMkol4WqbhvlFTqKuPd624ps62G/SiE+JekgH1Jw/
mPU6gVgGmXMXX5CghPGUOWrGfyZJHXCZGuEDyZ1OjTJPbk0Jn/0M/0MpYEW5W6x4HSykxyAhKL9k
25WcuMuneVyFoJyZfECjjwvNFhheMG47XLGHI3653QMM9VdRN4EWXOySc+pWL3oo/avOP8xpYKPc
//HIUPRYAaCcQd4doVja97+6LsY32yCDVx41veJVMCPSdU/lDFVESyyXYFl9KsUmD/0rt32UNr0x
th4boK43lJSXwIO2uc954jskj78id0Pdc1he98AQT2FaKWXRoriCAesKusMi14JQnlBYNis3UgRW
HGWXsFO29QqBugOsrf+ZZ7t56RRpravkSflnOHjo/C/6w318/mSk2k8Dddv26cCegdED4zeROdNT
Ollj6sBRSXoZ7JeX7M3ETMYpWINrAtZMT1vrACpqd6h+dXQG1zFn/llPTnQ2OQ8PbHH0nrzcHnkO
q7i3WfflKcVjoFVhVjMrJbdKtq8HRvcpZEgoal/WOEETHTvfd3r4CaDCTgutNlff9i6U/1PHRn7a
E1V/APXb2zbx3tHBT7HRbYIkT8dQ4KLRHGpoHKTGdAnLgzHN5EReVgThmBFgEuafTT1cgF4qqd6I
GopwT8aHFr1S+w3H8Y3wDjluSP7VyYJlt3n+cM6yKc/8G3V9k6Qe9iJ+EyV+S5b5aAw2n12PlH63
7CH2DCABeWHKxa0OtTeUJfcRue6uBHJhlHZ9D1gdZSL9JszDyKT7xqhiQcxwZ0csE+UjbSdnzmg9
14DRWnAWvYgZGuXgMeRihmTvcvYB2UOE5pc07ov6ltWHdkj6QP6oVVEFhY9LIiKt2QAyDzuvg1pH
G/T/iEqbipA+MxYpRV3eDcuqgPkkRWmb8ryGT26BMCJjnK4lysVSiHep2iYVrnWLFs6oWkjpvXAZ
C8Cgwu3iDO1at/tqNZdnCtk7mJTGDotsz91RY3zjGfDzh877JsoyZ/4qv/my3OSIz0YPKIYG+WT/
DmIU3CBvB/PD5bdn48HLaXNlk2vxRUpB/mEFLaP7DV6o9AQTQntxsccyeoYgEzEdEL58Fjwcm7x4
brhOe12iyCMvKYAcdcHAp6TM8J4FijW36Q0jDL6m053vylsjNwUPGEmvd4c6ngIHA32KuBXOsP0f
Yp4Gu/LXnMWSlhu0MeVOfvOXUWo8CMyaphSosxdE02FfZh+nS40ff4MNrzVmM4gen7IKF/ruKkK9
Qvv7XhSO04vyfBeERTIDgSbautEvs/+rIILEMX6spCeixH8+Qe1HEOe1PexPFmt0nzGJlmcBwYcd
YgK07lfFNXCx28XNnj4M2pmhDUBPbnaP0Bt17HgnmTZWaHILeDm1xxgl2LwDKVQfSLLq6Biy645V
O1GdIehcgwmW6vLtE7DcAyXcpUILKX92rlblSNrrX5hunqrx4t9aaRQcrZ2kllzS8Gp/odDWPA4L
dH3bO33Cs0+s1acWCOsb9enmLR1+IW6Yll9babHKpNuxQ4nYoHwaVF328ec70kPziawOP80AHpWb
2qlCB4vL1UXuwn+uZiCK69EkkMItkN8/Vz3Vs+1eZVwatrLe3Mo/bmmNhig9lr5UFtTmW2tqORZE
yaenHoF31qaEpLrupCMNM5DUW92XH0gbktye2ENaXldRZxPl4DShWwf814VZxqB61vsaWbJfUvHI
NsKxTNxIWrVNGaQKGJSs6T/1VFLUy4IdQsKb/s6AKWQZVld7A9Gs7jhBIRdF43gPHL892uw5vT8e
B9p+WM/nPBEDiSqgHpPSz8NjM1DGnEusZMDUe2MxEIEhjML21u3s0PmYD3o9XPa8KC5sfHzZU1bh
LpGb3fU66MHbA7WNsNP20zqqjXf73pRBrPNKR9wTSDUkiad6abv5JuYAfgdnLyeUbgCHz3UiIAlE
HPv+5w2ZqkTETP3v2wN+ENRu7FYPu2Z4CW4zYC8o3QgrDPkEVl3w9hVPiDQWIbz4o3hvABgR36nx
Asmo/86FrHxk0l5i8D+x+lQOlxn+2wDmA7+oYo0NBE0M/uLFsUV2dUrHFB82xdcWA7dEOnpxeNq7
8OEVptGA/4x1JFlF+0CFfShqjsfKZ1AbXfVY7oOu9XfE/Y0uksvfeIFl34962f2c0GbYRyKAtzxy
2BJ4/b3t0wbW+xwrE0Jnk14b6v2kKrI/ZVv2yjWLA4UaOgb5OJQ/ZGE3SpN0V6Yng97g3Fap4SCU
HNTSHE6FbRexfma5qtKKlcfiidzyg4eidb4uCZZJ3lr1PgEI7KCsvTmCVGQpBsYu4qV2mipAjj6O
u/Qmkjta+zCo2ZpTqP/q8LMkp6/DK4XzEp6vSKnLmOa/hul2OndUqtiRJuUVrIWr7MBGm9m4Ypkp
vYT9bAo7mn0RxIklTWTR8OEIt4uomHCOiLqM9FY7k2qlqkNwLl+EmKQ6EbgBikZ74tgTMpEnJWl/
OhilG0a5qGT1Um7bGjgRFa5TFxN/zjRfnWCBZLs0oPFlonOGMNfgpL8hGjBJteqCrEeWFFfxuyPL
PCjbiIghJX6tbkTWyShU/50iufCex8tr6kse3IndVWoPzwskAF6t1hsPcenG6BWWfzrjHRQIHblz
oju21ZMyUDV+LmDQ4CztTJK1yS8zcp7KqDY0De1+FJhuSrFXOLmuducPy99OAZWzimcIFvjMB58W
Cg/cUkRXsHqX3dlfl2Ts0hIHmyjzbHeUoTVReoL0lj5LS20kqpybTf4CPv4nDVjzyiucUrItVEsB
Mo7kCsu2A81YTJXtnGemUJH5yaab8W7gSCY12dJWwn1dZr75ZSK7VIqMN5LWo3NJL4lb8ueMKhrq
nNP24EMn9xdMoxxPWlaZyKy9cWDhRsuO6SiYlxAaroxAavka8Ul6SzmamW2Xiqer6KaaLPVgsEX3
6spdclfMSpoNafIYYEof7ZXf2Gz0dn0ysFz9QgLlY/m0K3gHDz7P1XD+Q+C29YNH+O9jgrKEAgEx
jMZ/wx4WeQu6SXFYYKaQEYb2YMhsOabC4/S7zHD1meFl6195AHy4MXO2NDpzNhejD70AIoRWBiNE
Eeqwzm56ciXaZDf/vBF8nJEinl8oDUQL+ZKlE3r0rqpLHPSd1vOoQeCZN8jXWMf/xcYMHR3EHeLe
VZfG2kwXB5H0KaZwXAQmn0Y6RKoNHZ2BGwDA3llNimFtYnGUWZ7qivZjrOtguD+pnuMDiISy/7cp
B2h3KZHWRlDzaUFEtjmwoBARtwsrr0lMU34jAWISZrlWQN/p421ZxkYABYwzUraXoCVfAbDc+7ej
1gxhT84zvLzuTiqhSXGvuIvsPXWaMvW87Ci1zTx3dlCcQqqaPcu8l/6j/GgmKxLOV7S7/gf0YyE5
6GgfHxptGJTcoq/jnXvsKr1tna/zTEi64MwwF5sdSOP3Iz0RdMXC3jcQUN+hsSqEyXoYxZgMo+L5
sGdb8I5BJAjSQeHgmcfA02gCLbYMM6gVjZPUclHc4qenuReU14XQsdpa4rnudfv1yt7Nyfk2F8VH
uKnxXpsw1OE3aLWqvVKhSu99UMzSNXBRNxZNM+xP5HbEABJvzmVAQl2Gpf0XhO7mR+XB8xt7LLkX
O/zPOafYpNNBef+j+V+PA8QeEppTl7dFHJO81Bbn+O3vEKJ4hi8WKrRSiNfczRzdz4RE9uF+lf1I
uut9yIYytgDU1YF3tb/MWHIuMgABBKlQLwOwC33+tikHksF6FHJxgFozMZ6qp/MAnCCDbqDuK5MN
yQXsmo8W6wFLpEjIiMOhs4qxzON7+2z5MtUnVoqPHSZPAn7q2efULertcD9UOC1Wnim3TnL0LWTx
1iurM6qdsFAwUCoJiFLPJhK1iNVFn5cEwE0MIXTdqMYSvYpAgCKgRos70aSqiafDTrcercQ2E5/t
lIhN2VUYLbMkSh6eL8m8jy6FCx3hFKhC9lcjxDqPpFxOQrPopO9YeIkdL39O5d39xsfk4YIYZXUc
z0z+Hqp7TgGQgxp1DkmKD0lIueYOZMcpPWzE2JV+OlXDO0l5BWOux27kCxOhLWXEOdCAyG423WyU
azKGSA5wEeFzW2GZD1/TaOySf/zqnXH6fSLllOJssSpELdebuUJ+Qwh03ujCI4cHwxKZqatdvnl3
iWWFRBTo8aH2e2SnaPvavJxZej7OvZUAjRICs+IATVv5Lahbc6n5YJTAIpJqv++UBvoxKLBwnHs7
/9MjoY7Da9FvLGJ+xLb4XI/mL9G1Oyjt3uLpkIev55P4W/uhn2Hf2GmVcZZD5jAn773l8/9/nIVr
n2EG/I/tSMmZWJikZljMuuN9OFbwuZZwAX6dic8/0s7qnL+uIhFV9ihXj28F/2MMTWBqZnBe0vVH
CNSYaCLFzeGCXOMmpUrP8wFrkJ07YQGx1TJ51q2JBePlK/CIDfr4dKU7F6Wiv/WLA7v4oExjBHF7
XeO/WiDX0sblhmU3IEtRY2vca2wXCXP9//OnfR+cxOsMFcfxvP5QD04i5sDR/U03ksI1zbOjDqjQ
I1i/IDtUmV/PAUGOzEoqCLc3MRhfr1MmQ4w4QR6/2C0FRgS21yXAx7OdrA8/F6dYSoq+PyT1Wkh5
KcD4mSUEQSPiAzSwhpanIWWduOBpd0Dw8xSbwsvK2BI/Pkk8J3/dSj44TOt/2cZXNFW7AW+Our3/
TOI/9/lwDNdVAOYbmK4pmg8Us8FxID5MzmFA/3APXs/dKnQpuGxwlBAdgW2g2Sy9jsHjMWI28zzh
8xTbUjl8t4DdPaJUg7JiybHLVrvmmdp+EgtuQU4SVaGjUq+bqMGRy7yNIe2FDc0VJWlXCs4Iw5TG
mibjiI3dV18hua1GRAIu+2S6AYagswqnCS2iStZVfM8p3qKUmr5RcVGFM0B9TDkRThvIv9/oki7F
J5g6KrcA0lrn7+DJFnq38Rrkh6dNAzBJro+zn2EAMoMwmYHpqgohn+oJ06FvXjkpfQPd91iSu0uM
xcnq8jXU/3NDVvNs7nLXAuMIvEphWSOwyDBi5kwxDfbiDaNa7bc/KRPcp23w94F1Y0H5bN8Fj1k6
x2uDj0nAulRWkohxEjcY275ebJnISIampzFFpjPtuPRG+Nbo3wHPhc3Qg0LW9b31nu8XBW6Wb/JM
6Xed0jtt8HURGh3lqe7BA7Q3FZnBRTi9iZ4MSp1R+8QW+UQRB4tLHMcxtuzP3kqF1/tWB8PJuIKC
ExaZHE4PPCbgOjM7OOpHCP1XatyPt3nLwlWbmN2/GAEp+iOoVWxvQ0qXXFEjMoviXvfZXlQtaktQ
MWlTdA+VTkqLWScG/OkpcufY+ld/JXJuvY2JHB8Zbxaep4v/cmxURfHUkky0KdOTmZME6FLmS1Dv
HJMbVnDEcHsGaDhwAG8UaZLkp1d2Aj6QMDrI5AjhmE3EFBSRuQnxLmpZ/Aap6pThhFxLZ85YyzFn
powBcRUuWeqJMVBgW5mgg0pw1ZVi6Vo72ShUr8GgaRpre7YjZ4KhvHelW9H74p2g2Xi4oIqeZZvL
mVlNLn2QONfTaLB1EjFRCV88TZ2QUWi/xQr+wUXCUbSqubLLBWvA8gvvggChykSeV3zDpSfFyWrM
70LKcXY2AZKDFC/FNXT5uTtjOYSIrjyg6TiUo/dlTpTRSja6SE1ei/YSKEcsSwpTgs2ExG7vQFwd
XadiicG/EkXrHRilz4yQOn2y8dSAKk4e8Oyi3IIMgYEskAHqV+hPWn0DAmeSS0hYbx0P0IfhzR7X
aFWhubpy+A4NJS028mShUsD1uwzIUELyndbGLorrJsyjSYpAprbWucGEBXke4qzsCORw+Pcqy4Ub
3YIof6I1541J04Oxm4IhzFGZyBRGKWgfnWQ2jm3VwnCukhzqsuxdMsAvEjg/cFy2zZiQfxvmNgwe
NPUeXC4DNRpJc7fQdvRfd5u2697YYU6Ix6Kn+abHIgwlDRtJxHkW50a3RqgDTXaL5b8run6RpqAS
Vmae9Iwch2Do+B+V2j9lT088IvALQP01G5roJJiSlMLqaEJAMJ4Y0ewm3r0TdhNhZkxcZ+R/mQs5
rb1qVdsC5q24jDsjQW+mnr0evjaWOyECu5wzMmVvs1B91GHR4X5e2do1CJI6t/fDEVt315JtM13m
Tu4A29SI68fwYTyCFrYbHhqONL7XOntkYVKMosbIshAyjeLy5UZwF+Y1rzqonpIpq39vG0NyaYbI
GOC5jvy80T4xalKMv9z8bw3kzym2f2PZhuqb4ORiN00m7O+NpyL0znK30EH2blCLSLd61XmMrOa8
ZxvMlVeSWjRDUMSAfzm2IadI0CGBFuYaASauZoJjwvSSsCxSe6IbLMTN8/uUhPPhnJOCNkH4B2ai
83QhjeXut+hAOeoM6qvv4vz05EH+myqPvhB+JnjZEaC37KMluxavoQa/ub/6dM7qAdiB3YepmKiZ
feGm0h+e4WmYGZt9NV1iazmvpezoPP9gifvyRZIB9KNpXUXsCJyz1+T4u8f82fIXwTk+fSWp7XHE
8vEUeBErGZpy/nG8drxixESi3xc123mk7WcKdRJkQB9oqSmCWWz6Axve1/Epbf0KoMcPesiZMQ7T
akcZtrWn6X968KVsS58yLowBd6JsDkgTal1KiX1lcXJxEsiyeZipOzmD3iWFEKKs2nTUow9h1AE6
qBPh/8x3RIbUFk96p27gviwrZmI0jZffDJ0vAnxTCkTyrYmPtrC0wsCxpcalq2EBDzjKv2L+4abK
bOS9klwlloLPVCtIITE4AKu1POotFVR+og7GuooThCqUGAyTSpgNxBKkcruTbqeNQBZv4an2jGui
ckDpbfzSrC4/9+H2wLXn3fR8CUrJRtIpUB8tvm6iUxBafGa0qRcW7F16Humn1uZZ92eGEA3A3ceQ
nC8sikkNOYM6GNYpLSWN7GYoSCSZwP2C6pMU4j1kONEABnw5CTE+NW4Aff9xu92/o4fcyrdyTSoK
M8fa3Ae5UbtJU1Co5KeIey/E9EldXtd7/Wx/TsBubVfNGKhbxnd3SbN42TZI4CxDr2axEW/HT9Ep
xrdSlkIRst5uMbKVI7fxE81QrJhtzM6U3xqN+/5Cwt4ovt9wpxziaC6EbwtAam+xeUDiTEFYA5ch
RBwo054TK2ibT82rThbT0bRaH6WQq0Mr3qejxa37INhHsqFMArX3vZfEfu/r7AvL7z7k02dS0ETM
2+mo1jQ6uAws7v4YElWWf0YYKaY4OpSwIdzuUstduBxqGzLFbSumijAEyl6jAgBAtpaLBNUIw5xm
24J/5nlbOx+y/SDm6Z7ki8rmFOOxOqXOjTTM/cy0m7ykrLdbSN2H3PmHFfAQo7nIrGtvjyLSIyO4
GaOwEQQE6Wz8Zq9K3VAaBVzDp2Yr5tgtR1WPWMQ/FTynB+tA5MSCii4ckjURiY5gLxlD3Dnvznu1
9zdm607qyed+e5Pu4qFp69nLqhK/194rJumbGKwRentyGDFIaeh/5N/BNNprwqVT8CPOBXSAu1fy
GzBnobW/UdqIiEZDhNtcjj3wQuSeeUQdArAoBCznPIjEEJdR5AY+fFopPfN+8P5f3Lp1WcpiAkso
T8Px6HeCYytaPyyrJ88J0sFZnvN3EBGbTW59Sci/7Sr9T/uxh4RS+RmWjz3UTOhS+13RanvPtdSp
Vry0akW6iiVuViIYxQ6qxWuNidE5H2fa8gyEfZo4uT8oJdnk01pUIvaWkj86+AUzxXbNopQCuQRC
VWGHslz1K1PPJegzd/DsRFrFf48S6TB0+fkbxjfuiDiL1skMi+CVeXEcVGsDYiM3yOapI+oEZkSK
Pzu6ctdxe3b9IaPxgQoFV8Hcr+M3oVltE00C+1xwrOcFHEqL6mPLXrvc+VBXf6FLhOu+fOqJF2ZU
R6Uy2GsKOB0DM6E41ERInKzhcWDeurFlADZnWjk3jMoP9l3GMJ2apX7oBsMSVbdEIUr4Qfm2I/yU
kKDujrzJG5Ba0Xk99Qj/6rXHxCimbVWecagmoeO48a0527eDBwUi1OgoMbTx1Zf1xvcZPuInIpzj
CtInGW/g6rnX5TLe5oh0Degd93LWRFprA7D5Z/vbMAuhoNU32sBvZOMmHC79lpVwzJopFTr/9Q+E
XvqHSgxPQJxowEGXVt6Q7flrAaK+8ANdLF0Yv9SLTIpUeVdSN9MjRIg6tACGP6yX+whlE37VcXxz
VXtbOzdhgUp3INKFhXJ6WWDTBjNcOytEcXmuXJEI6fHNM+XNHoL7tPej59U3y7f2M/166XrrfqLF
0ZZl+LRyvKiKovPIn3C9EjCKOtDQiPQki+yY10jVnmLvujs13J4/xLcT7S7n8XUPfazItc1NJ0+P
RXrNBCwax8VFOVkD+OjTREQmco3xQ/kqT2pjIFX+CPUQUX1sYmJjMI6mcXDJhg+qRkqtkydGf5JQ
ectcDiLAlHDqlzuRe6lOKV7vwuxJ8v6BTO8XRJtM53yOXVjx5gLdlxROgA9QvMRpoGZPnGYsr0XF
IA+6OqjPoQH8rdpShCZPz1YZri+yRJ16pBZ2UgIlv+3fuhSNOiA2W5aZkFFIc8UQWGYn9nQG9G4D
sZV9ndX2EAa/nsELX+1rP9t2uwK7bN5G7fewx5hmgNZ+jnoIHt4J+ZVQ2aWfWxLkKEEkDaZFb5rM
EGNmpPrSzbgebVPOVpzys0+QSoNrszLJZ6HmPmwd8fHsMUa2y7bKEdYLAQ3NVblnS1f/LJ/x9OR+
VWm/QCXlieWWv8ma2bs8ZPukXP3P8Kw/ZeGGQchyX1X3xyxxDstKoi6Y87qmL6fIlTwsTcD+SXR1
4cKHioyRLhrx1fwYl8FPeuA7m811wgclo3zQ3PMveou7k1g6y9o/NbQs4KlKOgRVI/BusqWB2PRf
eB/A5GhB5NQAOusbk5IyFP+hDaGOfIG22cum6zqERR8ukoJ3y0D+73CzA15laUMS2goMpAZJyH9W
ud+27LPmX3MxdmHbGBmlqsOou+EvjGrfEjkHlubp4O7XxSn0g2NSXu5tlY8l8BqGn0gMTpjkCeTb
RBSqf1JsmkEW+13tgrlIpoh2E/OeEHQHRolh+iDwFvLs2ljBMIPQfa15KROb2QgNVJswZyz5l1cB
SLmeC8j9EDIhBfElsF3oLAdvx1JT4bVSNVVMi9vlR1/FUDIGmxe9mtVkARrfFA9OKOjmiGOc9oC5
9YGJs4iP1iwJx9fEtCi4I/0Hky4+qB6IXynK5WKlA0pg+e7G+aVRzmZMMAKKVwrVImlz/Sda5IEp
R9FXxaNszzbjiRQ0ERmU6SPLbyuBgbjmkgm325grgCgvkis8Xj1MZxl+rYt6H67X90iSjSHNXiq2
uMe5X4JaIiOzUL597EjbiE0sIG8eUQg8thZvl2lEa5wTMmT4VhD0YmxESzVnnbCm/BO4fF6mzdyu
XA+n6fG7T9UOYvy16xoaIPR+dcfLApaEFsa8Iox7ehek6vahpUWDwLwTfHngcjgHv/jvdjDPvz9d
wsy5DvViKzqcK5+r0P85rCahXerywKEyhOkb0ZYCStCe8FWMFW7HgNzlhFnclOE6e/sJj98r78pZ
ZZfOpBhP7zySWJtCIiiYwECrUyCs4XA8VAdjmyaebqedSh/hMu6ce9Tsf+6gKJh51PNaFnOrbOai
uDCvwHK0F5KkZ505p5Z1Ay9e9xWnPYcw7wKj9ao5Wq7lriZHYslKOHtbvHFWg4GXlI3WT+40cclx
DLwkZLkAis36vCE/YlmKN640RRqW6qRIUIPY3AAixBM1JNsaeJdvTcRv6D09L6POdY81RXqJj4g3
kd+HzCJip8pQVbbgXCwcDzQ9/UBJ7Wcbd+z+7s/XSiiepsB1Zj2vuQkYh7k0T0JXe2SvZkc8BFW2
IgT3k6Nymuo2sxfeDNf55o3IXy5uAZlOVj8dO4j6aYg72YHCcqc/bXt9eBlFLaxOT571AXdV7Ic4
/x9db1NpxguSC1eciNJ27lXrMM72Lyc+RmgbUcf1pwZdEfWZnFjuaSfrLX5Xrnp3qHpUk6FsLhQv
+8qfM8GmdNAMotT2OoyZMr5Shal1Dix/r3G3dTWAYaBzDJl0uFUA0BW2OaUXtdBJ4T4cW/WYLHH8
tnwvFTpfXTfHUBcPyFYKXkGiACwdTCRMIEwVC9TlMq3bNo37WxDDDh+5KYS4/IGkATkICjM0ktjt
00PiArUCF0EhikEL3P5ZyamWuyg24JiKBqf4OVHKGQS8XW+laJ+2QpWUbA5/sqtRWBYgto2VOQRM
ctMZKAkw5ky/YMh5b/c8bASIYOmql4MQ98XZrIGvPX8xw0cLtQXw88uOUPkdabFJdpZXccgpAegZ
YQYDt+vEVpPusLJqKM46Y5vJUxeTj1rPujOKRWVgQmpIOEiUqjYa1eofOyMIuGjAp/t3i4lK0poZ
PZvYQt1m8Fw7djj3eEgAFjlvX25wo0UmjV41Scu3e0eWBarXPK0sTdTl/IIMw3rw15m9kFqA8ZmX
aFSW5R8A7ttDOFL7cZehR3b4h+Bos0EOCmGSXyHfsh6QR5QPO4sf1AewoPk8tJ7M2BhA/E1XmS4v
HPP18NxhzecsAZc/zKXX/gCxMNKfq7YYE+agH46CXlvOZ7Tak4GVOoDOcnf7Ra4MCSkPcWGED74T
45XBs4vMWANkb3c+aNaDBs0QIupT4tD2IWUtZn/ODdJPXcHZnHIpLsSvDCVDodOryMR1cprAat1/
7FcP7ZDCG4q4kgnGeSSQbuGwGP77EkkVxz5oNGHRIu2c6JD5YOzUCazF/1QTC3i8FeuRugdKd3PH
Y1gmRWN4BCv3mGgph8zpWVHew2eUl6f6Xl9biCbaJ8Cpwc6ZCMGa6infOfM96rPtFdjBEXAFwGOU
npLJibHAEP5EOESFPSJKpwxnWq3ywX6EdRVXBjRty8qvzvZd49XXS51yHNNXg/5Szy9VwnDm2LDd
+z9LOrNqLf6PS1ZkMFqFuvuV0dbJZ/sSjjtVJaKb6/v0Yf28ontdJDwXbVWeaWaSnYFv6nhoCJRz
oo40GK/5vrYRjVoFbfC3P0J2BmaoqfNyuUbt9YqExFZ4xE9jvq+yd58lfHXPTR8Z0dnUqYbLUwd8
nat+nzkbbEAqWeRieXHA3gumkSi1XmzY1GkDDOW8E3/77QsW+vt0dnvRKIN/+FrcnXIsf9DX/Iby
cVVAOE6cPUfrFhQs4QvmwVUymYrKLgLwUtRxqCZtuycm0RuldSvhJpqsG++ceLRrfITbioxlrAhm
3DhEJ+UEhS1k56SRS6WhnV4sFGWuSxenNi/YVsxe4qRrYa1dY8OdZRqxz+UQqmr5ZH4A1A0/Tm6q
DIWmySEi+2qUwcvfHEh5yq3IpQVeiyGNH1VASQRqeu30cmxyfZZmD3dvDYFArxc1LXHUiDXT+bMR
sBdGwtKCCmFKz0Rk5Zq3BOeRk2DjxLY/dlfml6dy4YTUotMcNYAKkIXXuOQEkxftYUaH0uhUfkIJ
CKdsHwsPyJ/UGZizbge/BT3MMJvAqmkFGL/zGHAM2kElxndf0+WawHD3Ui7wg5KnBlc8fnv9XgZ5
U1Jk0/YH5IyiYUfhAV3IHkqkAABZ7BWVjvPO++mNQeq+8DW92dd2BswWfwnh1+GDyv/h9HQGobTq
d82qRtShxTjDrlLpFgly+vPTVaqmXr52lnaFLjnrsRddG6jLsc8yy48yVF3B7QwwJ7pxr0E7BykS
SHtI2c1X+EzBYB2DGGQcTwW1En0snxMQESTB4jyJmMXqHNOo37EZXwkHGrZh2EWLUO4Avyv3+Cgc
h+XvgEoYpI9yqiVESW3m0yN6/oCgYCwZvykx7WFdqsC2348uqLEVk+BOT0B8PDCmoutVEaN4queu
WLMsTp4ncyQIGaVkQITN6GZ5j6jpey+SJStmT5aMUg4RyAFQdBofRSNleGCiGGMPqwVWX3riFdK/
NtPBCV3I6FPgCCNxOX5nuNHLuiGgWHScOXGUn/Hgqwa/pdWdeUrgcZdMuc+VcMniQWavI3E0uyrB
Aoc4IEC2Dl7G3uD0qs3rbq7eqaouHIW7Wm7CYATV1Gy0opxd4nxyP9/Idrq/9ul4bo5zz1ClVvDd
EEaEc0Kzq+NuqeVzvwGmaV+85jMcaoQezMfoIHlBNcuWRLKQ1lvsyzewdAHXl5uHrBkcJGLb6Zsc
Rt00ZRZCZwYU65ijr23XNO3/Hoyt4/T5x/9hPgOUOzzKwYu5RBWgKWYekJwF/g0Gvt7b201y8EJk
SjSfFSCQ+/bWyou6Mc98jWDm2y/Q04o0uNk4h/SAKsYSsHsx6pOcgtINRbCb1Mdi2tgK4S/IpIXw
Fows6Npfj6HxArswaFJzJYlCaqP2eRvmsfpunhKQjwoXCGoqhBuwHqgthu7bRviVWOaUovq+LfRz
0OhtCfTx+ZMLkrqgeh7ujKJS30PZTOAymOlLXdTebaxc9Fipbg+EDOQdhinj9xoiKsKSFlJgVIiO
5ZdNXRKQhZowK6uFnHOGs6eKfweO73kut6DfVKymyndV9Bh8kOcZI2e6pVOP43wR+gAS+1bfu0kV
ya1QutAk+tc8WIGMts26aIAGfnwM5x+j+d+hd9R+UumSTSbFbaX8fx7fFm3TJ8D0SkkA8mO6t1t4
1go2sqMW3AaKWlCTFIJjc/kdb5M6s5vQD2XZ0jFOgVwgCikDjTXVYs+F8vmMsRjuczhuhtjBHdzX
vbeUV1/YFA5x/fs7seQwFO/YZyWMsarUag9w7vUpLQlrbdxb6ELjhWfnKnmXu5YiURO/tYa99JQJ
gHDOhIaIhyK1k9hdHFnBQGu8dX2ccjfhtdMg32O/iUNUzJOF0Sql70RQlp5qYhB3403yELH57IQf
dmDckJ3Lyug6c8al2gunYhyhe1VPZyrs+u5BO79dyS4gIg6dcVihFbmWZRhB/hhlbM9oHY4gVP3v
EiDKwdYHp25ScatdDcDo9c8xVZwd6qo0Cj3KUM8ksLOi7FsKMgjxFFrvn499IXWZtCDoZlMT4XOD
l28wjOSiFnIjKPgM5W90DkBPZU8SxB2EPwMQK8NyVD+V7gt7b4nsJe4gIhqplaeX94b5EUKGzf2M
rKBJPOwfFzDmnxp4a9xp/5q6TvNNwDL2mfmx4mzy44k07GgUQ8USULNVsfxDCJe/ay0w9MSbzYng
Ph3Zc8AkQU+aPwxMc2yQFTL5ZO2b7ZrUQ8V1fHjNaW+Ki8D7e93GgcCidavCGfdf+xxFnGqnVH82
614G5eBxFb8V96MCGdQf+IEq9hkH/e3PFlTxrvBgNGZu330EPHkj16MY8Y9DWU2vSb476dNv5YgP
0IaoVp7EFUWAO7iH9ohb8S96Kf8oC7OHbL6yVVtzfuOUkAP8VQ5SOYN2jSQOBuAlNVKdqVyvhwTV
x7tXekkj/eiTKvOpHnkpYLYlJuGPjyXIRlwsLq7Z5TDA2rcHifuWRhdcLaoCqB3xPWA/BM3eR1JI
1PoCq6wv6RFEHaKAvXjmm6AxacNoRyrF6i1COhYvix3YUl24zzZ3firFCbFdDJ27fEkf5ZLxEGNA
GBils30pZWUSAmpasKwRNvgGIQ1a+LaI4i3R3zTcQmhYDY/KT1CZ+xXgnDhuePMN8qiC44au8vSS
5aDYU1oUj9VtQ9MQPiqrlb4XqKcLi7YLAPf4GAiNko7bwHtcYIvzu+QD+W5wrkRoQTjP2sN0XI7K
mIIjeS3Rt6fZe38/1/n6+wmgFHE2Zj2TRo2zQDGUhk0uqXeCWG86f6RVGsM4XAm1pR5WbczG1r59
E+9x7d8Tr/gBUM3tVldU3hzV5VXiXFHP7W8zPE/tl7FEbHjR4GkB60/T5TkKTXqQTO7eV7Ru3o9i
G64yWMxF9BbkPYXkfgTxIEbWZXJzC+Fv8RI+ceeQ8xztO8D3t0EnK6oIW0YEkVO72qvL3GaG0Me7
vxo8jG+m9r7VCoyNffnBS7Zd2Tzr1c6ff48aSOAs4Id5CbjFio9e2d49XCPZd4FuiqZ8+tlxDBpd
lty5Z/UVay3KGxWi3nKl3iWHTw0OnirVYwEmoK++QspDIKrUlTEGRzp29D4uLS2GXXzE78YNyZml
ARk8DeRobHd9oN7y4HrM7taMnE9Wwu9NP27QUBYElctA3Vvl35Rej7YChh8+8RFBGUmAQc7SPI1A
vUqQwpbdCLB1uUn8o0WEC5RsEr5ceXYwgj+zVyz15W36Xi0p8du2uGxTXO9mOD0JgaIoKVCqwNSH
w1jIbmrGvk2PJT1JVkAUQ3ATYQXdsscZbNZ0oexiyA7twRIY1UJMoB1/Ryjk/qKZI3VC2rSBoC3A
blNi0V4hb7l2il5BPNuemBSeJNZsJbvruIHuOJpUUoIseDjU2sS2uOZotjnBdhjWZ2UFbbMoEH/I
XdGM7GyZFuKEAnSRFIJ4azbEtpGwVBGUUPebzDzablVAvkj7FIB6WKLUZXrgfO28D0Z4nDWfwWhT
v3dAblM1QjsJw8CDY6OkKlo8/snpZQ6uTtJ+Bxnl/6akxKMtknAEpTeHpkX/wZnKVsAvPqiWASrn
7XmYx1zGAsWCHR1YLwVae9SMk8yqeAR+VXvCyHwb0RneOca31LXeQuF9lbXCn8Bj8fQPbpdCpMHP
Kjb5PumYnzhbiYJn9WuaftOWSYiHlJcHE9StNiegww8imWjckqnejjV3fp5b/j8uokFjo+NSs4/V
P5RrBGW89KysUTUAqFCucKZEFHRbLIGzlOXNHt9njcQHXTDVfLkEKY+PVgHCvuPxDSvCQP2izv5e
gtRsNaObzEw76mxsbxg0xmHd4Ml8CHOrMT7dBGB9kgaCka8Tt9Zy4aDLC36mf5tydzPPpeNSO+1W
iLvhGEQKD48L5MKw4DtWAdP6epa7+onCwtaIJoHwsjpObN+1zFdU/P53+ErLZaEINhYKYTCsUTBa
zhcyaS1Op6Myr8uGVZcyOhqYhcaEaO33I6rzyeBaGewkOw/baX9Mx3hgiQhw/STrx+2KKok9DZs5
VM9+uOuO2Erb2RzPkdyp3MkcsSNcWi55Z75th1sc0C4d9M4UC8hte9Lw++rx+NT1kk4rE0HH2Mrx
WkBUaQIu4mwgXfSPkPpV5+egAPBoizGZIkSZ7ZjFdRYCNSK/SJbrcA30fXjvZ07Wcp4zAEIZkYJd
7iZjoecXd2E4iQK9n9/c5IrSlozewLUpx2InW+YjOdy/7MFe852t3+BdcDqG2Pn478oXsXc7RD7O
kpYfXa0lIm0UWcSCERQGePKT+OaLw0kGF/HJK/Jcre88uOgRlHqS4GpgWnX8a+PWv1IOr7DBhssv
S4IWazilAK7ssuKIUUDxkmyDI0rsRO8S4B0Akvut+qdYa0jMktQPK9CgztywfVIIUTTl7NZF8Sep
qgaTN/80RARc7oCX/iddABdshsGZ1TKt8LHq4SRIDht4ZSASOI5a4bwfeUN9VhOvs5camC80dPKr
bVJUia6kORS4A29sr3UZIOOZAS+xHaC+o3WpwQXN34xCB0YSKUBWABBn5ERLOd6hk8yGg4/DPzNG
q4zgHUy3MDmMxG7aRorb0S6+P+1I5lEdugLGUxOVVCFOZiGkp00lA+z57XCTxFbLTh6Qm6LBCw6F
tKMiKCm7IH9+/6D8AABSa1RqulIlb3/Njy/VeK4pEPpZtq2oeF7Oj9n8SHmzCOrE3GVIO2YGs8HI
zPyGXlyxUIoVaf3gZB7AfMh1SraEawPyy/7TMoFJsJy7d7lMsZOV9kzHjFx90N3o0SveWKJmuIsB
2lYNo4T9MtfRoyJFYWlbqRJ8lB0fyszGDqr+R8u9AmLwArFtAMEggqg/TXq/Jb0rtvbuJtRBUUs1
oN8LHvpKO8lFGC9eyhcZ6Z0cKiomUCa+8xITW1IjLlzzLSh0avag/XfjJvHb06hcJgvcGs63+KJo
WkuG/o99EVTN/qg7nB5kkLkCwobK54AcFaXSFindECk1V/7cmBhqCzZl4JYKufRcrXtQPc2/OkJG
d49DVZkOkNjVM8oJa2Bn7a64U7lxjXb6yBemM8xuxi3pH3/vxtCCbcs282fnjBfFjd9FMwAfsVlK
08Y8Col4LB84Jm/zh4GwIEIrYs/Ipq0yDzZTaYHPwCp3dCJru03b2klQ50vlYjF1r4zZtuW5cDJz
edC+9fdhdO3AfyrFBIBip49jlAWeS3Nh23h9HxMX22pEeeBPmsCjvSJd03roreOuIixRu3aCuI08
afo+GOVqIRJKs0vrBFjaFXrQYO9wZRRa6+DdHDKD/GaV3wdq6x3fpHSSo2l4mehgzcsaAE4E4yFd
zTPJGg/Sgltejod2bc3HajKV6BUgtQ4ExZCkUFJ+dqdtQuY2xGIZgyi5g+nithFfNZjZCCzwe3sL
bcj5FcDuOzZ/fK25pG4Yq8iaSbGl/0s7iDJKOIzPObCmmb2+wytO9RI2oD/hH7ScrR47k35bR25O
bg7r8DNcu30bbFJjTXtpuQd5J5uqH2NwKReq8JFPToK9O1h454RXF2NynO1T6x41kbJQTYx6CLuV
Z4EAWhJTOCz6z4oOuRkUvNnxmkTKiwU0y+y6ApDPs4+/JgUXfew4KTDcbB3k47ng/uXqIN+h/uyw
wqsRNTCmZkw4BoYebMwo8hKFBnzfqgCI6rhy41Ozl8zdrBORKOIEtwXrNWzLb1WWt0oTLnOWHbEV
j37sVXUqqgb2zaKJ5n+r+bWaaXt9WqxQNdzp6ktTyVgrj+R7LTQ6gyxKONC+d00pxq4VALoG3L/M
8/Lvt3m6mFGhAcflhwNbKNddjkbMdpbaSBnuLfWZo2pA5GrVPFnsnZMRHtEYMP+xu/i8yxEriwYn
h5Nb41AedoAz98rxwYVip/bUTS6GtJflMRPTq6QytmLJpeOoc4mlLhwvx4RJ8y9tFUFll/GNFSg0
lB4x2sCbbgbCcQwygyLGr3czUoBQoA+/sfqqzx0LNsObgfftmwqFQz1LY63PhCCl60X6abFNZprh
snzkPeT8KuERNdo64CZHaChGG8eKeB5+oV8F4SBDOi7gE4H11f0ybyTW3h9w4wHeTtnXJoWN7Bbq
tcf/3Src+hdmX+3DqMaiHH8h6Jc0WR7iC4YChoEMx6yRT2xyhC0MrOG6X1aE1kdpYljvxr5sXROS
McAejf6yX8WOerRppmE5vnz2GqEYEeJgTBpAY+HEheT01tI7QKS3qXp+SJSGuSKjeTHKq0ZKqTIn
blStdZ+ChDvFmNdKQ60gJeuVVb8kHv9ffrlchqqXqVW+Acm1jcvYhUN/lScP/0XnfgHIMfJxD2EH
ojyYMYDM49zHHVMLTzXguEMn9DH+W58zc9sNHrtc6tQtIF8oiPwzycI0UnmrMUZpH5HcteRoUhfu
uFW0jpK4CI5OdKQahZ4Io5XQZEwM1jZH/8bHqMn3yPAh8Oqwe259/QGcHBPgsi+EFdb9zR4Ug/Wd
8rvRpCoeOZ1ZdndwngzaUFIO6Y3C6kIAMhoSLrI+BtDvNOrGTKcNQWO+PCB70v0DYDz5ZZ2pFOqU
UM8GKTWdhBEv7law72DSTPkBQdrVPDd/uxR+5iBdF+K1LTFu03G9RpYfZIMCljpVBi2g6WmaF7eP
G4Ok9ycTPXe1TFVohWtMcAAFJOdy3GHj7wSV5mQgUU4BVWCsTryQ4wL20VMgVnfnUk8NfO8VF/U2
JzNaezLLBL6u5dnmgAanFIc9eb0kNHr1ygavsodB9QZPKSYWhO4SFp745f+bwNy0x74yd3DOMLnV
CAVcDtTAdF45B0nOWYdFxuBUiEMjoTgZKIjsGx41pRYBxRks74yowl4uqxn4AcKxIemZCknCmqEr
BtJO63/U7/N1NQsqZxDE8DpEqv6lZ7Sg0i3bVcHh+eQDyZG7h6+Z1cXw9bvGDnC9wTFDlA72XgHe
DWTxx7eO+ZcvTllTfQURMK/G28W1uPmkkE25M/8KjF1M7a+/3ibRAa0bgKlDeDSqMzI6RDEyzZQu
X6UnXOx++mQuldgzc0EwsCP7YbjiPKeihbdEyGQesVtVQ1RDec9bmGjlYTg53wjoXSD50pKmnrv/
OefdPnvHtH7VjeuUQC5bvcQJLebUnXJPQaoarU+duwJ6Cz3Ww/+6zuu2EBqAj/phaxjjqMMgkHUG
K5F8gJC34eFBUrdLQg1C5p3nmrpiwoxsnGOUqVurxrKNO2+78OO6oR8HMvuoQ7Ifr9ZvMstB7jKO
l/w8vN6O0d0ISeO/l2MwrgDXzBKxplH0JAJFQdAoY4Hz7H9Zo1Cgd7FUQWWpumQULHsDVKHg2aRi
YV+dBUBn9E1pBH0i2qfXcLsWqTom/HxzZYQwqfcCxIACRMaEwxXoJOe6onfAcqKgAn+vJBOUEFWG
Px7iC8a0yOLaGsOfYFJ44eSvZuIi8LulX2A4FaOsAwQuRA8MamfwkgQeFSiQvM3uyCSmHdcJ4jz2
wQZwBYatgZvH1hsmZLYIpGljGZjJORy5z9igGFnvppLX2UN1gzKlFoQ1wf7VktsmEEDEpto2e6W+
LQwUwzgwNr0vFNlk1cssGno8ThHmyEIQ/181CklbitdKeMU8rA21XBe1zF98/eBKqfZAjqBPX2ep
lsLLGFaOnwWlvMNSmihRZDVUEnqneizRTD479kXn763gkAhBFIKdJGlP4u/abl3TIgTorvZ0gHtd
pJzs5wIHOcmJbsCjNgrOgd9e6QGlSzv++DPZ7WxVorpLEdHi5zxAAlPAYPVlanYnCBKy3pgBvKPL
ksG8MGfIn8ZuZfOnOoVC1YJEp+8AWLcQ8xDvLz/I1auOnVQPmBzY4bTQWRrPR70YnRDHJzqaNmnc
pf5nP/xNmpFhpSuTxLcvVzNqci+iaaQ5c2ohmp6cMckZigl2ZWtDrHOLTkvWDJQBVXEp+JjYNj+l
IniBq8LtISCTRd31LbZBSMdT5ql+rWcI2/GTmmo2g12CpYiBd6/C/osMIccxtv6hHHoZgdCupg31
++quzw9zVQeXne8LOj2BAPAhjTzU2KKjzxEHz5jUfK9kuiVftXpdDErjjVfsOjFJmvNLVofGMoHc
ISV7q2iFOIWoC2d5HWk+RmmagjlXQskwbvrbdIt+376Hnnmzb6+O+LM1qkdso1h+HrUt8BRcGCni
0GbcjAOFUNWBH4R/z5m2hwiSnoR+DVIHs+pTnCz/EWO1dIozfmlQ/uvLI3n1QUNMjWMj6qPb/d6E
74JVIhLnjoIWLPAynQO1dplcKBLbbx6ZDKYmflzkUBY9Ur1YRcUzrjHr2KMBAuHTjqgaSc7c5qgm
EdJHhc12boPippkIRgA4xs17M1z2blvYqc9XZTVl1dlzU8ol+UHoKEF72LAzMdYBimZqifIw3stn
UKxQ/bpIzYWaWC5mhVeqCM6Ze87dFGUStLl8Lm7duOZ4myICe8ozB4J+VNZoI0/7/z7dmLsTa+m8
tyjX4stywKEhe8McaKoSydJuwtJLoHqMwLpK1WefC+Z527T/FT5IvynbZVs+2Nk7KvcMGLKrDqDY
FFWBG0n7Uklt9ksgpD9qG0sXUEyzclMlnCduCP6FxM4kP6JrSKuGAfZYTWIG1puWPdUYqmG2tc6t
WxF4k40nlJjc2asoyBui05HmM+1gx+6dLgOhEMw+BBzsR9/F7FZquAxmOJDAEXiuKrJElu0A1KdK
iueQU66q6B5zrQMAaJYnmAzmKNwM0MjE7oLJg6lOQk1B2Nlucno3ZiHaPBxfy6MBekQQ5wAG2L5M
dRfWkwYBMdXmvf5l03g08UYgPnIXR6F7HE47JnBCfC/vTmGD/6eUx4+V1xNVhZ/ZtKA4yS90Na7h
QrivmbZMBmmRtHNFa2u6YmmbmGf3MHXP/6zFlmwLyMW3WfVRu1HQUjVYpnVyj9dVJ/5yTubMXeGH
cMlgMDVLd3HUPDtjPE3xkKDc16qCdrNxqLdqEBLXPIcQDkXrtvWvcI3XM4IT+uFF/AHlKKst15gj
sro0NeHFWatPgfrZXsgpvnm4+bDKNlxnCj04G5CCQB0YFKt5CWRSdBQ0m6ENcFWxKl7shFee7pPT
cxWuGHc2sYVldg8IU2n17s63DMuK4T6kDF3t5zEoFhJ3QL0I7N3icATM5FSAdnQyr+wCjn7XvyFS
EMmymDfuVDNippXqH02ZF2OPuZg9Xx7IUOdmUQ7XObJ8CK2826GGMWPrK3POgZ4EyRZt3wRcNYdG
TaCEOUosD4JDYw4AyRTvwXLjkSIxl1k347plbHh52z9J/WS3MJef89HsPmAjxEJNMqXyrgrS/30y
JUPYJtIsQfc+0ELWCXqEYBezbHBSsQPSGjvlq6XHTDpYgPW+bre7prruGP6bkD0rn+5Lh7m+BKqt
ZC5acA0LiQTzNw3GaUwkHZK4ApmCXTlPp/VgpYRyzUvRGFge1rkd2B4TAbqvO1SwJNm2ssmxMclo
ji36M68N5UeLu6+s2SCW8m8+AThB2PPWpkjCYRPqsIhPuhQU0ymZvhDuoYATncKZwZRrLt6ZQPxp
5Nals5i3CQVC0GaFldVPfDKCgkpQJdcTWv/cGDdUdzRdkAaZYcHh5o/dp+su9EMk1hukSp14quKV
oMM/OTJ9uEMO0L6WORwspVBLrVdL1XUrK/QxT0EeUD8GP7c/i8PsUKUIfHwYxI/9l2bfsYtoW97L
cWyzQKH9pfGSbQj1bQ4DCdprkzoBkDNjrFS8g357QvwxPdi4EG6KBZmzz/0JV4Adhdwkmp1nyUzR
Uez8xs6L8o4WpmezRO774COnBlzprOPWi8pfBVhUnHcKVmkgmQjpH1qoInf25h8CSBEjnyMwYBeZ
Ems05UxemnwLZPejgKSDvWzFYvfm2ZNneKfoFzMaweE7ZVfRcfKIvtEw8L8c+VdwievgLUfscYu4
c47mGpyci4XZcTxgMyLbDZA7qEQUIMLCbCLrcGTclsqZJi3zdiqUThP7Q6LAbbaiWCcBy2xkv6ZB
KtgUNK6+T4XkKUqiPEnYjbXI6SFGkn0DDhqifeJGuZgGkfHwK8Fao511iCNZ25Y3Fd7I3M+B5/um
MqgJeHDrRIgK5h5rPvb6dlGKl0hy4wSlMviHy4lCDO5NExQvi8CVQsJipa/Qa4I8ZBCcPomPzRwk
KYmUHTwLVF3H6+4fVzsd99kQoArdsWnskqFZHoRKC7uodo7AsuMZgQLLwc38S2DU+bLnkHdQC25h
ay1T0/6brwfVPVnzp45s+GRX43reADvYJ6UXQlsoK4YhdmcKZtLTMuMBTE1ZYxkVGWSwevnf/6cJ
EPC7Lx4DxqMWPLVIF3OiTkNCR/A3aMHmDJF3olBgXtknKV/64+mU121fnxDbFSlWmjwwRlV55UNZ
0yIYUUPxM3r8sck2nM4ggY+JpWQPkiKVBGysnO/3g/Y5VjPGHDEx/irQxkys3uxj1OR8aENRY9R3
/4/OOzfXwI3h5NXSXVmDwNPvHXFIrmEmjlt0lZVPeJfTPxNYfwocI3IeUM9ohCb+EVk6vkY6wUz2
UFA8wyz39inAH+FirwUIuQpcrtpoXX+k5wEf1KwBsAMY5YXlOXQVNjagWsolJDbMPa1yZMdzb41q
fdqtMf1fEKw0kt8cFFEo8AaIdWZey3KjeHeR4VcfcADoYkOkaK6h/CeXFlq5xVu8Sp8r2vT9E+29
334G78anrt0qFzHpBQ5v0SWvKs5XY/t6pDu6hBov4aw9Q7etcy5Khz1dUsITaU6wftKvkVmN2b0E
DuINoa7uNX0y82de2wnjaWV1aXSQzo6c/mt/+pHrBDUS9apkav8NTRUepDoxYvgpVnt6oUc0afU6
2XLcDWKKJiSwyFs+4r0QffaNINkJu9nRaOGs+AksndRifx+80ph5Pu4daFsz3ZuHwnSsdX40DNk4
Z6S9Y9aZ4xT7vH010CrCMTehYIa6NI+Gu2QBOtyaCan1Crn95e/q5f6N6iH9NzLbsRrBXnIhCkrQ
hA4uHDEgmjSebCsEebftcrbSqIcbK0HJ6BUXzkDLiojUmlbqnMsFwapknYBTVjocuNXqNndSSCNg
+wEkpTMIfpjqQS48AOlNjPwVxs/FSYb96xlU/SqiVUTh7+DxFCTwDCDHro9fcDik+YCd/evN27be
i3GcTSuXHiKfGxma+2MiMbpW180960JDd5Ff/2uB1RWLZTwWt7CDgV3pIvK3+NVaP6s9DRZW5LtJ
5kkqpagGs9ydkacVJFJ9iJlq/kv7vfWPWLHpigrbvBygYG5WSbFyPta2EpBZM6eccOXgVuTzfvKd
Bu47Yu8r665HDXp75BkQSn/Ml/yXTeoKrU20DQAwjKT7x9EeIYHjTuayjt2CtKC70i6rnyMucy5b
445Zv9rZVM6hmxBofdB25pB1b7vfyRAn9r4hSJ9Lhv9n78jnQbNKyF0RZUDcRk3x/ODiLiTgzL4Y
A0u4taCvIQMAlpOW122gS2sRQxZ3yzxZc+urArFdKuHIbcMZR+6deMS2RjlrUSIL1vVytJyWNH0G
dQ8gS6CO78rkpOXnIuyyeqRABD8hS7sJVAyA9bkrlp+K/psQb5VKkHKC2SUcI3zTS0MbgodqlYgm
LXi4wb0jEd0KhtuxS02aJaj8OS9KacRlak8Fon6sQxhhWx9xM7q3Zb07bqgUW4PsLbZxaDcWkq35
5rYUohXH3KX9kWcA8KQJ/sSxcWZtrkPu0JxWcFHp8bzqqFDgIk/SjrNXPLNCgc0VKLC0sqxKORWm
VhcWWGWthLJ3OpHjABZL3M9UsThJoMOxxh2+OzNTAO0bjPEa6suJDLHqn0zyBlZMeQt+x+wpkITT
6U7OYOgdiJhnZ3H1oo03eN7hYllkP+lQYsabrx19OOWyg1JMig+K5gBUKuv5pFKo3VgWH1ccpPZS
p88EVLUIg7mPjMqw01xjmExl8GTr1u7SPw3mVYQ6yV6lfKzkX3pjoJHap0AHbAA2eKKAsE/JSZ67
p3dnez2K0eYKHKIEwbjYlY4AVCwlgFpAlJdmOu3GZWZIXm5x5ruJyAUCkNtdM92BFt2tfxTjLCH+
rK8nVIIJ5hoxKDrLHxAEKqwtaO0aJLqijtMNayh90y0xXLO2NDhZXlf5JUBru7xploJFtj4MdHOU
qt27JQyPLwsXXvIKaqWcFimF6hFMeZTYTJo1cdPI4FJuAemp9MhJKD7ne8Ebw+ZiSnOBjMirrvmh
wYzm/nW6zrrsM7PGp7xHk83L+aXxUlUt2+Yp7AiH79bGhmlCeQnYjWSnAncVp1jgq0tWjAj6eehs
noCOS6VKMRzWv8xMQuOvciTxkdymapAU9Ge2+VZSzhFss3FifTzBxv4EcQBGwr2IdLmWpfMb+81t
hS0UvgBC4M9Bn21vS9bUp5RhfuZe3kZYOlTemTbxSqn4gDx3K8HuezYTxMAULs+gDULqLFFQEEZX
tB2rLEsMjH+CqP0eb7I5jpx+FfUfl3VVEu9dDN5MVF8fSkd6WRPUGgPezyWHEvbxhWwNX/GaSx3e
2EM6BZAk3CsApY9FD15L9U528kb7YFo2tcnh5zhusnwhJED9q5Caw+PGR9N5vFlSs+wf0WVia4tD
mN1uVKPyJqH1fbeez9lvqidlVuhItdZPlafZCg/6ImjSIgnukrJpX2OFK+jnH+qkpIzUWhZfrVRm
xGIJEUx2dO2RuYFBePChFILttzQyUAxqePeIxNyfHpkBAatQRnzyGNzAITKWTHVy6vOZuFoV8mcl
c00SwSOf6rrPRYT3VEwfLDpArm42FT78BMVGemOlBMLeK2r3Yod+cE/XC425IK22mH9wGoMNvYkU
cVd0JLx0jrVhgciDRlYTMNji2UHWbvE5Z6mCr+WFBAVD58Gcecr8uBF81SHYKwVW8t/1XNiCKLa5
PlCKOMHUNGN4jSegwc0+fLbUGZap8IApCqnaGCmTsLfvZQ0fWENTXg2ovY4BFdyAN98AgIIWYtCk
K12VatgU3N1Pe2vK/JFYrdtzelHB9XLQd+R5n44Fjgg2+S0bumJqUykq8KK+B6acekBnUdJKDyi5
lzgD4XVvEW/tcWaZ8/ohn9NRN8w3PueaolTZBhVVGqMSVWJwvDtDE4vx5Rkx1XRJrnzFtZgEvnih
WKOtAaTXQse3uHEdmOhg92vFF9MIMBnp8jEUxHSDpD2yGkTiKOkkHhMdWGUjqN0CJiPJnZXo/AIz
cd2UtPd220G2rZfODmxTMs11QyH4LAa4wTO+BM+wBYq4nWOliCIAE6Gc+/tFn4np8yM/NIU71Hrv
ZmgVMOJlZCoLJou2D3U+fn4EUXHqTq12d5p6xJ/KJXbWlHzklQWWAOf7k87ZOokAgLXWA87jmZBi
5efYWkEWJcLlqoOt+IGC9CkzPsB17aTSiGzHGL5vGnZ8OEq0S3yZ/zi4hpDqgmOm1W13mVj+DNGP
i8WmmprLgWV8MzhVb5ENVWbfZjUCNuoqQLuYq4x7+tn1sPhm2In9rrwuq03yCeINmTw3WIwz8W4W
oNpXypkuj6y1EPPwpr7py4BXEfK8G8HH2jNJ4Uegh813slCgI1s7e/2lCVyV0oIFxWktzSrQBC/p
6rZBtNTtI3N2Y5ePbxaYPMKIjLDR91pp1mSlEMlM7P3vyBC0AcbQXCA9Z0a0OhLtk7eMMRKTH426
oO9zhs3EVoYWEqCcrSm2rdbTORQYZTtUcMyhyQK/9CEB7r+4/IHCIH5jxE9B+gyour3wpAztz98C
KKiObyM4eFJ5zz5k6vMS19Ezl8ek2500UbX6pjLEgb21dhyb7jIB9Gh9hweJnEJkb+WQeqeHD1RH
2IaKdRg6Qa6dAGK9xFU8mlXG74GWWgFl2lFj2I3iTikf1mNF0A8W7WQMs9ZXKjceresU6SscqMuU
o7Ri2nNsrbZtIaiDBYEfcKVHINChk1BfnVtp2TUU27/y333yJNC/sk4RnZQXGXcHpEGIAcgrBVV9
1wAgIgWvEmE1K8ExmcHLeg15jUgRmkyFwyGi/cEw3ub1SbyETZvx1J2pEXzQuJSmq61HIN+K0vEz
koe2LAgpori4YpmVwgDroIulqU+KJkNxDZ061ISXI+o/T0q31chBbCC71FViZVcAqBvknipJDVOk
iEiKyFRh/9FPJpeuLQ8CwFiH7HC012Sw1i3E1d7WvVzQPhHY19FFuxi0M0PoI4OIYqjyTKbltnVG
QKr89qVg2jhUJG2Fa+C0ddEJamr8JfYMvnHqV5PmNX2w2gUqG1lSE8RDLYteANnP/MLvROzFWGko
3iPslgnQMJkvR5ltaZ8CzvnrleSqzHdoPJGBIYrWnRs0pcOlZ/oMYlT5rgJvx2vGEPVLgwCIeYGD
Jqp88INpoCufJaRIN1J92PZHs0Atzd1qptKP40D1DiRx38pQuZF5eFrTQw7dRX6Fr1knGrHBjchz
vcccJO5wNQXOHTld/MKEeLZepKPW7/OTZYKKxKv06TQwH5mecqq5PCQH0lqWNbvjiLBNzbEfvZid
NLZmuJkuHXxSHsaAqeiUg+DSwIYqYXbi0dY8SUDOTR40nSJREjuSHPeJV+RwutONwa3Jt/VVhUgp
c2xUzTt/S5oVRSkSlvt9Dy6cFH4VihkTMByP0Xcz7MkBXEvxKYrIz0sMBZx8tb06rvwSQdhI0RGd
WQ+ZInhouRkSa6vIDrwaR92kaycznKEmgdaN1sWsA1sDXQntYihfnIcFUvDIm53T7SXTFC0dqYzi
QfbLr8jx0aZcBcIM1XoQr1d1picwV7ljoFRoalemrkeuktWN7mY086sWlujVMkSwMF3L+EEDnJSk
jDnG9EU8QvjuYx2bEbfycwrYoXYOmcgvIDsStmODFtvC1VcXPNwo+7P73A8eebIK5QF5WmGFpF45
mv5yXvjKkl097wSbLBLK26b0a1igP1mW2CDI6z7E7+yHE4socFTgdIChR58oy+205B7QwYDTD/E1
fxZmD9TdNyyZnOWt9kx4S9LoHygVwmn05qMsZdob4v5uFHkv2dMH02q60xciRZGOxSc/jOk9CGCk
sGx4mrcSc5uh2pTPt4Iwi/RZoP6o1x8choM5rgSoC0fYqUpSRiQFQdFrNVfMqliyftY67jd+MIgy
OxniU6U77xzbMWnqHZzxzSR/GD3GOJsgAUSl5YBHfCRVDOGDrBJ+VXwPGl2AsUbr8Z/9k1iLWrGw
6bowUd8R7jatQo39ia5T9IPLiQjXbnJVyoNe9civLv88Ih7QudcsSavnwpr/TLklr/NQZBgWJprf
nI/PVtF5yY13ETIBDzya73U5+dq00z/dWG0QKnPcq6EVqr2H8/Q0Mt/6z8hy/jA31raSKFBdAJnX
TVl0lRC8u5NeE2kgJXG7EoxZaevenca/jnKHs6e3NYfwsb5xV5aEVXX60tR3W0dDX4GQnGCAndit
OAM6yYjgoPT8S2SuZfrcqVPPWPx2yBVECYuJZJepCsbqA5oBFs8BKMK9B49EjbeAnkK2S3G9ZX4Q
i5uAYrBJJByq3ZZ3W4CFyAxr+FiAOfld+M5aZxNAloOBY7qzLw3CGCrB1Jg3uOCEKPSdaionqEYz
l1loqZCuvZOk+krY/M+awzRleUyRUfA0N1TnzgsF1dnajiPPd8uGyz4COBX7GX6KDtiLq+grlJZV
s8GMb83csk3FepHQuv/GiLEze1Xf2P0uwwCbljUju4C0IPUw+ulUeWxDP5srDmx4ZKv1PoVzmvyO
h5pbraYxCJDy3CR8ZGQN7UNERQJn8jUE33Sd+W2B8B2DUPifFQSNeCrh0bnVItDRAPa6uuWtXrFE
Bv4BhM2cQaT/3NtpKxE1l1WN1mPVhXCrNMn2t83HKo/ZJ9UrxskoLGDFjZAujQZ957WCrV5jpV3r
54bPImHFdFEbQeiqG9gzbl2BKxPZkC4c+KiPTsjjZwxpGnob73hcEsV/JMmeXXVq6rA5G2GrRrPf
SmUXF/F85bo65CpZowqCIoF+ayrkAWz/M4hhpaTBRFK6+vOQFils6oLpEnBukAQsrizcx/Q4ZX2H
thk2VozwcS1/IY1A4iluNC/Y9hVjJPwDaHOlL4EDP4LfKUJWe5JbWApH8mKTgNz7lwFoYV7Ce7hQ
z12QswkmHG9imdd7+oSN98Of/C9LuSEDkYEp76eYzv12m2PFSafYGmjFafawzpQRtv60da1tpWsn
z+O3HvFrveSnfGsPDrThoLFm2kaxLlu85Lbcfqoy27IIaRbm/xzO9RnUakN8yNoEmpS2/Ug19SK4
xlW+SaTzGkNUUIXawXzFqJ9kqQ58YVetQnhapoY+Ermr7q2znL0cGtoFjGgGKMvvENe/R3bxo0F0
gYtkJ9LJyjLfS0peP9WPALEyrZzisDK9YxCLdeZZghQ/SYBMgkrLD8EHQxiz1vB9fAIcIf4wjC7X
+o07XIu/uI2Zaaz/6o4f0+7sb2soaRy1z0VowlOZtgs6GVAIjecYyiwONoJX8vCuo6T9J7lH6nYQ
BedEO8W26IRArk3N6QntiYFkW/cxK+Szv2mESAlsQKI6cgsXQap90tJLY086mPBS7VL49yH7qlpy
G/3iwJoDVtoswoCc8qfKB0XmtFf86ByFI58bj1S4+jNK8a1u1raEtBmp/QuApOmPtXnGwBYy3mtk
xd6WQ+8OceJABvVBWza3M7/TSSmk9fzed0dwgoKAVv572vhjWB8LBO0Za/7NSVTPqJGkgMD8jgJL
coaV89bjiPa9modsOn5BZLvXNyvJMgzvCoztKdWUEFQoxEqxcmmf/BSBiAvC4Odm3zFj/NSvezuX
JSk3eZ4it3+CKUCgykgcN4ZnSeeGhzOuuEYcogqOVlGOXHI7WJ5qsxGW0+P3KeOezDp/X2w2lqID
HM4mh/47Yr9hH+bBcqrLh/9WXlMmzeqIEM9JekImtAIHMF+M2W+p1CPN1LJwyU1+eDUlgV9x4iv3
F5DCnP0Sfmeo1D+U2BA8C2N7R4pWHl0nSBVd7T5KLyvjR0RkyrwpRvSYXnveNlbaqASHuH7QSPfU
udSQADIH0cyWQ5+3J8Efiz04dqBV/cUKVTMrFKOxMP6ZHaMMzML7opIAT7h0WoonR/PXxSpmAt4W
ERCFc++4CroeElNW1zSoHjjmKfYqKPabI7/0+QU/jQ45ztsVxEKAjYoQUhZjG3FKdR+hyiHXT0Wg
P9Ib5IYUSSHPZH7X36OzjaEbmRobA9oj0M7+7YEt/+p/KbOFJdbAhM10D2PC2iLahJ+PWWQufYHu
dJYPav28bWnlzDY+1CqGNmDgW22NmLQtAi0bpxt9j1jlb5LDNs4df3/O6QnFbtkqY5i5+3r3sfmi
1+Mhk+gdJ5ZiTan8bWc1lzMW6Ets1r/4SW/eaNYsNI81WhPAW2JGeO/qFd8Cjwtjn03sAagbG2XL
+zd1eSxx56LxwtZ0oIeeOi2XcCpS8gkQnsbXG6r/+Uqm2f3HVDouYqbBzOr7ZJDSczPpGfIoJjiT
h/ovEUVDNAwYon9zBc9zkqy0OyQfTTEDGvn8VfAEg3m5c/i44MdK9m51NvJ1zFFUzJbQXumocxvp
7mVq4VelsBIDDlXuofZ0HV0wvCXgErE8gK/ioVdsYPwp9GzSBcWWlyou8/Vv09em/XWam8o1hvD8
DniQS0wHHazZlIEmOhQtY2ZxgKdQOpCTGb7yzD0raRcKQLYrn7PVV8FAlGCZhMOcKb968yYNsrZz
AO5N2ng4rgrQ6gCU+qWT0H+STaNrEm4bD0QctrkbnTDdUKbmxXKfNGKPR3I/+ewiCfIkhFYn8RMA
ICtePgIzQsDzwtJv2S97a00WLbnZZf7IQloJZuDeWZibMZK09s4+hmezKVGkkpTyGaG7r6WZnjBl
lPtWLUGFGhXuiZ8S8hBdI1HRKWqwYSsTnK3s2oW0uFIzUz+lK62VO6vLygjLIwSu2/wW8kH9X9mg
XMrmy6yakKnvoU5+hMmKExrnVcFhiF9pNTxRqlHwfSoDLxiZnUeq4Agq64j9qVlEA3+R77aiQwqE
3CQmqGkqMGybJ5A3KhnvNt4O5zJH0KGistbl1N1VrR2HLNPJineoMwmw49hlFiTupDWnL06CvDMv
5L0XK9Ln4mC4D6oXxV4x3qXnL2t1Q8AGTM2bCzQmiN7mUDApCX+k81bdEQklcyPs1nM2hOgeb02+
6l+mbYREqYa/GN3q1npFevWLj9iGxEFuwAm6i+BQ93VHRDJdFfnt/Dw0Y3Bu+KYQMZGIPwuy9Wu5
zRApNooVJVKCKEoIuFudGMyaohvUQYyq+TYPgd5YsLhdBf7vmjsyzo79FDQKG6KwrCDQU8Zxg/ot
lopQ7s+y3OmAZElzbjeP3Nylqmtj+kq3lzY8kepgij97ou8csvAsRlYlyAFKZG5nHVfeqgky6flb
PBZyME3NkhlcNsJfOaKFu91j8g+oXVS0lQVyPlYeOORaddepb/p/SpxQo+Y1WoqdwS0eOnEjOKtt
ZXmSNiQvXkhx2P3yZMMw5rrT/zBBPzL0vc4oqyTdmUBPO9+A+vQ7ZEMENH43i0+JEm+UqAz2h1b9
sjLT0n/XazMuhOBO6RTjdXpYFU3NOv9jGWy0l09hxnalpE+0CORDv5wOc4zgKn8WepNhwoNBlHBD
k/iSbDKB55RlR2ZuA+zQFMVKtaJXfQNdg6hYtTygMWmATtWn2CByDvfZuaHAx9TD5Sa6UmypBHGD
VPAruFs6RTfqKdgrsHLzhfte5BznkL6WAqj/E+ILzyP0bulK/i7mf1+COnnII3e/SqPzS+BZrgKV
Z5dbnrknKY/D+0XTkCgbtjJbG9m1dPcIyWQMHNZMJPMc75vNGxbbrL5vsSGN5olc6ERgSwnNdNu9
L4VT9MYD4QAmpjM5zBgqLLvczq2lMFcFbuBbqobsBE2ssB/q1Ava+nIQddGUxSbG4ikLdpwjvPq9
ArqfIOO4ioZ2HvkRfUQ9GBRpsnDpHTuyUQ+Oa+et9b5JtdluXFi7vCRHqb0eDkUitO1Umo7AgBbV
U9K32IkX6qDlhdmFiVjJ/41zT39HdwfFPeDEmQlyxGkFbe9Q9Qz36l0L5gWqqQSxVRc9wSCGbcOA
V1aKD87l7DArhufYgmzfziDEQOvzQE2Qr61Z5R/+q0AHv64xcGr/ap6HSjp6hi5VzAwqGicrFAsX
2cBHkQTL+aVsQb9fMF9A/9GMMjZQMSmJQlZwDwdn3YRALWNYCQrHshNZiFM8NMkOlC5iuFZ47vh8
ZTvwxbb+vKYrZeSdpIBJjEL0s8aGCexTb5cZ86Cug++VS2mS6ob+wLd0h8H6ljOxh5xW4Bb/y4Av
3iMIZT0JmBLfqZHuQS3LpMO9veY+kdb7Mu+yhOi1wYDM5rrKwlAH4BbSQSEmlQdcw27UAKCVtch2
khlnggk2bst4KCYCr8zi1LU4EtO+q2DNDNGK+kylW/MujojeCjMRk2hrO2SyiUSucb2RsEY9xgEL
Itqd0zgxjcwkrbzKZf8uwvG7W5+7Ff8ElpEdOZweooALTlnr1CJTT9PHLH/HUa0HUslisdDZV3ie
fko8WbtZLdY+SLgzMcg6xREWzE7IoHOwj/fO6cZ3mkRTkQkxm5d+xbe+h1QVDVA/45JAYJ6KWkY0
RdMSPPEAoH1YlTKbbBvxlig1fc9AnF4VbIALJm196sJzCtEInmrxkhqg57mz5fSt2jUZq8XjHIDA
dXZ54IMcpRencPVpB2NzUEu3o4wR8edTI48NQBlDx0SiL8ijzkeqH7TnklgLe766J0t0mXLO+L0r
nA9lUM1IKCKYPpWqITA9YnTqJHI8XdSltZXF5bBUIgeCn3m1g2xxJhf/ymrAzLwQT4g27XVeJmlB
VxptE1Nqib1cKmBHhq1lrDojx7y6y2NGqfTPiXA3C+djNhW0dBJ9alWR/ianQFevZHRoHzykkVZO
LIyBLZxfk9jgElK64szaUxoOHDydTUifl2pzQK3fmr9HZqnKGmQ+urYYcnfOI+JtnvnxfjClqxZA
JQUF2fE4MSyeXkoS/oKLOUu3jMros1LZGLdsjQAtiem6vVJJ3sO1/8MdwXCsQGf0lTrZjuM5eIQs
Z3snp38Ivn6C8lwIxrAlrlfdTJribmi297yXyNyTtHSuuDXE/r9hUed7In0QAtyxQCKPs+8e+kpl
GzUVB296fGb1rOVQJTNeSKDfF1zcvZarOoK0tJhlWv2AkHg//7YbfBp7ApZSUAw1rVY5GxhjcLVh
tg7RPvF3X7lufS1tgZMzgPlqp+c9OOhEptC6B6+d688XfvSPskSHWND0fXrK/En6NvPu72S0YgZR
TGrKX5+Jzh0ZpS0XTJd6w00esW+tFrWBoBrCzLbKNi9hyR1xsVMsVbNxv2Fmnakq/uQ640oHgGUX
E4aJ/Q4VjjjrFyS3MiYmCNG3cNFaXz+VN3upBnhxmdKo0ZRCRhHyCgzPMFRyasKHdZVXmFz+hXnQ
PD9oRj1PbiAc2ShC7GD2rxYbUVKyKeR1/Z1MEuGZWwncEVwsuOa8YCL7cBTvuGehXH07PbiA5hzr
Vp/MMvA7n6A0CetBJt09c+itIhmB2fWkOzTMxrqd+nMwf42p1Tv7nLRhWR5n7Vbf9WFXJdTMaKsO
DxeGS9vnznTi2yPjxBkCVTFBAMmRvUve6Y4Wf3Rbg5VEgMqUlObPUDsPdLEY8h9JaDieHksUP4iM
+3DU8iaKzOa7QLDlyf4NnFnWMr9cIaDHJu7q0KsKZmLL7yRBIJrFxUFpN78vfR40Gio2dlry1ZPK
chfGLi3BGSl1aV5AtyfyGk7fymSmCdLQ1mQUSOCO3m6ydBN3zhTdF92vziZiABfhM/uO9NW8+Luv
avWS62g3gGAsXnTOGtm+JliIqN/RIsXB6HARjwQqwBg+NELP1tF6G1fcIGgjQCKNeKfj5s5v+Uy6
FVgfUFSCvtNdAnxpj3YhiDHY3APG95nwHi7Ar3vyZ4phDrRkaXe9618LYR4j6QPiGkeZaQ96C0Lo
3lkMVJIXgjq9lSV/mq/zjR43ng9Ch0Ps8GpsOK8D12qoAvY+y0eurbo6PlHM4H7W7HR82EvLHRbk
F8jcmITRW95T9J9ECr4zWbvz0P4k2svhsboY4mS+gvqEyk8g4TV+NKXeY0UtzLOgMsqcW7iFOxQ8
VMlNSzmp19YtPAIwUhXwuaQ+/3ekXO1fGHJg6LUJLy8MjT3OzER09u4jRWKg7v4RhFROebj5w9dW
5ReS8R6u2RdptORzW+x1BZMpMcxsPk2E8+4Z7ogVlCrhEizugRZmQQXhTQyJdMr7G9XjPTjMdEX/
zcj5q3pWSEba9fOojZ/kGaXazMaySYBv8gmG4SFSARULsP1s1UTTSOJpzVf4WC6YioUZN2kCQDhC
h2RyjV6v2urTPFQHVN2x2LnDiu9iZrvQsj2+AlCtIbifgnpp+r9V4NFXJmMwJ22lN/+59jZ81DE6
McX2CxaKjB+v6OjZLF91sEGrVY2MmvzDtgXI22putULhqxyuGazC8b4CTGL/pAxfdWN8AK+qWePT
zaLy2p0pzwnBNTWT0QmDA9PR1qnU1cogeWRgHgB/wc4ct0gWjaJ2flqa+JrMYoxOnTWlUts4iw8K
f0NOsZFj4D1vq+KrxhL7V2huYD2y2a55hQKJxlnhNU+VcNnY2QMIM0kzST20bQA//KAnUjC1M6Ca
QeL4Iar5EcOk4uB+fg0R6u9NaNXYJ++9OY2vaxF3NJXpBnoZ7sDlxK90qkT03seKRyXtQoV5iCWD
zcn3db/oxuALKqyzteoRMdMBpUV8yIFSThsIP/8bWfUzHz9/NAxPD2QmpkMXQtLHTzEJe3Zs530q
A2HkaruB6WFI1v7FwduqJQb61Q0eLMnsQ31dHCv+gpi4BlT6Y6i2RNCrMGbOHNRn58Zj8oUw4lar
ornWKGq3f9BFrAko+PfiZUpp01C6IwZtZBjNT8TdYIArrJQgMkSl4kDwwTalF++DJf2ZYuoiYZvM
6QPp8QJYGSkowpDm+qPWPakLxXzt0q90hNRda+5Pb8WxppTfF2RLrSv9fYqmjOypbGFD6sRVWFeZ
I0K+V2EtSYbGgKxzDfHES88HQ8kvl0Z6cMviy/Xs/698y1AxVtp5kk8paMWQ46I8PrYs6x5cGyqk
PyofTcfCS30WSokMjG9eP+6M6IDjRIbWQklyG088t4C/GhHvzwwh17BKmFMyjw5x8WADRVM66LJm
kk/4rkz/8op9aao4BOEk+NBulcC/UcusvF9u6QrrBDifc8UkVpwBkDEYPIqHnGbM/n1Er6TtC6x3
6aIVTPIZDgmMlay9yfMSp8mfNK3KZcjPmD0BTSvkoYWOUk2UXQFcqo7c0J7KM3jqW1G8MKIKpcNi
r6pqfjM1XZYEyMQhgOHlaoiP/cXMd/ZG8g/FayiXcwiu0Go8I2Pq2iZ+NTbIDMeyNFo9o9wQevxJ
Sk8iH86UAJQryQfyI7zMnGMN+8XxqCkghfnT585d3HDLPMLjarTxbhpWgeppJj7tnujKCzQbLt+K
UG5j4EPI7UFBxXpT/XMtFCBJe3Z81e1jRArBuxKD4V9BnPhYdiQ/m6TmvjuOXa+pYMeUW/7CKLPm
bI7vV/B6y4jHMzKhyaIDSzoRdOYaWZSRAmHBvua4p+rr4Ma1I8WGF9IbFc3gYhd+TK5dlmYO4zzo
ID+h0RgR9rJce9RsWtftJOoyc6P1v5Ojspam/ZpLJ7cENt9N3OHJ6DUbLHJf8/Cv22SRTgYyPHDA
z2vU3cVRu0UAAco09keKfOWxdPnyCRBo2eYaA614c1Q4kPDhV2K3vPWp1qke8Z9tNWulxGu5pBBp
KMJyVJ4GGwU2TvWBTqdmwwbNSDNjW9esJFJYjHhXXCiYG79YuX95apOLgo14MQhIaIj3ZbydU1em
mwGy96fHLuwGFckr04jZVeviByctzeEhfh8zP/+hayNWuyILCjYwetqCn3W21XXWL84b5A40QXD2
AYcd2ZmPBIRqLpbq0nYPMHXG4DjtT92WoklhZmKjsx8iiQzfc0LZL3NiIKKrBAgtFw3/idyj/QH7
y9L8NpAVkmWE5RL+vZWHTNzsaNp6Mwuj2UsGZQ3Aa5s8xAtmiY/Xhm3JwKd4eHF/ASOdKMhYONSx
IGGhW7hCa0LhnuhSqQATG0cWi0VkbhQpKqaz6zLlHCCHWNxeQcdGDDV7w5GQqcqIFOWJ7SG6V21E
rckK+66ZfzgvF8RKdUfVENuSLjZVhD0Oqr5Py8VlS9BvdkwcOefM5lQMLpGPBjTGw+pNUUT5lObU
CRntYlJT0kVPN3ygU1WqLicVbOlq0iXj3HP/TCuLlCFfnqc8NeXMw7fbfhCZ63rTyLwpTvCYIAgM
CSVx2r/cbotEEUA2byDgrzjDyO+owB+hd2TV1oP24AWHMfeoQPJbaMsTzv4gDnO/IGunQV5y+991
3UFFmYyl6aIXm6mkvEoUVmyKAnDuem6Iq5gYawKJ1IS6GE+g+0Fg4vR/+3FyKLBxfNe8eUwKwa2A
UoNw8SB02s9WauN3GKGkWJjLQtDfkrrk7kowp1CIZYoYMMf/+5sf26LjmjYhDt8gHDo56aU1ZvJs
IyrpuNTAUddXd100sptWrNNgAulwUFm29LfAgrZERUgSjiaahHqfkDsntQfXDKf7QS4Ufr+bgrQk
OVG67zQ0K8s1r4YkSR94NqwGrHINLfR/PWN3lquaHlJ/ncz1hSc697tHlYZ7bTHiXEpFVG3+KdVY
pHo1aZD4tRL5zEiboFzCrQbeQe+C1nDzqUf1W6Y2CZVjQKNxpSfHSIDZmnzo7wgqFyJnSJdDX8ob
VvPOFRIfTmrS4capyCWcVZHMTzirCsaK4nXEmpx4P3pHBXRgTVigH/4HXm5pCNzZp+MEyRKaV/Qc
6pSkr4XInBMvXH0Z8o/9vXTlZrfV1W2UTvqJc+Y7ITUf9tngU9gVE1oIKltDEcTc8XS4UJhEcnLa
qr8fdJ75bxfbzFjMekuL40Qa5fLLyGaSWIE9bRT2cR8bofWjidAo8D4VJbxDZHthQD+wztoHPpvP
a/oqC9N21l8LO3rm4J/1DgKGisouqT2uyWdj41LqtrVe90dCihiood3bBJTLCMjRBcxfxnErk0ND
7BAp36bWlMW6ciOAyZG7t8j8KGkOJ0Si8oyg0gFNqUvFelbIFTts5fhRxr0sn7gF0hspeKZl3alO
7/VmijedDl1cq2G7pif5axV0bPVzeWCm9b3y0ibchVEIdUESvxV1Vu2ngsyTT2KASk3Kc0aDUguc
e2/K03skv9rfmDFRaYuwIHv45euflWfaQhE7eHJC7AL+UF8KUlJRaPQ0HhaOunRNwQrZNUmirWvF
5LRWhtV2ZSo1AObGFame3habmmVnAZ1/hNCgftf1H1IdTwzkwtVBs1ZunkVGYctzaDiqPiS507kj
i8CCoZv49yl109/3GXtL4roltmWmL/NJB4SAAqy2BPxb2rtLofPwI3sOS2Sx5iEPzdgFGJbJK8Di
ErNThv8ber87dm18WSNup0874TqJbdcdJp1MjTacqniFEcctwYB2SUNN+1VQvysxsM4R/uwMwhFi
TbA9GW6j2uxSXmNYI6KfC/nqchDlGFvgUwmva517MFtzF6k6wgc+/FWiRX5VVIFIR0+gb5W+30Fl
LirmxFw2ZwvcGUZt13Iemk7Zt3uMrrQDI46KjAHJatLKC3krp9yneSqqk0wCRXlTNx51kDwJPmT+
krt/244KKF73bc0IA3Cw7omUIrOrbFAW6PF6g2fh5x64pSdmot2PG9m2KutgWxb1mbileUFumWE5
gDZSelQI0xMZmUDMBYPlDxaApN7RcpeMFVHD7lPDETHYmhNKxPFxObvpDsHmDwL68AeLEk42naEH
pOozZMQ13hVndKlhgRb15m3mWqgjMXF0nZMap13b2sTqZmwPgnhijeWObdTgC65BUAaFZDu6mQ50
rg6s/OGe0lqwg4SE1WDKY1MNQAKYML6hg3EHPdaVdPraScESQpjsNqz8HU6JabBDLX6TihJKV/YZ
eps1efWhWcofYAMHGKq62hVoxpOiY/iHgVMSj4sSXJSq7uy2++V52/dH8tZnyWXH0/cuHj/F78/f
du1vLuAHAuWB85HSIi9saUvLMQcKco8gig908B4d0oZ2yfPz6rhPdiyChhCo49Qk4p9g8XX/bTpM
PGnGFdviVYVL/XejOVaBqScPcPHxpmq+K/LHyVwIJZlgm9pHCVtV7sPE4ytsYZqUfz22s9FjEsyn
7K8fdHTJM9ZojOJ1AKm+OKWLwcxBQ8Ll8PwjbJw5f8L56/bB+lbfl0u00mir7fYGF/jX2rH3q5Vr
BWnfnhSZAe0Mo3FE3yLPDEvR6fS9PQCc3O9DJRu31FAtyJgiX60Fx6SCVv/aqwoBOBvpTr5Om61s
12WiLYYzs8zbFITtYiqrkfW3Ptr6OOYZ0cg1dg/80UBFZs8R17XnYh1sDC89r6eH41usb3BAqzB1
EaYy0P1z57ZZ1eD8Q/SqR5eZGTaJmNpIkassYz6pcxOYSsfUeunhS9XdLBveg0b4WQ3esPFgftpr
jumB/i1G2HIfJfxrMGnmmrNf5a3nNGD0JguJMPA8IhaWF+Q59BSRbznRsQnASluXr/Qm0GcSPPlE
oLJQJH3jy1Os0TpOsYhUEnlRLu0w7vHy87L0WrybbdNgv9HRCykQDShfb/tJg7gHjY37ItsKDKTg
glsbuao458Ea0qxk7TaJ983A+D93GsKWzxO9eXxdMKd/CWiHeDqHjjAacxk+cB5wxNHkHvacdI9H
BkbAqel8n0ABFf3OGFbLYNZsE4ZXp0ZVm8eLJCCOs7TIs+57E7vE0+ThBnRUZT1u1N61/OZcZinw
aBh9/22i/HLrtFYW6usDUlUeQLfAtrkQrsbZRy8tgqqvg/h91LvtmGFj9kPG38/6Q5jfpgnqoD3H
VvS5CEJNG55a3QBa1KuJ015HqwCxOy0SrypecxC3VnGvfbHZlzdGgdwqU2R5ofBMbrpnY4bsLy62
cJB0bqD8IsguEOoVnj+BE0tk2RPHZ06KGvAmPWLhGm/1hqMIkhd3RRpKUP2X5vqYHnB+abO/vati
JJh2/cUq++aibN3VOdMiAoK9iDY5pQNY7X0R9aNdJG/ivKESMugunj8qgSWCAdypYYYXwzuLBxLj
cSn34+PIZmX2fkSY0KUX3kchRTCJQEbq9tjciWp1fHuezi6jVtOkMZS+aFmptfjuEFXD1jOEF2jz
IUouaYJMO4S/s75iZIWT5asd0DPlFpDU8tVxi13asRQbiaLoNdT4NoQ9Zrv2MgJ6Nv9z9xHvKwhw
DiaI4Xti5qpJTagvYEGqZ+4Qk5sArfJmR3NBeDW4oedtFK11Hfl+5LcEinr31srnuQCT1lXysUBT
oZmCyHShWde2PARgXXtfZzFKdKqIGAUpSpCua4b/pkQaPkd9UfnITyWRRdmY2FAy5dEVgD131yec
jiDTT2SxwPrfj+ysG/lzHOY2fVGovg53dHTClYBg8jE2TnmYOiQMQ2WjbxvBg1hHm8SPuRdmAlOj
8ZJosgxFCHb6y2B/4fKX2iRU3A6mPBBMjrKsn00gqKYUzyCmDhHaqoRVbEDshDuDjNTiHlS+Hofl
4ppnmRdj29Lazwfzn9darHrM5Ci204aEeRg8+/6YXnJeb5OjdBKbMq1JPCPVBv9zV9oM3yRrlo3U
BgUf7vdmZ45mGYmOW1qOiYmJtaBpuuk3tCUfPGRDwojstWxoQWrUBslYdY6gYk9XTwOkg/RBQqHQ
U0HdHd7N+2iw9/vXPiTjlOktjgNp5FIKqw3otp4vKINhxI093/1IcpE11r0aM+uFeyPwzJyUz4e9
Ar2+yW7blh2iLcbz1mD/ryUCS2GXtFmg1Hpyre+ylKVmeChadCNwsLct5KZkKnkk8CSL0E9d1E5n
pmaeK/sMlC1BCtZhWBXtYXEeatpSFbMbH0nwbp5c2Ey90ZI29yja7EzQBbacHi2MyIRduBrg5/ZQ
G8UKQqMEnARkX1MIaSrlj+TBhQn5HKcAcq+ncEUz/dlBc1aSA/SuH7LZramLV510EtS6siDT0rmI
G3VGPJYx327NRsJN7hj52vIESF6sN6y1p7rKA8mMJPZsaP9UY6D3zCCcyVkI7w9c6LiQoctxBdgU
eri/du6Hsh521GnlEtZMdiJ/up0tY4VlnNbW2iHcyuttoWOzHUx9tlmiGK3t2ahtDCQ1KLk//ynS
3Db/+2nKjOze3ED8oVLhxDWJcrTAMzUaWLbFOD6149UIVIUlzx1cASnrU099CJsCY+tjikETrVtX
T4KL7OFh3HrQVOLMjGh6CIYWzcyFIOGY+wadYFLPIsJMk+i4/Pqq1hbP05a7LrDMmpsrjRqkTr4p
RCP63ifbYR1KncurQwkOKwNtxcDEsZNXmrWxKiB3XyzPVsPMl0fRqIOlfOXEuqoSxVs5kpKraZ0J
xz0NROhqgTG/dg/g+sQj+7dYxaSZeZ6Wm/TumAOwbdBQzDtKoVSBJut9Zsf/OVPObLx8RmgMTrqi
5jN+xP2mXAJhH+E/mrZjK4gtgRd52V3QQDv58+ZPRnPQqExPutcPnOPTCgOWF+O/0qy8gksFG3TY
r3VB76yaapl6qaEygEmYCdJZeVv2a+HMvLmpLB8MbuDTrlvx0YUHY8zPlAjPbRK0WCBoMCA1rg4d
mpSGkSinvKh3EIWmh3UZZ6gxJrP2sHc14RBgNQHD+Ps35Aiphc+xKAqcwyK7fu5M/BmhTRYrj1zk
x74WBnavQTT/QBIenNhU/Utw5Fij5gI7O9H5IbApQGhwgGIBRVwkP4DFbuxG+4887+3fWTABaL4T
WEHBFIDS4TAEewEByAjJqMa7i48EYYgcUsmNbXNAjvGebHwMS4MvcRmdHDkkD32D9IbxKNxxT0Wz
PkromC5wxJV2g9KE4QV0ncYbdkWvHBuMSGrTikc+u9nvCM3HecXsZtL5d/rskarBtJNBwSKWpc3l
s5mbIa5KZjZ40jpiLTTICjTnzYUrSNQZnh9GZEt53LqROOyCFwVLvWJ0BgcTMtq3ByNoVQ9t2mCB
6iStHNqXb3hucqQYAQiEDir+6aVa5lOmSdebBr9iGq4PuIVYhOQlmH06aGedfoj9xOuY0qdAQWfe
sGZKfRHuIx9sa1ELoLG47wJzPNMh+I5Hyt6+VAGYA8UW3RrNRVOm2Mg1Ydykov87VvbqpsjAHICr
jtzPaGw8o2qdL9/RLeBCDJVquIBXfwLQOHcyO1Zkq3PCYLxdXp0F8rpQmrA7lcUIXF+eAGBibyQX
N0fhIKJoHv0clNXleezvsuoAXU2q+mak/+37UcP8ApymvbJtCQchiBGKScehj80gLKJBUZ5zYj/g
MDMyL7PC9blT1oVyxOOaYRjZvBlLgUULTzRRjw90xXIbONWL7IpAh4PMekXQ3DfS/fWvXdtxlrtL
1AyxvdYiaRnaTQBIlhsLzktFpdiShfdvCAm03saKr4l4EOnihwDL3r14POC0AMezvHjNPWrEsn49
eZxlb7tilR68qI5MgBIYFD/f5u+yJZJVE6ZwbSu0xF511ZsZfK3Z+VuSWCzGA93q2gLokLbTlnUN
WWUKjDz25qEXF5LQdDDjOdxJrPgGB92yM12YwEKq1UYj1eUvbyqvqO+z2nXkiUguV1DebvIlz7qy
zrnuICWUcbM1frRH1TkxyX7LDl8l1JIq954l2J94lsKVfSfZrlalrtCtGX3FQKfdYctoy04kmKHb
NR16qmZ+ow09nn28CKSASfysUd92PXCbnyTUWCJn7fKcusiV6QYZmO0fsnwXOxGfbILDtG7nYqoD
yqQLqZLA59f1UZuGaYi3cy2Z0nXTUezd1G4rtPWMBdO6Q/vNrAi5ksQfEPLV2VIkPB2rgI0utRyK
gWvdbIpPp5V0Kkjm+vesb787FG1yNpdva/GXfHQT0km+jg2sOrLwB2CHghK9+1WTLSPypmmm50BL
4rDIGSjyqiB+Zy8wuLFVVfbkjhJavtMMCo/+D3ipHWqJ80akGEAFajaw9YAmL0y22jY8WF4b04Ik
tUebXEi4gkaORqarQLYkOVFtWal98PcFKDOdlI4cYSWHjALhuzb1PgGPlALE58tDJfHAvY42RNQT
tarMsdFYz1V6s14jTv76vEBKRxtWU+l33hnqhLoJ85NVFNOrk1DV0A+wFntr1mBGWeTZvgkxi8bY
IEr7I459/XW99uG16dxmEhRcBPoz0AtE7Oh5uEPydSIV9amgbxGFK1hmSIlMQW13i/H3E7J4mKQn
CwDxq1OcZgos8E574P0hvNrEvD88vA5kvpvfHLYj1Dy44wbh7Jr5o69OiSIB/4c5AKMKsfsZlsXJ
/F5wcFKHU2RD6MxuJilDnCnRY14c+NpAjnc2VC2JPlQNi5FounBc4Vt4WX67bcg0Z4hayNB0X/oJ
e+MQVDlbE5bkjDs9CJeOgxOjUlFrJRPex3qzTKLFUG0vBMRRiRpYayH470Hd9iDpV68W6Ji45i0o
LmUkL68Ok79zvCXgTWS4ngc/kcoxtUD1HJb5sV5Uq8XmSj4+iwVIulSP9AKMIGvdKt6PJEjeUYB0
GV+yr6bLlbdB9oaxso0w8qDdvKZx0TqtugApOYHebPcd+wOn85mK783ZMu3wP69xxX5xuOc6CU2w
qzlQAaRTannLQvWX0HAR5Fe4yNTdRJmDKbQn5XQhrjYGbtAQ2CnUn8+283YYBVBpxJ61tRUprULG
5YWDw0dMOLsUve1z5StrG2lXL+caS+oFP8TyY5XxYCRNSLcXo221qyn9++JZegbk0Zqz9VRXPegC
tCo5LCAI1yjSMEChZ1ilLUlNJexuZcu8p5Y4BEtHTLl3PlWEvtwFEcKeal52iG7Rxlfa5+HtPEYV
dRKrCiPc+qjXlgHPye+ITYRWLzUHTzpooy349ikQMYtIH7vEYiEnwlS+uZofntQQn7Jns2xXziah
3ska0SQ8VVvR8nsSkNR9iUH4VxSspGw/XVdzjAuqSz0HT1n/v5AlOV8K8W061k8CkbOI+nD7hW7H
MqISSAGhvuCPjY4vXjhvARCXf46YT1ZghmWMkz/nOk5Mnmk6xj7t8cS02Do8K+6sX9ryejyVuXSi
hhf3nQ2g57X4mHsjz4gnntesk5NO5igKqo4iw6YEw5ub+Y671yL+28zadrrNXJtLNV06FAg6pYy1
iummrtXm9apUHCbYiXI6A6VwdNSzHiM1tQlE0hdxlOz6Deglre7lTZYuQ9uwTqAZrWvv+Mh6Gvo6
RAksW3b95TKplEmcsUex5poQBvsMuauhAXT+Oj1sOfEKrY+/Kg0Qf5zj0hpgwH3OBQkKJJj8JgHD
NBEi8JBxdC4O5V1HBKEeGiFKcI4TpFHM6Z+vPTc1jTxBTRVMQm1rW6tzc3N6vXA+GVXbVN2EAvHF
PTtoW2OS40YE6VGwcPeTMft6kMzV/1OpuPfaoLZfY/LWw70ky5mdCKAjHjMpQu/yT3setHMphTyo
rcG573MLKI2qWjh/szjiKSQXqx6qaoRUmBBOSDGcUD6xUXjBtGZ5MFBqRPNC7KkDgYJea0yZIWbD
XNU1uTnWenTZiYlkC9NI4/iLeL0WDENihG87JzBa/SqE7n7J96Nq0iAL3Gx5gjpBsi/t7outphW3
cShIZzQndhSDFNsBUKJl+LUNHK5xu9NNKRGxKJnkNgH1UbWx4A6O2fa/w5xIIX6kHorp3KcouPoH
s6Mr2Dy9nZqLsvDYFAceTz2vGScDWDsrOtFRft0/Ev+m94uhQ06Ir4gsgldn22lWgLo6NbeJEa0B
j2GVir5M5KwT9Vfwrht66Jo+JosBFLd4U7IfeQiPD3lxzEFCM6s2j5dgN4KEGyLtMyA0fdWevkz9
iulkEac+7w4753qt69NxbIxnKmcYvu7ZDd5QWGcJrmH3noO67/XW4ukOIsdgUAi1zk950AjuRRlk
z4D+UxGOTGh+slg7UtlwqFi/P4O3IxxyBHu7+UsYRFtkFD12huoNsOzI9R168eNxMtfztd1Xd1DL
n7xthlEDaLsF5sbvE/unVNDIqBkDavUiTADy8cXy6PlulrXEk5d7XsGmUNcbjHHFmOZADrqYMHSv
/uQ+DxvdZg9/6Lid+Mx5Q/r5ibfCx0j9w1VY/6dd5I+F8s2t2DarPnuYvn6Zr+pcogR9B0K9DL3I
Qd0n46Si/x0KreN3Y7UO9N5Z0/mZ4j3Asrh0PSAFJqOrTbrvHJ/+2KNAQ49wWeHsNkL1J1s/WVkM
GcHDAjZIDxQsnGfHWPLK0h2wSWO4EHLw8nySP+rPNeDj9SX9u+ekYQD6Dks1lGOyOgEXJEFczn7v
3tXjQkyy2tHPy3gdjs5fUfeJycBUsx79XTo+86rbMq4nbOgd8gHVgL7/TRqr0tSEqH6MNUVqoBFM
yc4q/x+EQ3FNwBea4dwg4rYwKgCgXWErfCLkhDPuBG662WtmpdmeC9dWbx6fNokLznyXUI+xGVsx
yEi4knsvlre1tfwsusW8+yc+JOSHPuAtjYsu1K++QdqjuKnyvfQiK531F1poRuSoi0wLWTYZu7TX
JB3mQxQ5b16fSvA9xg351HzCrsy5ZriyrpKARLDTjfMT4BajzF/Wz59kLRt0yWX4qdRuUMcl73Bx
pP1BHDXMsONqDFdZjERHZWnnfROl/vCFSqn+2c0Mz8yr40dNU99mGE1snwWmIeUoTY2bRhC8lACL
wi1Opt5VWunolhTzWkhfW74dFMRZiktuky0c160o/qYRy8lzlar23SZY7WtnG4j+NbZPjnkogQJD
tjua7EHK12E1OdR+Tc9BvvACNePCUsoJ96JW704jkpiaGZiejoYZk49/DF+hpOTqyRJkk0Tq+9fK
LvQnjL04xxqky03WnD47kN+BrUuSTCSaGFvxQp95Hq5i5NMiXg11Wg4L37RXmOKQBTNqTVpQk9I9
iqFHg0dIgFkv4ufLNNW5A/BnJZ74G3JDPurzgTWy0NHF2l3mLLxNVfG2y+tl2VNn10CymxDKTvOX
dx80HhsOWWnomady+hQFjy7i/xdOwmMisQVaCWZNEleVVfsjej2PxwUg/tMfXYeu1xWgCmq943UP
OlNayBwrlsd9lzqu6LHgkYzF6Z2Hpk7/V6HC9cg+igcLmq8tF059l0mnifU8oZ9RorbCxk0qtLX/
xuzHc2sE9H9fLyMsUtdYsbIGnbP+JJyObPftqWqBoOtWwwDMvRS4dwOD0aGuAEtJzjgmT3UcRI79
IpHXV2l0WsgBGnsxgnFrGoUBnjafJ5FtSwKYjfHmMoFll6JyaHa4rSJ8Q9qkXK4kbNGx5zOewr+f
hVUUjWUFtfoJ2lZkIDAit+uUPGig0hIpsZNpFlNGJhkM0YM1ZD0Wcmac1zmfwWXYwake0/MJJo4V
aTNq6ol/X4FLRWytsqQiiA57fcLNrOiStE0CFoHaPxy69S+d/0OZG+XKI6T9/qCX+Gf7H5ZEhyZP
hw4InyiqFqw4nemsK57SW3ivKvdwVW7cf3DQhPNZfye8c/oDtqmRLyZgKjOOyIsZUrgj7z7c9kBC
5vYu/KGgd2TJe3PM/QH5OCfihA+TWMioSSU24JNv0sF6dO1NeTeLXC2KHwhCsZNUEWyamGCluP2B
hC8MjCUEmKqv2nC89Q5r1YTg03f7ZIAAJVg/jleblDCk8PSWEw/+9/PjsfVYVDmmqWwfEtHQx3BP
OD/EwPfgvdj/gd/a0iahpsYLzqmgPgO8MQKzcbTLO9TfgDGw3xDw15fW9MvmJM4OOtNUw4s5kD8t
10r5vZokCQ20y/PbzDUgwDizsub47EDL09VPbGfd0ylVwgdkM2oSBf4DOOBavec1KoxBnLQQXqS/
ETMXdT/vjGPLzPfFpXzp+pr4rfefMHXmWpjg+YBsD4wJX7s9nWsvDJOp2A8VYSvOk/r9L8TiCC5l
kYG3ooIa/vnA30QIkq0DUBdXmpV9NTWNAI2UoS7QwnKjVKM40tQxBG1OiGNb4v/ltE5mn0mvTKEY
ytLacSq3msFkaAaGhc+loLvybwYm6u5Is+Khl85lBefgE85TyGT653psY5aJD0R9qq2NDbkRjyQL
cqHCR8FIg9BCZARtgc1I7oOS/8SLbLHr2QSsuUOGVQZ2QMr4ueDvgnNAoL4HXkfIrz6mlYOH1m68
6pKYihHNPxBKNImS9TzF+RmdoeVh2bUbApn9Prb1y/geYm8k/aVsm0SdESOJTryt1KtApLjpn2Nz
VuQm984IE0PPdKd92jQgPZpLOPRD91BF1C3RmAwcB/m+w+COyj4C0F0eHjsCEnCuiReBWhms+5nP
hWUjZ66QHM3zRLj4EWKTOjGMmRYiWjXGIOsQB9Gygce3VkfE+qJ+yRUOOfwduw3E88NY9+z2KtEe
DupLAu8d4U65MmkxAlQ5CFDfqmYkh0sE7RkIlsvAOFhN5TeSy19jKfKBJooXXPeGiJiQ+HCutV03
YTNBIyqrOxwzRlyBb3zwZAazssiu8wclXECRvJfvcGaggx13Eq0VVbJL54lKhAG5zonkMlrF6ug+
lCvpYfAqBREzUhfgt4Y0dinQssW3RBjo/U5v+LK8+F11H/Q88Z2dj/vht5Gawh0JLs5mznAFUWyR
nOjVz67eDAR2AVf9vC+r6M0kZx2XoVt0RsiXm7r8cABkbnR3Y5Y/lHRQOiGrLJPHFqpjLr7//Lfe
EeRdbVXbYqUKqNIvYgQYbv5Bca7zSQvAgWFI36IIFt7OthOh8pkTI0j6uByRnV902oAoKYJh/PSM
jYi18L4WlMv7Lj0wb82wtKbaxx0hA9HDDuqe4rXWnq80KcQllYgaGk1lqWSSb5OuQ13Qj9bYBpdH
fjYa2v984EbFBQjq7NNH4vpWZZqMcYaUJ5uwnsC+KI5yyjQSMM2GyZqRt1b4YSyNcAj5bQKxrpS2
0YU7pf40vv1lwI1+lNcvO6xWDMIhgS4tV35UwLdRml0zHJTj3F4pHnaxPLM5AqKl+WsNdYv0Ij4B
bYMIVvYRzQhOPkWms+r2/5JanjwYloMUNH/b1fcT42Spny5NSUEYWwCZi0dcGV2gGzs9d6rayTY3
Ai5JkraPGItLnW/cIL4TevZShVrchiQiJAiBBJ3PO6oLlOij2MmHvKnOPOfiHQMe71BP/14cqbxK
2DgnOVWcj/0AqkZM4i/DtMD9qwN+eaw6NED+jqBVld+TSMCDsWbtqfB1oC+bsaEh+oC+uGtkiDQW
e1TLu9cRbsmw9PlzjktziZtDx5UtcdjxieFNEwdOVnsi/x9BD11hzAuf25LDq7NYzpmjJXvUlg4l
VUGgdr6LZNEQlEjlPDYIm9HOfKLHT3R5baKgvzS9jlU2PHtOt+ps8ZGcQuJmWzTmPxXsFx8C3tJO
NfTPNmhDpNn9arc5cqDqIbbrJqTBut6KuWsLXa+L6Epho+Yv2hq/iB2Vq9TsunN3s0HB7lamQqBM
10YS3p8jr28XAgz6Devq8C+RHxFcqF2jxMJg3Kcqt6Uf11mR+dBtxGc744V0YnNBNa1S9u6eWI4n
SVvksF+Lhzz413vSZ3SM7kNZBZSJQ8B8UwoR7S1pvNQV+wV38taC8P5b8ImzEtSHeTvnGbwDFt90
0Ml8bZsOk994POdpKWtoA224J92Fx2QJT6arev9eHVTSb9CT5FSJp8vO8RqRdsKWE30rtXayga0x
9hbxyhuKibjH58BNfSr8O0k+Zc3hZbxGV+jKyULaXOY2Suu1DmtH5OTR9AqLO8kuuZ0vfeoWaNAU
Q/bEmgINZBIGiUur19ICBAqWwNQUNp0Rn/UgnOWokNpXd5NDAeOPkPbZu71oGHxldU4SHq71meX6
st4d6Pb7xhjycnD1e65uRH+LT/YQnQaw1Tn2nGzOlYXjtzIiBHtG10dkQBpYQKDY/OzV9I96HOBQ
cD7ZUjROX7v46MJ7lRHLJPPp2jTQ3vmSo8oa3ZVAEXJpSWk/d6EgKsrtK4K3Vx3cVCy1Li579pT3
71hEtd6v40X6H1PJydzlxaGS0apK/8A+5ZKDPWWJfAMmxvfRY/A2gMAmk76LqGiYNlCq9kJRp/tl
ldE1KLYYoa78e6wp2y2nxFekaaCHcFiAh20WIjwM4EHaTVOXVSUA9GuZE4IbQSFr/XWFd735Kl2L
Sn7K0xdv7vHe5uMZRrrCTzFvBz5frEEpV0R7uGiVnCvoynNXCzi/BTYsH/Z4tPeK7DijbVvshDJW
JyBTVucAoj0+vZdQcVZ0rxcH1EgRxIR9DZnqBmgRQCAvnYz3pDjwwQwwE4WWqEeUijrQU0jS6Y0Y
Hw7zvHlIymJVyJAGUrXe6osW1GWqJxcT9d7xRFsjd3UrAIziLArEPYq6MFV2tlN1b9bt6Tztvudq
o8TB4UxJ733qT6YwOAiXAr9BLBnjuutybc0p98dYi0kanuy9DREN+6tJrZP64/ptbzCfTvjQuDkF
gO2tF5d+fiqi+HLWpNXhAfioMuCwQX7syss1YLChsEca8WyyM1l3oS7g4wcQT5b7NS2yTDyqazZL
9kGWEtbha5z16CFUtIG42eyH2Jw++8Z9VPGL2K0vqqMgmYmiwj12qY1B4EPTG7CKMnD4yMq6nuhE
JJO88TTtLIFMLm6yyEQEKSsvVvSUWfjRL3xCiXM/8ZfqxM9kFxmRqsveF0mNtC+L0zWr42OqylUQ
UHMM+/RDvv8lSmIgUZe+561pBofrmVY7IF4IoTCGHm59iqUvua19yX5CoIaQIFTPj48+m7PgyKvA
61aYbMyWLw2DCJD/1S//6Ut/43JPKeEnLGWLCife6CqOL/zUH3QnDRmR/vVGyGjm/0mdFufZlDdE
uQXKEqRltZDWXF1ee08vevHizHgI26TNCIYf2yrvUKAHudJHiatqyQ+J3x7yhRO/fbst1DaY84YK
1aX3yg+PQfRJ2YbWuvzK1MHYH7HW7lGZRNYxeGGR7XpnPjQeQEbBXwldIx7cbu0/LcHjinqHk6E2
j9s7Q5bp17fn6uJyxhwDSg3XPoiTJNx7425lPKCVsxeJddXviu8zsSQnAA/EgOA+zameU7hR8YdQ
yd771egQJIwaDW6kJz0ehomhtKqO1lS7+YSgaw87OxEPeG8mZcCZeHe+EIrsBUOmTSDhcp2xCfe/
QzE5pvy58e8MiVS6dFp8CDrRYRi3BlnTp2Pho4zSEqh6oHSl1Cqvvucg09ttPoynkKhBGGFMMDdH
uklh6g9mVJlfnbi/Zx6owBhCY/a38v5aH+ZSAYUe7Sa3ZOkm4czq98tdicjd8ROUxmB2Wgpz60YN
jnePU+Es7z9vXUC1TUHCQcI40/U2XqrFQdvyWdyG2idkOcHiTPhaMo/WUir/YxdNPw8WtnWgyVCB
THeNOLkDHkDDQa5z6g1pRPcs0WbZ5kI+jxByOZicOV0JfREjt/fhfT9r+QGOmw5BqX2NaAZXEVl3
2Lx8ygWimJqV/px8mHZJKgakAbofqrOYMDTH7OjFaVPH/gsOngRBabUANSaeQYHtdKovnXW94Vr2
ERSjZrtFhi6rtQIqLqeGUABnA02ch8NHk+DSTrf9PZKONciy4AaFzrxiGBPeRRI+BH9VyPrpQSlE
JwO60kM7sRP65gsA6sz76HlIMr1Tvyz+e1PGoAvD7YvDAJkVUo48Fxq9hhop17f0YSgSgbDVde71
52ZErnUq5KEEZzhhN6MzR/ov5Vh/Ls2l/VersXyfXDRDwxHXDX1ohgRd7RPVlIuhZXjsTnkc9bgo
1iJkRTzfxz18NcBrI5bCtRQvhmtBssIf0GsMaekcrQQm/wXyV645eaxLjP1OeC37YlZYJgvv8ebO
BMe1prD594jSH/jbCtpWc80Gcr3iFxhpzYKiaq03cVzoTPWYLcDO+XXosZLzn5og8y+6W/opG0np
mSN8kJiAMYv8hHQwgnuM8Q2xyDE0L9zkErvq9ZgxxTQQpELrsub+SAi6P9jjvs37XrC+cmGVDMwc
n80Y0rg/+hhZj3mL955CsNzEmV0RKaAuHzDxH20CjWTvWm7+/KYEiRlMkn/QDyzcEYPummn2SMhU
tdraHLcNm7N1+5cu3HbcU83VLe+jRshIKqYWu5nc0Fj+03zyZmz3ApHKQVKNELgY0O9vx1n7HmkK
59DoLYgTRUPuaLxHCevFOpTp7NNf6Fm3Eu6CEQWjPjxMdbcu3OyfG3xArEZICd4eHgsHeoJzhlEr
zfobzg/azVqEXnzrSKxYVcpGX6rqNcrO0/D7uGOynw70aMaXHguzZlGVKtfGHEKmCciEn5yjL/JD
a7jLK14cy+wpc6eMwy5mqWjzbOmW4ocP62NmANZnJ7UddMh+25VZn6wzLV5sj48Rqy+pN+HV930l
3kPVyhkdO+he+qTTntemvwCa3GGCPH8njCCKNar6z03aEEPo92BhX1oWNYCzw4oYBgAsUmLBeudV
R26pnK0ZyMOgvj5G3G1uGRrHkqAZ/+DTjjY4hC+rzTzQPlJrEuusdAW0YFYMzrY/0cOzXRdYDGhE
OrHhhdyZkQQo6hh2Cm4S7cjsOGa6CpO5rgypCRgSVDJDhuxEcq+GNtJ/wZc5u/84TN5lycfu5rvd
nf5dks8dKBbXODMlM3XyO3Q9AO0CjhPoG8FtHkeiz8/hy+EeAU1FNqEkhVm43a+e0MMoaAJLi9mG
w/YkY6HYqut8voUQTypeg5GVcYjpBQAnjTqjEzqOupu4lyEMhKJyhZIv1lASg28KyGeYqU9FN5hs
SvnzPjVncG4PNdPP2LAIXXlHRrT6tMDJ7pR6df9vL+QtWPimK40Zua7bOj/iHvNdvWMypodxKWUo
+YEqljj129wsqxgIzBLBetakPXJAlcWR43GK+1Xz54lxmzo1vAf0BwDM3Dn1pXE0UmHVZG6fyQJ1
N81XDhLuYbnnmgk5SGrFW5HRCBYnGv2usv2BUS3dp9jWjKiFi4DJ+hFKwqDoIkxVlsRkYD8DvL+Q
nYDNLvSzH6FRNG7Z7hgGq8TIoQq2FNVOL8XcOaHYr81UEWNklYrzysZGxThQi8s/Gu+ZuAWxuyaJ
VVGZOwgVltlHBoS9OD/hgkSgXoCU19J3ZKiH8/4OtpoSekB0lR1fsDP1bAbgxuZQU1LG8cYlSywE
xRNDNUxE3D7LjvPjjGknpKugJE4oKjNENBSB2FUxLxo+yQlm9Lb7j46mb6UZrRFjvm5aIO7JPvvq
moJoFYIGN5MJwAHIQCaqyXz41CfsH8BuXDvkKjcfEPOeiUYs9m9UT2lN1+f84kqPZUMyCFXmsJnR
Z4shLq7hmCmmQh1M7dPQG+JY//byRjzipf/LWO0xQdUoQycP/N/vlxGgTNgXVddWweDjwLIe23dX
tQLKxVPOPXqYQHP9f+E+gYz2/Q9iNJEOgerjvGcV3oe+sVAFXwZ1+4ql31zvHJLd+KeAOCdxpsVN
sYP579LByZKMz57TD9MkTCRC/MAgqQtqlCOek4f5JA2r75pCCOrFyA4qmv52zw+ebgvucGO1l+6G
8MWy+g+8L2x1kKGgLQLMSvS4hmbWiKCfYb3fYYhqJ0G4/mwSZiv3E7ZmzDmFJTbXnqsuwExGIS5/
9lyl2s7AmThbBGNgpqmoKgnYgnn7NojVAKm4M9Xi7gc+ZduA5Csd41ImYv71xry0yJnmbbIKVdO9
l7bsd4jGi5ZxhpI0zr0Un4o2Li0lrOKnUEcDdpgUOhUtpOqwmFjZTBdmo0eVSYNzhexAgRw3eKd4
hwLK++ERZ9tujYduxTZF7BqNvTRziAHIs/SWwgdriYXjAh9+WjicPyKffmVAkR6IPVxbVmjVHpx6
5mL9TwhMRVZQnoYVuUJ7RhfDbTo27wo/hcr+sX3kkrx5DjxrrNoGl3PWotlDJq6KqYeHRfgUY3u9
clQ37zlh6M83B6QYt3wHPH2HzDDJOo/6yFVZGajT0S83ipXy2stAYzBfxEHZ8j2aKzzRK3gG2skd
vGqzmAueytBQzhr1PH5NnRMKm5xmqHNI5GDT7XxxpUGC5FOW97BW8J0PCm3vTjvsRFHQTyA7ONyn
GMKYjSLIQnbU4iN1t9CfBo/GMXcEipwYrGEbttbDORGWrnHIoaLDA2v1a6y7kloW1rQXuZc+GDe5
H50hAIiGL33IidmvjZdY2YzRKDP9B8y+5LGLPj+2iLlQpvaR+W+aB/9n/UyUl+DJmZww5wfjJPW1
ML7Epy05mwwhgiEbVj3HvUic/V/vaC+cisIQY76uVipP5ASWh/moQaKVZrWke6m0dBzKKpai4Zvc
6hdBdf+bz4rgjJTd5VH6uO23YjWicyh7XoVMYBaqHO6uG0QhhW58zxHNF/GLT9Fuy4cIDe2BvGWA
nPApv2+sGtlE+vlh3NpR9HOVJil8LJA44WkorKvYrJDSaQBUlUFBKK7Fqznc3MtnlZ0SYH9uMe71
hEJKqhq23Vssq7uy4wtfZUs6Fq5iw2yKWIT8k8s49HrZ8dnMUe8jeJZdlcookWOvD8Hr5rtTS9AV
f2yR6OrTcDhOb3k09JxPunN3RIodRp7+K+CDrOGwQoGB1M5fM4d+xefSNvitDOK5XfvNfvzSNfPY
r7B7cmYZBv2INnsV0eoW45rKCfmF8lSU8J/tCowjMMky6JiwP4ypDtaj09RV+q1gbxFtOhih6vX+
OFqx7rA1uJbBc7vB0PP1xM5MWcvEu6VDnBRePYZsBhsoVVtGt+6QeoW7L4pH9uLWgMUPIJW0vx1F
j9qBkFXP9bvQkH9n1eH8cIZ/2bjPDQ6NrJ0wCfzog+V08DP0s4pM9MYqeQ+C5j00aCKE9JhG/+oD
90xXT/oDbdISbvP4CWCqX6S3H24CWEMeDbNW9UMYFTfdbtB2w141Tw0/iZbq28+bcEsYddUBJnd3
rtETgG1C+KPLFWcZGPFeY10AFEEgdNoCQauiHUzb96zORjMz01btr3EsHU9vW9N+3ik0TafSj4f/
h/nR5+YvDUc4MQ4Nt2MyC3EiCOgukZ86c3jdTsSVnJWgqKVI4zo+1XcP9sQLNSvO1PZ71u7XaST8
1L6aIi/gAP71NPq4R5/Z7+yYKPo13XFCaV//q33UYAX2ZANfGbWFXq5gfO2/H5lZa+JoD4HO5mxl
gup2Yex3qQT+XJbZ2nW2zy6MxTPaY2n4Pe4JiLMS+K1jDWLy6G6cCaJMmpYUOFr1201LVs5v7fq8
vy6K0U39ZvAFmQloLDpX1VzzlLGPrJ5LMsBJz4ZDr6QGEDpXq+/yCYg3LCg6edpCqueXJDknH2gw
C3dzigtfvSPGmPXSTQ1B+UahW4pGmWuYFZUjDqW0nKcM7C1NE0afdOdFjgUvJmbRMahKBU85QSrP
RDmSYvSFnjbCaLuhABZhC0Ef8WRiISWIFpnmqSkvY0Js15+8XasJu8Q4lX3Jw+meNku6TF18KynX
b2E9MSIphdfTdxBEd23j3AQYC2yItYXef21A6e6UwSG8cOIMNkV0y/k4uglj59LxP7VgwjSkI649
UFZsT/87gRiVZYjSWXx4WAYXHQ+j3DqoSlQvJd9zwXsr9RCsAb1mn5zZ4glu7/5k5SiRqU+1ianO
91EfV+7FS3C3rK+4dJujyC0pTpWXCPjvy4tK0YuLXBnwDoiwVCXO8XEd5wMYr9EcIadKpHmMrfu+
itOmfA7QIsc0KE4hfYk/VL56My380WwjwnKWMP6q7CNQMqJ+gAWw9/wK4W8F+SIlkhVvliduL948
k7FF4odESiu9hHhTz6+XBiGeI9iuRv9qzX3s2PtRcsHqh9aiEsT4iBhw1ylKXWKjv09AJq3jYvSQ
02J3TgfI0GtbrD0ODkqkZEUuGjPbodgClKzxMzDAoe6cd7TZU8aOYQgwYGcARgWE+LnybxWR5vux
ZzE8TJ30W5vbQDOeGdOhTZWacfOL8Yi/YnkpqfiwB32xggotvrcWsFvoMm5Vg/4iLBgmw/gEOFuA
t0WEC++9NqmZb+Az/uzS0XXbUyBX/fA8hjKM+wTLAWzk8wmoeYBVlFa4rQFQORSPQNttwMJH6dzA
mrY/F5AfvQejBd/kwefnPU1P3cRbLqr2DP6tHZ50rU22ru5344r74QKq3vINBtluSBIu8zQR28+p
yx9IpM236S7cVRDqTcqFISrOMEImD2BsnJXISluphuIuBsTGKo3GG0OSAm6LShEl12zJkcEjRhwB
GhBIiA+JNpAV1/a/lFJLKbGcvJToPTIxHPK53KTQPpUGM6h5f8rT4uSrXZLWdjn1YPU31oQvpXO8
AV3fo5pTYXIFG12EV4/F+QllOiJAsGils9CcqQQA7bNGjybQzIpZUjw/2rVX8h6myeOYPC63igVw
0UqGPQedPNXt1YnoBgQAFQEGZZ+g284ygFpOArp+7s7aerlZ2cM9MGbPaGXV8HQwW0UoFrDdreR6
Hlw+iFOhEIdViq7NEzCwmAn9CesiNXX51z5ItWBYj6MsfSBnp5egW10lY5kMD5+gEMk5kw1hpctd
jfZNdyneSPUMgTNQ6oddHHSjem52bxjoGOMBj8MKcihRBT21RIcOgw5dyYymvqgmVt8l8w9CK/wp
nQOe66qNjS81z1jE2YFmLIjAo0sKu00h1cqW3UkOFXeLYK5lehIb2BOOIrE0IpV/vQPtratGSqXO
4Co+kwMctAspviRNajeI/ZBxF2aqSHYR7lhnhGpFqfqlEnVyY9z5+o9fE/ZasuMuG2Gw44Ko+Tj8
kIHyzXqTBRC6u3IVP9ZDJvmbDZ5nQJIQaumOHQSRwK96bgM8IMlx44LfC5PxfPzpK8cai/aKuJMY
18s6/LRYyGC9mwMNqsXX69rzbtjpQI7t2zUlV6SEmC0F+UEyhlyXrJuArTpL0Y1ijeRMszAN4oEX
GwUQsPHzlhqX1QKHpLOC9CMTonrEsIuyWTB1VvfoDWBU6PO9Hms9qA02sQlIFLrRcib7CzdY/2+T
c+Qwk/nLIDFtUEWoehO3k17JpfBO6XjkLzboS3Vv0dfFhxgPs7WyyYObITjrVALCz6zvTEChsieU
sqgBLSFNGXt0YAZwX8HRTBB5TmxpwRx4i4kcfA2shgNVAr0gQ0KFqRj4bRzOfpIqDObORV5ZxyBw
5UVwBOE0Mgaw8HFQCpfMgYwT9WaW0GMGIa1yCtVfqemp2oRmWHtf+DIsWdLHfudZTsvO9YD+vbHX
0nFkgG9OKb5WtOb+nCqqWCg5WvY5VTEl5sLQVaaQMAPkVLmcLvtKAHX3DiOqCSMabxuA4Zg6Ptjy
AW2pUo264zau1vb4LvZ4Bo5e0plKnb6z6UkRhWC7cZ8RZDsrw8uQL0/I2CcDuZbVFJiP/7eb1eCQ
hKSBgw8JsMt8mVBICk5vwasNpI8QauAMHSNxNyrTgrJgB1iHdCvUvY+WSEbpz1rrxN05xUT8BJlm
K5aRLjJNIC1R50Fi6zANZYFO4NiaCBJaj5Utn+GbLrd+u2ExrkbrLWGzbTNTogXEifYJbhrvnn5/
JdQzF7sVYtWvxWPMhJ0m6vszb8qb2FzMkw8zS6JCqMNhIbFrk0Si2ngOAXTbd4DI61YZoB3C424X
3YrRyLdL3Nsup4EiiG2gQW6knRdIKyBmWtup2f5iOjnx96fQH/NPPBh0dRfweeqsV3FULUAw2HK3
cFD2f+BlveLwiXJaOh4MgALairDx859hxWSzi1rq+dbhzZKcQLANZABTZeQ8asBZRsLArDcm+XhQ
pY7bhJXfFt5C0RJ43c/X5Y5SEGyjf4/G44OmDDhp77Btr3qN2XX6uEIB43h1Pr66JN64wpVXEXs1
b1EgUwNcGeWb2pCVQzs+ViIbVPeUqnkqzw4TkZVCmVkOo7lpLfI3JpZ2YlAJ05EtCFR3GeukLg0h
vZ9CZZs7p+DTEhhFCKkdUbVZ1JMPg7co3TOe8d/Aea/EVU2/vPNtjoB1VupGLgqPkgJOj9lNfj6x
2wLQtgQYV5NBg4hvit1gokebMBfDDBJElMs0Yx3Cj9m+hS21ONoyYf98jjIyoC+Q0qssSmUV3nks
ME9MuLYLflPq7cXnlYzNPiwlqWKI+iMsqQWByRsX040aX5iaKrQ8EWz1BxIpY0qJXjrtdhhkJwtN
wXGZVuJptq1GcZPmRhLeEqVsZtXBOoWlNO6HAnPw8INw7bs8VhJIFrYr+9BqjAoLNxop62UIcBsW
HHcWFTZHaLg8e1B5ba3sa2d/OnfgJhE0L8iF6RQ8QH29v/ECWbRvMLAaJ2D1qM00cTvozrg8PZmS
10C2OJvPdj24tsKgc5FO5hoOc9QBzQ07+dT6WU9FyQ+pfFlcxbEXM5jkiJr4JB3THk0f+pGz3Weq
scPiKF0dSS4qKH6AL0DT/VvsKkaIpRBi8spKRniVRgje5izl26IhiCNyEi23lend81oQx3gaxOYH
ZoSUIiGkZO5afr30038Bk9kCBD45XDEOdqSuHrgKIH8ugGZDSzwjAmdY+6Qr5sZV5o52BWeIyg8u
f4kTgjSmmWKzoZYy0T0qIX1CyKg9h0AJC3HIPpp+dvoSmHtyr+gEcPua2PsZwY/+KCWrLsgBQTpQ
eOu2pHkVnHzEL+OWYiecILNtb2jpdMQoP8KmRwmoeFcBhsJpzfAPojAbowObQQTjUK19/xguuAz2
L2SopGDSqmnFzf9dTbnWPHQXEAPwzPeikQMiLTmNATOdsR/30ayMTnZ4Uwx3oyVuh3pLYT/RDfBy
rTg3/+sM23y/JW86yfwRQS4r6ulSY5XoCA/rhK7VHh33kO7pnpDG/UsVYDceA8JFDWGb8JJMfq4s
IqQ89AR3QodfgDjy1kk3tpgrHdq43ykY0N7cYuf4cAHtNR8MdOcN5DrAvuq7VfPrxk5D0e88g1bN
Fq+XuvI+4nQsbZizL0scs+xwy+H/ZLwaTkOTyuO+O88aeuql8s4iYIhxQlFSLVgS5KMSdUcJk1yH
0p3hiBGSdO/qfHKoTjSbreAw7UnlmXARwzWUvE9gxhvgIiEXBp1C8vLwtF99KGUb6rEZFZGiKzxx
35yaf4xVzVmMURdCdR9GwjdfBBRBtfC+F+HTpNnGnJMryC+BacSAMhoCbqodPdiqPrMsLHGJzpio
ikZm6z6axX/+RaedRkeT8E3XTKSLFpuJgX8cz+gDRNm5yK1CG5GfYh0lYokVyfZ4fnS1+H9bLMes
bmnNKbFiBk+PSMssTWgiN9TNeV7JmeNyDgZrTzZad9eSWu98qqSuIm1EPKlYMKOwGBDablC9tRL6
8pChR+sWvEFfSc3w6OwZem+L1K1uJibu0hPWKESfIDHP2WWnniUJZaI2apEV2Qu6G9yDPJ8RZUQR
aNznFZhoTI41iQo0CSFDhglWs7lxLEJ9mDJgTUFS22+37gXhCtZQJ60ZOFKB1ZgozDnqPwQauO+d
/0wg4R1BZa1NMKMiBY9xufDkYetY//XYohGMvLNsUMgqXos01A/1u4ULxs4ZptvwJqGoAToZVrI4
Z7+QX7sC8vyCcVBnQGaqyDM7DrjBQlBbVKLot6lkPE1ZwAD1hH41+HRQld5V71JUYvUBjrWkSGKV
X+VsKY8UJu4RRwtUwHDGMgDZqa1p8HVPRDTotPLf9YYFXIsQ1ns1Q5vQ6yk7MHP5+0SBMZvCUMHp
SQLaSghxlB7jlrJlP2fErivYjVeSQZ7NjPIaBFfjZT5gGiK37mwwLj5dICM+/TerROVp5/n2r9i5
6axR/4dc83ZJ8bkfbXoJQFQqYg7xexPP3c6XiPrBx3nvQGfrhg8aw36mj4opOtPsd+ZASuHtsiBp
01xjZYciH4aDIreqCG7DCpKQULePUgwCL2PU466VJZZ7Af813v2NidH+RIsHUwp2f76KLQyMb39A
eekrcOW9m7WvTUC2Nso9hgw/YC8fObT5Wn6px7TS1aoruXsOcnJfNNqmRSsLYUIr+ljCutGHHorP
RMjP1H9+dM32dZ6dDfn8caCAlRZrTS861a4urMAdMCYYtboTrhqXHtcLKcAef8rWFsDWl6r1FY7I
U/8HlMTnELkoXKpv7vN1Qd5mpoX0p8fsrXQpGrSLL2VbHrCm/dAUgJAHld7S7z+qpyUK4829PXSV
lqSofW3APL6fRG5Y8KmfeEJT0xjiUsgLieB9zC2iXs/1Tr0rpf/4MOo/Pvwispmp0gWiUYpmY7Gs
jLX4dYQIhKetOU8h4N+U9fQWYDIbHMpVEkdqTa7/f5ltYpilTELAoi8ddQjkMMruQudxCe5wo2hl
KmVkzSXa6okyE6r99ht6VmbgJgE374oNr2Kc61GdYvGbfWpnLGYp2z0dlfFHTZgob5U2PxYDmoX2
zNgOePvNttj/0iAzDhPePWlyCArB4Av3TuAq2sc0LPrTaWMJCPE6wxuROUnlrhCHvwGGScHrOImB
VnDe9PUFyh0LZXSWMJMni40+WghhnKz07cRq9TEF9GQcn5kTwaPwBQUVKEy+i/W/FHPd2ySU1mDT
To0tHfm+aQ+/vzVrTMWVbtLvSWHvPXdpy0nJckM70xCBkiMH9g520gqlkuDBwdaYNzGCkJGQhn4e
myrifHzwzW2LWkTXscmcsfaJFn0YFwuRuHuxfbGLTPEQwv/uJSBPNN2TcyqNF9gcC/TX+kjtZ58E
s6jkqfwU99EZtbVHO5XGMSUEf69nSkZ2EpyOb7TQf3DYXsu0kbxh6diCKW//kbiN9hJ3LIOCXyCi
xSxWzKjuSw8K8fcwx11CqICN59I75IObSU4o1dxJvqoWbnNFLvFNSXBvKQg5VhZQgiQf8cADofPw
gDb1KNq67qBU3RktOO3f8Jj5U0JuWi6iJE2gtIR61UFZiKcGGcwjCwAvxrBfsHvj5WJ9LClNw9qt
1+H3p7jgOUknMOflVjj4VK0k7hP5Er/2Mp4ukN9pb6f4kK3jHA0ZGfbldOm2+rHy4FdQDJzd6ISf
sEZpUXXa2Cp2WtHdmUS1b7l9rsPHRvBCt3s84Ezc+bSZ8BKaRN6DMCTZsW+Yd80CQJEut+0z73tX
9VPPECeNoJXt22R7FcQDda4sBEda5fxkOfEbamwkThA1cz8xRO2CJam74G5mlcyd0jED7D53rHVF
w3T5r728LREXtE8PUFmfz/64Z8IH1LzwrVBvduO80JpcN5oUuAMZUBQIs8MsIJKi7ZI/3oPZ5i9F
jOjTcE1rd9ud+XRLLDZjy8YXYhlwUwqEZeU6VKaI5dg61N5CkpgU8bvnzFHmLmMRTMJDNpDDRns4
eB/ABmaD0FLglmFGOh04XD17BdxemEaRy+wMlxSgrtM/iw/t6kXuh7KfeaWHXmK4DJT4di6ElGD7
RglcSKAgtIkrIoyp6YlVvYO7Q6CcJnoaFAyD+kpVoaRFunjuQXwwHgXgqQEDgCNXBBXPBiGF0vq+
iQYF8lgdGSrADgZsdEfLJd0sKQ5dSllz5OkNhiy4ZQJM2NM1PFMlrAtHdpHi2QlwmU7Vwwpu8XlO
76nHeU0y3wYFvYU568VsjQI7wCs9HjFq0Oybkuo8d5ZHmifWOJKUeNAX5pePb6a3EWpMPIhIKmyV
P0xHVyT4SQWwzRqe8JfVxAmqN3aDzcwmgx9cn4WSNK7wLj7u72j1XjXm4E9Gx3X7Bm1y0SFEWXIj
0JWl3ozcu5jH1bbk/PfO7l0T0RihsUJTRhtJl7CHG16S9GK2Z130WGj0je0KkT1LW1onXR6eNfbl
j84r0/0zGuapZJbwSfpILjRUR/iDRke4S/ZGgU7DSEeeX7y77vFEIBJDG3zd7GIw4fdEbuNZS4Hx
HT9POpdOpNM3x3RgGKMNvuLxXNm+qaNom+W3jRUyXjZjLMaC0od9KM5rOeOIebFrX/ohaZl1WTog
0o6IJoxbLBHlD/oRifcSeIs1o8mXLUWmkWbySUrlzyBBdm2rq/qU74CB9FbJmfGBQ9rdpeoeKP6J
5g/3PoymTd4f56R5SpMJLbCQtEYcwJCSLrpyTOzgGXLKpwI5rpqrvFEgz+aNhFL60+fOQVxCkfID
NAU8kg/2w8zCzwGHgGppo8Q3vo5BOM12ZRXOGCcU+gQTUmzs7wddh6C/GXevTsUg/8cPT27S1jUL
s73+yQAMVI5GZcNu54gZFUvidGsEhUu+5n/JLwVx5tHBW3MZPz7BdVcspjPy7V0/hsOgRUjjcA9z
AXQJrRlWosqKew7T3wwnMXTkvenkprQCG1qfp09eovZKJv29bluD0Zem21AIHFLMUy+OKAED9e5w
RZqmUEAlZDbVg/M1x/gnvvYpgGS2cvK72cCtcLHHAnSTcFfLazarYK7XySgXI0/MEpM3I7TN959h
prN0JtuIthNPnm6a4zK3D98iVTedrkphA+xUu/tInLWWJdtGUuB3y56RC7rfyq0diQG67OR9lRVl
LOMjrHet2ifoulGzHc5MDdlFCFAuHiz3YWf/+8jBmTsOJOZgBNcLemso2Zwex7D73udOSeAyRM/4
Bdxz+6ZXfxR5/6NCySsbZC3HVWRHrjXCASjIMrKAL/H1M5maVtB727BdxL+Lk5DO4puLYvw9J9rx
JDcjewGsk7orjrr/Kf7BpLEPAVjxjt9V7JYDS6VyY2qYgiYh4yFO3PCp4RZXdQFIDb/dsye2j+z0
sXxGb46dpvhr/02z0/Wsa4smDRyt6n8WyMCu9yFtX8JDRWkfP2oVyQVTbpy6HRrlelqWVPUqZntw
NPUYbHrJ+3wSr7IpFq/emm5jlSFcWF+tooiUig3GqqQ7spHiQuR9/NDJbe7nyC7uWeAN/ZxpcqjF
faBTuJogd0BaalkIjfSnPeTGRW+cKISiN44wqxA2IFLXb6/1IArq3Ii+HAxcT4VJDdiOh21j4ytx
XQi3SKJJ8HqjB6UUMVpZhzbQ9b2p2ttADcKPHDn+XBIdoUDKbSLFpNgZHeuiIDwm+UH/Yi9zo85X
Wct4z8bc0JAK+GvHVtVaKzdC8Wxwm1M/scQZ7NIdOUFAxL8DAABXi1Zw4ENJmoILeBb+/JN+Mhvj
vibWN3YdnVIsrz1mWj1vfJqcbM7/8FltZ3glfscaiUAiXeaxSTRlnpWXqwPSmx9fEI96ALy1PqKI
NaOPXGlhaaxHEa6Rd0fJv8KwG0ogti/JKb9cz0UAF90BHooN3nDR6GTWakJGYhqxsL0+2LDi+JQW
7kFi4d3S3GkiWzXZg/K0xEMKNFmUCk8x6PrjMgZOZlvSsto1aIGzkRy0movFr+YvEVFzMCknEPC9
8AJ9r1Abi4dygQXVi3KDDgB538ekZ9jCooh3lMB+Rm2JI2Lk/8BLX+FM5txE6zqiGX40FGaLUl+J
W0KL8Z1NPQOHKdqWHfrLqMy9qm2aAyeP+TYuNU0mbJPAr4CysGu7lOxSWQVnPigiG0mKiLBji1+8
J68h3Do9fyADVoCzPbDFLLo5Msuxog7twpkVfvpD3jop+oketpjO+m+sdRUAJoxYY3+B+APwsPbB
v6ZTNGxKO7Y7b/9ut35h/jPwW6rfUWsq/jJqTcEDrWE8xz1A2m5347/GW+lJ68uoIcOm5ubeBwgq
TYMAAkdk1cBQziPmcBHs2iAXLyHkN9lv1mSidTqUQ1ycRie4f5g22sWTrqemFELkCIkzKTXwN+1M
MsLJGRekSPCAjoi3S6+BwaaMYpAtkx2nWKMw6D8odcx4Rpi554n0vTFTW/KZPNx9dUg4NZhINiRK
9r+ZROY1tGnmgtCMkwp4swzAQXlDALpSIprp50Vg4cC4iLPUvN50mVlA1JzYKhdOYVtt/D8KBsFq
zGR9rvHf5hC40D0wSvebWNnwuvsOZl/Vr32dWEajGi1lIMIIJuRInzpZSQClTBs4Oh2xRL1eNaJy
lEpLw79QxgQuu+2wbY/uoubnqUmzQLXHqziMxTVonF/gaPRJNI365SShJ3Minhg8lMpT3ywKatOq
75PBWTe6et9rqNCg86Qkgie/4JI9GkyyHr6mcDTC8S/RrLGya8nC7NhO2LIxxA0nOibobWCjiKwk
GnvhHfmt18Ki1Bk+/fpp4/X+fkvtzfJkcVCJUdJDgBknk5/zP7/ttVY97A0vOAqPH619A+nXzkVB
mp7lT3wFcrRto6lykSvjEvJFaXInLJiXGXWhJepz0z6lpMhMGGSCXZAecSD1fxkVlowL36fAv39/
aZTQWDPHP79DkyaTZO0nCYf6Z+GHx54wkS4wgsqxejZsfh/VvhlSdfrJdJHeyS0iRccvDF24FKIS
HbNFt+2waxehrB6vs6jsgJfw9Kz5fa+zBGzRdhhgfnAyaqfZ6Ka/yAOs2wFg+cglmbvc/8sXpoCg
UV9jazvLRgMapQf0hMJg8E+0Q8oGo4QmaLoqyRwvWvw2bjjxxxfC7jWPHLu/lPIxy6NILC3tno81
RzJiFLcwOfABE6ayW92J7IVR3HukiR/DCsPANdndOBAH034/LsEsotCr+8Kn3sKUkQ/j7blI5e7s
VAviTtlL4DSAQPHMvM33bqBLyEQ4DQ66Xk6BMb4GGLBLVrAnzVP8hXyNrQJaJd3u/Ptb8rQfZ1BV
UeALeGqdmwPD07bRdQXy/qsA3MS5JtWYiD12aDBx20maPb4H1cIN1ndLusP8GD5V+DDlOzFP8rlb
FapyR1ZjCqnWtyx3U+sbOi7TJDQxTcU/CSqT3O+P1g1/8hLGXZF6iChGvcdQmncnAzgO5SXn7dJ/
eAb7VWhRunovaWVyVjHbjQ5zFwjNu7v0P7PrXjHssKfD4smEGECBqE+j0peQzxn6J38PmvERbfx8
uflKkb0NaExP6TprfE+F3VLy5RA1RVG9rmveD3572c2OKVGYXRk3S2ZtAX2xjfn66dcyIbFcm27m
iKPXTVy6b/KG+rcxKTWCdAoqFcClSIPUZxSi+ugzKCAN6YgSUQi1mQr8AGyBUY5F4gor698Teeya
x33o/iCITeJFIruKjqEK5coqv+JAF9bFMzCvosVlt+sCkpMZ1TTmOatae9TbdxghagA499pebp63
0AZViE8t8pIrxSe3a83NPvitvoUMwfyTtdKoJIBYnA84vLrJWv/odgY2viiN3U4bxZSG5hToQ/L6
XVkYTUbzk3YqjefuFvDB107B1T9dJ5m/FUvmWpj9HOeVNNN3bElLFzX6Hp0EQ/RTU7JW1T4mvIyx
9cuRY2H8+uK/3kw6axqSX/tLH9oUwBahh8E7EZQDyJQ1rCQlb/gnX1YWI2z+zlV23p79QfaeiNQY
3netEjOoVzlw1RfZtIxJHLxkenF8Uc3RfR9/LNY/H/z+i7mDpMFobexWRTfMjlaXdxpl5sV3xCUY
P23z767UL8KYnvjNalqrNruERu6MfXPqmZZQP+Mikbk8Pu3i/aM0PvGwNy35OuH4Z2q+mEiO6dmP
lpAqk2U3NbFGkf/Oqv34CQqijdhQJ2z8jH6PCo5Lbtyxq6d6AnxreyAxH9nMdJJd/lC6auh+pQCe
uysZFfOYgoRXwG131QWU0wDx8orrsUHHvCyq9ZPWuorigr6+192WUsjw5zrSTZzBt+4N+aaw40C0
Byz0yeykU+yuebRUHapW+vpEL4WVJpGdXc688upHKnPfE7OV/E4QTl8D9nJzAoXpP8ilGKTAFaXK
cB2m6uElW2BTf5MU9bmz4ox6+n3O9KY0dsgmKZ3zyJAWmJakhvmeTPmnADD905vDtwoVB9B6xk7l
O1cWvtjKaGhCtpvHseTs4BhP9ivhVHtpJpl3RviYunuiMvyXcWjdYvxMx+GOTPAz9pbPaLNhxlDk
MRUbRZ0TsjpMqCeVgjbLm+v/Od4bUZ6N9PrV6Ewyl7fuSxdoNIvqzNWenQTE18xSyGzN3kRARssd
jnvp48sZKrmMNyaRRH5iaWWEFLy48138rnCRYOOtD/mX+NXN4dd5f2xsvZ+Kc4IOclFmRVPUAagT
YhUT9+ctGyRy1HFrWCJ/hK0Q/3QjIq8cfYXXEWMV9x2BXpqQ6T0zjHxr5TJEti4oYaIwYd/j2kw9
tgAGZhDVOKdmEScfcnkJqCgWq8LmWEfXyT6kRUtJxPnG5FCAII2HfZKUk+0X9VVgXLXHOtsaFB7b
5DWkrsGVqd7f9NQEAi7tsfQ2V/FHx6mEjEBSMPX4DTVtWQ2gQa4OiOSdr7QN+oqX6GS/QgEKjTOy
PXKM78jmlKU8+sR85B+Mvq+lRtRlqV1zWeIcFkwX26Zq49um7289+nKPQ02yPfuJ45aBkNmNy2al
dn/3NM4VX5NvZhaEiHYBrKGz3MDMSSTgh0G0ItRJjNqYDURX7wlNLHS+KPbfBWMs1ulfEna3MwFr
P5w3+GcJWch/NdfwaOALccokT+HtcApUO9kBohPGlYkSjrPdaJJUBNbnD+Y0R6zYAJoWNRRM7bJ0
iXP6S5kbDQgxoQyRke7F6erpJX+2fPZie6TD3+XDvoIS9pN50l/QxHtnJvdq4+dgX27Aa/eFkSRu
GgakfYWoqC51+mMOOwCGUjZXK4mDGSi6t9+h/drDSNczzJapxC82SN+FYAljaEqZz1ExeFULgZUp
07k0OqQ0TeMLTKmcj2IjAc7FjZUTQyxkjw2h0zfQL3pEeiTuN5j71DPQphha4FKEBPLQ9E6SH066
riNvtLB70LPSMSRRk+ul0wzI6knF58gXH8uAr/+YjKF6VDjDR0XFugy1uTqg9h1GWg/jNi3OFOdO
2GC0/CFIAxNujV1fitQR5bpCwlJTiGMnbpS9L61TWn/JTxRVQ69c1j/dOcfkiDVSCmbAFebKfEXV
V4igwS5kILVpO09MQQLi+81Uk4v63NAE/NgDuUXwNEczcGcoMCLX+I3px60L+i2/NdT7+HYw/5vc
X2viRmZUjKLkiQfMCdbdhYa4JtHGdjPtsgq7bA+yaMqYWKXn6NuZGrSW500Vk5YSEv6BI4MXAP5X
4KR5G/NybPc9fBj4x6ob9Nrhe+nbKPS8RU3/CYF8Do14gZvr9dPZ8ogtavMOI2S9kJ9JgtZKMhUU
dasDU8LfB9hMWYX8Ue0wdR9UC/R2cbtNebWGkHxh1qwr0hBomUh27D+V5oh6fFSlbB9D3r1umKZL
cpWDd7A+Shw93TcUgAB6JJZgIxg3ZPtwI+yCqEBwVRQyfVndg5CQxhYOmOkHqhEtZQiWNMHMUZ7b
4RtuvzrMIcrWFQGWZFoNbLyYq78Qpu64QSOCv6jrB3fM60lx0qPjkQZ3Qfvnnm80U58ThV+ZOD38
ATc2zGyMFTK5ijKUq1HNEJ50Go7h6IhTTwCESrl57E6XtGuyEFfHDZIvV0sbiLQoL3hEUjGkiBJU
hINJoMy6DPi8gqOk7W2/JA/z6nmwmMtFwi4x4nEdQjauO5AbNs/KUu8cTs6OJKHgmkY1/t5AMmYX
qFoS23CrZVvTwr/38d4S+tH7OKxOIhCIGTwVR1LhCEF4OZb43S1mDOxq7K+T5FBCUG4QEkaX2Avj
ZlZpYib17bJzr70BuDVdpx/F7VTxjUTaLRYW7H0p3m7+7XvdszQRU4SKA0HzDDaqj0OyzHhIlHVg
x82F3HR1fxeLu5f7c2OHdPLN7NOpcnqEUq/WTGUVFVyOt1+duCJQDmwtneHD8XJ15v+eVUbYZYq2
/eotovDKs20TpMIpYh907X6Mv8dEjNshMSavDH3rjzhXD/R2NE0+Gs03r7slLMVuCWHq2KU5NckJ
4v2MZE0oXpxKarBogw9AP9+6I6Ba7zTTVAy084QYe8g8e6BUpRmEzOILJ1NO+++bg5ww2PF+r70J
Hn1Sb67uTj4JUHY1iUWyG9H94DBpBMXyRdEv6Fy/am53NkgNHjbCnxgiAlFx1Yozpx11ILxaCYSb
OKz1NlN5R2vpMB00YhRablIQ5BA4Mv4ILHEcnGjcwv5vU0MFKVoRO01+O12uCX59WunXlrzyucxE
b1rfTG4IwknNC0/q2xPLxd3DIwoprtWXsWUsewBhiYUXEbBWA0CLUYfBUFhMp+FM1cC7hxBj/NPi
fAG/QIz4sazDnE/JpJGwgEt2u5o30KF5F0dFNF4uTdszgFbl6760uz7B3zAxW6DDmrp2Rd+xiDhr
zqEFmgBY5vZvnKVBcVmmgLMcUI2F9QGBIa3tMMsUbAm/YxZXQhHXUYQ/hjm2QmhUCBaGiz3dsDu5
HgOSV4ucZuMK4f0TDEoPbhM29ttiWoNJ0Oky/qCwKdBWBNbkKymLzWeEj4BJo/Ytw4y7DOCgCSkL
A8GrVnXCWWLbMGLMd9yujJY0P/Eh0219q+uYq8twzzLLy30miNbVEOmhYlCqORYxbVONZ8JKD9oG
lf5ko5afvpukn6VWvDQyDasMpfsHDq1yMPBu5trr26wQVOVgrMD6cQHxI4JJM9vvG3nuGTNRRQ6p
C+2IVCS3hCxP0AJyxrIXwAjuqDfIk6iv2FCScQhWhCxKqzf6wVHu22mvwJPXgsPKLlpVzPnQ7ngy
RH1dWcPR8DLiBjazvJ9TdfnLZxO34cob3Axy3WVrcKR4JRgBrekh5Hceg9hZbRMQ17r8TH6E8ELk
LDPAcxk1AeMpUWy7s/3hvcGGYs/hsnWDDcbSmQD+sOgU9I0rkkQmFGcScoZRkb6nnu5cIOoRqdxL
sgcD5MGVDC7uEY6TeOrCyN9t0ymV7YYaAeKzL2K45s1JZrrmxotJeIY69DqzMGKPSgOQJ+281Gd/
IutLIanlHu+rR22+0Q/3/JG3PoUonzkKhVIKyIL1qiEsMzkUDHuFiVPuNPyw/YR14ZBp1Ziq4HjL
OG98BJrB1QcouLKBpquLSejB2rpZXaaKIP/TdHVz/MCeUQONTPOSLwdQ+3KIOwj3SHBf6pEm4FPQ
zGF35DxliFQpN0ntgvVR4fcYkzughalUyUJwy9IYaaCqhydMC351euDZW1xJShvp/Rf440qy0R50
8Uj6rZeNYjUMTxJ/4sIhdHswHBgFF6eU0olJfE7Vx6sCPM2QwLEl8PHPix73d0ebCAv/zXpFF2nc
vfqJWf/SYoTxKX0YVISDztBNRk8MRix5Jfp460q0zqLo+E4rAvAT6IejP7mJLLAUhL2KcpbUz4iO
ZCmA7vvb+tUVVsQpPLiW7og0YPKFG/IzRuUG1KmWoq4vygQvZB4D1cA11oyZ+A5+NuQ+KKmmSCCB
ackBY644vkXCL2hkSxyTJKLJ5UkeaTvO3OheJ63WfSUXFfXo3NRdOYzfhD/ZY1pvQQOjf+JtkfFF
OB/RzTfIyLaROdPbwQvc36QMdLulGWcFAsJ32DZBDzZWYsaxe0qwHSj4IvaKCOqmL/W4ZenpBCzk
P9GSitJFCGf+Pc84xhJVA7q/sBUTqrWsdYbDOMcbkT2znkExHto810nzHtN01xuspaveoQPU516R
Wnqw1afSGgThyLftBoKaFEGV43VGtnouzuhSrfc7mc/PKCMGFWNHCJl6us0z+lMxoj36klSrAiwV
eYpqrkORV3eIBFCoJJ/NQTwX3bREuwZDBtyVT6ZabzuYAx2wvKxEeLOH6zEi1ZVUzjVGqTHWvQlE
QK4qC0y80tON+vvykeXLp/E8LO3CHuetpAcphojrFrs3tayJ519qQZZRpmTiHFRCIPVzmkL7Ns+/
UlvbGNXpezemELGBZXjUfmA6RxKbb+gUMgc+nBZES2omeOO6PUmIf57TxZX42/QfjF3JN0DBhvfK
GGU6FdB+T+KlJQ/y1QrlN2qq7z55iVkbUShKQYO+2D/HERAVU3BMx8xpoZrE+/m/L78KpEQA4itj
jlMVSrXikTaohlasNJdUBUey2UgnFxoZ1M6cKwG5BNMgmgkhE175ts7WbPXl0OrrDqdpkLXVu7YC
4xBxuExN1KkYH7BAEqDacV5o4itf0Xb8mUtTghwD9gYR3H3lm407iNn3Joid32+buWeQ0R6aldc4
bvSgdglZXvUux42DGl5HuUNoTK07tmYil0e59cwcDONpEML0ycu3EOs/984R7/95FQpCXLlGpSFn
3wFuSUGMpmT0x5m/MWIpjG98087ckUogDh9K7b5dF/2aFoej26Jdbu7pLlvvNvr/XHdYg4/LKAtw
KmdmpxF69Fe8MHxsnD0dR0ZlF2STig3MX3pFYgDUN9xOCx7/ms/uZGGIrlgpq3W3nIUr5nr6EF22
+dmc23km2rRd0tdDGBnsI2953CKEKT7FNggf/L6CKcUCHC54CewdF0s/2MmxdoTpbkTpga6eddXa
Bx3uNzwogmI8ucXiijVTUMOGN7eNWqi8z49aWWWI/Or7aWXW+tpROAT7XehnxtC1vM1xV1EDtLCy
/S3fKmPQOQemnaW41UQEGL9q6zFti3QZeVCdOvx630ctxN0LYgGqHYy/pTSHNOMESylOJVoSTxQ+
dWbEa2cpdJan5QsvOi30/nWTWQ1w0k6FT1qeAMB5Wf5VdL6/5NUEn5AbQXMjyNK9e3J+sr684ARG
kgaA5FKmp0TdKYGyvsmnbz8gcYuCwo8q+zt5FjjUkOaZJ9zaZpEy50Y/Kt+zdeyZi9rBzDaoc1yZ
vovOAPXqfrOxVfvvpVz/5xvujZTerwb5nU+6iQvBso478nJS6YRM8uckzQS2qjmJKzO8J4xE9pSB
8HHPya1juo8NNoQjgU5nWKcUUpuruppa59H0ldLGGqmEcqCOUpYOICmt5To4jA2s7YdQEraJuONE
Rol31mmV56V8dsr6o/sdlMVMCOKl5wvzHsvxfalDRtVQwHzGpwhxyhzr1iuEwKkPX+Law7aPMCXH
/MUuz4tqhLMn8sgLvJpqS/2ahtAd2/zKQJ6avsh+MT7P2cWAf2GsFbtxyCrA7U9OYCJBIhDyQrTN
cpkxpqrbXjTOrZ5n0rl4L/fw818TZEoZTdkyv0ofXENQmREP+h2YxNVnsnyVn2KVskeEL/6lMSBn
ijSAShCGqaLDO9Pv5rKGwtxryKnwVUvaVdOFC+MzJcLFex2oACZqNw8i/48ZNXLqHJIYAs/5qqIN
5eV+ao4yKFuEhnDISRJGuLb9ucmjQR6fmzNYpoUAvJfn0H2UDo5wMVtIJyJZjP96gGj44b7MEQNK
GvQhYgI21/AnTWHi0qLkx4gpa9toVHW+0O00Ay4cgCfp9+dCUfs7/yJ8fBha6u7DFDHxcuFYvoi7
S/gyHRrrhINOHt8bFQA2wN01oeLtcraibU2pKqIoNRjbn1bRCaP1Z/xBFSNJCjz8I1oDA2B66yKm
GLkrnraXJkcKI6z2C79VMYB6rpCEBMaFFEdpqk6oRfTe92rpZ4RDSXpInvIYS6C8qjeYNrU9G3IE
tki8ieN0Y1JstpiJdtrUECwDROjWRIZnSuEG+kxKEezldxZTS8OYvpFDK/6Diz4sUnYA+KI+ieQ8
etSaSZWXE6KEBs7jECoG4RfM1z03cHQLOkQU2Ib+NJGEWirPK8gATBVTZuyXgv3J+dX2w0la4Qlu
XGDrwa9En0K3QY7VmL45j4PKRMUVTXRaXGncOrvSkQP59lL/DQw5nws/9K8Z5Q9t3y/JTtv0w4QT
2tBZKaKjDZYx6ibdCyJG0AcD2PVZGc5Pf4p0+i1olV9ytO6t2dV4Beh0tyr4SAI10zYgID7g1vJR
kzi6bXy65qJJ58Wd0WzYQ9m4dprBmMpfn9DcYFC4+Q0S7K+tNQ6L56/uz5et4P559f2VtW91o+j1
WE3i5vz8ON12V3uLLkyPZxL9398rCTqfbMTJkn4bkSFxt1Gk/QD8CORaJVzrDPXI5dHF/TVtAPPZ
ymImNpuB1CB8S0rePunTxSsRI8yx+K5wLSjqaodEzZFhmr7raml1a3Y2TYAL2EDwySBfy21u0+6t
zaTmyt0bJ9UMKucU9XwvQYcdIBiUDJw9WLoq2VnTLHDi62/2QcCKojTq8ebg2Wh5dSxM6bb2gyP6
/fIFCSOY0/4eR2JGbg2AWRpq4e3mKQmXqvgs2gRRo60Wfm/rw9T+G9hSxU2ePVBsFYSB27aSaeNg
duY3CmPkkYxFKtEZ10kASueoQXhoa+2AoJJAtMzjd/84vQ+0ooG4yLIZ0xCJ2Aw7Shw7zbl6nHw1
k2PWL0kBxA+OFQdzrycq+fE3WCFcZOwvjuAjYkj4qsz0l66ShJWJijEnZXT4C3wjqBRlBI/XvaFD
ER9glOy5suJU2V8hQoIRUdefjyqUhbTwfZ5xEHrKfcwd+bQlaxEfGyedNItMkGfIE6nWbwW0XFbk
JGcrP36VR81eIIr4vS/mthUntgobBsDXo39dRrip1Terc+TWoMNHYQ87Hj94KMKlJyGAMkvzCoxc
g4XlSASUKZWl8ft2p0Q/r0SEwfG0xBT5pNIxSF9RrA5K0KErJ4/sgH+Xtp2T15GfD/VRaaaCewZd
FjCfAi0bAeJE452WehgXdSlrMylhFfR7jqFaDP6YTLfSIYKqxmAIBhxysahI1/pspsr3uUCASb7Z
0C2NOGow23MjS+hU/K+9kKhUlEN5EpdqGVNb2U//RDyBVOymEN3f2UaX8EKnAQdC1BBZEQeGoHqg
NXeEySP7TGPkNINOKqgHwzXKtnFcaQBoKXHgkXEhiVtA2dDKJ4Au6uiRmaGLT3YKoOIK0swt21dd
UHbvjYPmIB8h4hzu6F4cK98qUb7ogE/UsrPAaF0aw3EgCBuw7gksQrLbw2PqcqUVnU+Y2Tsy56V1
n/N4o92RCOi2St+9S1Edqw1gKlpaLN+SCdyf5QiZ0C0BYkEm8fjDqLGd033kjwXv1kglKnsQ8WBb
9GZRQc3RDv4nJymYz8SHvlq2R3SzUatrgLRXdvNT2S7XBYJAKAx8B1dHSYxYdVW229VlyZm/P6RD
kEIRlXYmMkVpAFoYaXyw5S1L4FriJd5N1ys+uTaNN2tTg3/VMSLfJxNlYhJFB3pd6Ecy6dy86U6i
j6wb5MHRTRKn1MoEOT1QbJyjgIEe7GdIM5q7xv1BV06xdWNSIkyhjOw09JcrYRTcSNMxh9phUHYD
t+v0MTntFMA8dW+80O+mdj/afuFgwP184l1GYQRf6H6cZCMslGIoFKRYZMaSazAuaXbx3u9PDetE
+12doPAveBJn8oJ42zLPsT55vgDyNklwXKmXgTo5M9sj1sOOgv+c1ycxDvJVTsbCg+ozB6XX7iUD
8MauQZTteaK2MN6MbbDcZSgxmFAJM/hhAUsYWjq9v21p/a6M76asoMOfPQPknNWqizB5E5JM06ZL
kDo24YSGq2qnOqwkulc4m3kvtqwxY370OcV9eiugLPuCuwZGXAl3JZI3UkgtBDqiS7pYoxfXfs71
jwb9h2GtaAmQFkKn5JWUoT6sWvMzQFqiCz39SYtu4mBkFWclTTNN2aiQY5Z3svU7I2masFEMx/8o
NVECzQsrulslaext3mlq9ZKs7nz3yXeeP+caUDySTTPM7vb8jBtCgPvEnWD9Teo92lIyUFHNJnjP
lYqao6Ybgjq8KKfC865cXUOPrW6yyNvYAjl/LH4set+sCGprBxZkUPq214TESG0VNI+94PXzRh0B
gNSjjIZ9v63eWxjEGRc1cIkYqhPwwL9dr7lGPjAfTX9RexxmLTM5bcOpDreYQQM94JFFjJYZZroH
AoSjpGW3ySa+2pnIePu5Lw9eDw4se8fP9Fk1+EYs0cqZGw3vXYwmcjIUZO2xx4NJfG/yskknbwqZ
V8N08oSLZy/nFxDfgjh86RmQC1sGQy4uJGkobAhbgCH7Jn3G8zY1iXoILnKusmifm3TAG773t6Zf
WAQRv98Qlsl0Hb3Uy10AlW3cOE20SRH3KwSIMpSzVi+fiPJIN2SeyIl5u8s1/OwaoF/QmtsIbcOl
dIC8gy0hkMKYnlM5ZR3yf9zHYSyDkoPEIFPS9fBBPjil7YorzrKY30eG0rKKJ7akQC6WZ0zHpLpj
+VclMaruG1Witq89yPmmuj66Wop3ulIUzDVe53DscHpi2gh9WmHs5z0YzRhdwwAZPBMDx7QB7O3m
ajzyNUAfi2DC5OzB00j74AUO8mPtDzZwRswY+qSgtUCNzXyXrxBYsiqvGj8eOCULR8kOyvpt8CIg
CGeKfIs/XZPql+xAoADNv4dFot7s+HIRueC4Z4X+NrOZyCoSZmUGS2ualm10J+ES9dKZK7aKHa7R
6EHfoNl/RH1YSC1MbL4a57Jy4YX1bL8/i+QuxLNKjc0Oa8bA+iNMB+UjQj5+AA2R+dIYpVm+1aT0
b/PoAOS288bEgfuw4rTy1yhTGVPedo5GQ2Ry9YykWaKo16ej6TuOfqUbDNzQnaoeJ0ROI7DQhIA7
RT/CRYTNlPSxnItIp371d2pJdHwiZ2DKPghh7tUGC5qriSuHN7gRCRu7dubb0a11VQMgGTyMQftX
qDj9yXFk89q35gcZgGKZ/wPwASKHnP5Te+XWLYdIZMg3ZsVEoxBWa8Wx1VSoEIz3cjQ+Omw+aH1k
n0KbDYiza3hq8Jl6yDR7SnxYDThVvx5qwwG1hCnX5Fg5lgJYcE1RCZ4Gv0Kr61pCFcFifPxoaGKK
lU7UhKa+UuCmF+Z0pAdKHJXkAc0GGOvV6ESYRjFhmQY41HFMNUFzZZwiylSNooOOBN+pJP9QvNT9
HzdWo4PB8T5WmRppRpD7aAYbDNAdh9pMijZpA7b/JsTkWOLez/Wyez0noDKqEoMVPYVZlPSVDMQO
IQTWQA7rAQWwi44813Y87f9cBcvXUuYBZsbJwt90Z2XnkcxqC7YwaulfI29uM0oy1ht6CPweyHC7
6BYNUPGy62oMtIBguUDHEpm4DCl+G+uH1vfyjSuwJ3JxFOB3lgqo71RD+QuHyqUOL0OTUmw5CEv6
0TrtGaJQUxmKCJSeS8PwdG2PrCkW//jXSMiadZM133UrUq1YNCsCxiYzfmArsWImnQTnDCIQlmN+
Uhkr0h1DSXHg1YE6iLVjnoadHJ1HKRxwz+dm8KNnaE1JoXVWC5O4rmquW55Azp0nHY3VkmIp6fXl
aWzuYFjeh1SgyPj9cEmdgCPVNMxI4csQuFXTv5mUBT2YbfBT7UsoPNSjLXejl38ZzKcD8BQgRm/C
yKQGSIvCnYY0GLDO7cauTLhgIDu5CdrqaqMzHwYEiVqJ4FYxdnZIlbR7PGx/uONiAeJ+pT2TEla+
ZC7EiDkcI2WkNEmkj8TG9pmp2dh1aYsnj1mcmQObeRqwtKt2vFGZVCF5YJ9bfHsVqLr2zrc4TLLh
TichBaLVrg1iEbZ6XL98DZps2KttJUKBf6sTEO3xJuwceEsr3viyFZxyc93+GMCcC6RKmJ5w5eIq
VhpcgeJgUH3xLJ8Ny/Ar+QITob0k9heZ+4HXOMW92ikbMdziTvRT9uGgyXNBckHASFQcYLJeYxDj
TyYUNoT16Vt6s7ien5TcTEcW8SiGPtDsfV3AR1PIqXK7b1MSDDakYNbHbL+k3V6U7pqBKTyKLu8R
MimJ/rqqGPK/91+5vE8Hr3SeebdbSB9BlEZ2xgIJc9I0MY/m7BmXi2FRG6W8bFvSaUZqO3JIIUhn
+MiLYm6lLM4ZtVVNms+3UUgZjH85MnQfNqgUJv/v5jRYsNXY0gopJqS1QSxUP000YZrSo28BRyXT
kjK5Na9r/cNpBRTJOE6ZXqoKOW2S+E2yMqQtqfoZeJo7w74nCwoKYJz6FavZYIkCFgDDj1TrsXeP
VmaUkO4F2ygw7u7PcseOXmr+TYV5zdDEa6LYuv2/OZR93IX/0GXBbVPkDVoLgwO7ujsvUaG/m+SC
PdberQ7LKX3XJhnNQ0CautHxG2XJOw7C1vt269ozJgf9pFD5S4yNEH3SfoJ+aTZxGv2qXud0u+Yp
ASo/c5Z+Vt34RCNSZmFAfLU8IFZ71DmjlS5PIQjtD1vFXkhXp6v8CBHgB0FhFOT7iEUvqwd7dPMD
GIbQn81kcztVum19PKAcoUCXBmtaxtd/GBnXIF2gQWq5d+rthSk+zrJwYqDjKTcekVwiZA6X+sH7
qQga/5S7zwbHGpLfOxIvhJZ6lHMsWnUTYmGcIxBapm0a2Rp0y+7k4BtcvQ47MwiEB34QY9/T0gcz
xmTPW0ZSCzIykZwNicifo74wDANn+Kp9Ugkjgu8LPfLEsksNIB/Jxu31N4q/l0z8dxOLwuT8Jf3M
7FY/8l8/wFqtlInVnJn7ULPuwDPd+hMgLJrMh4EFeovyIZWrS/yAaHnR7r9cAxuNO2IrG5/Exhkb
4d/IDNUb1rC3gDH6KGE4viYKDDuG5bSC32BGCNFCKPdw5Bmb/9aT+dQwXkwI5Q81A1scZcgsze4d
jD2mCaJWMacw7t5XWewszKsIVFjMp+NLEvld9eJD8XoFK0XhPv0dJozH2vxLfDZW4DL11yoGn21F
ItZ+Ncy5ujvQFAJQ7PE9fae0oKhxVTh5M69sjGNtY2gH1J968jHLvWCbE11utzmbZE0uy+2FvNft
1rnuLex14TEPN9W0n/dAHNL4nVp2uboSuJ82EGpQiQnYG80/vzT9fx8yFkBMv9suLPL4SY57r0lM
tYUIVxlNRYhwXtu0uQd26mWsWxNbxE85YE1FR1Q2ZFMxVaWEEwBSXpJ9qlSLxX0Yc35XDW3iBsth
qP96GggwnTBT6Q5geX4jcpkAHmRKghMI9MLc9KhWMo8hJqLzWpdn3rhwLT/KuLzZuXF2YU2yLgvo
c0MIhA1Uop3bLCUYTci4DFMugVEMRndGotbpbQncG2EuCxSwLOFksRhRM6DT+u0n1D4XcSTYYU1T
+U9a8lWFeTbo1RVAirYkZT2s6XQeviYMN+gXWq/vgtFk3buarn8f4XbC9rqQKfgFRj0AvxZ2Fe/4
QFX2KNW3y0f2cDFT4UEitOUTDSNIdI6ftdI7GtT73bCSTMzgbjwKi09pl6Hf/q7vb4WVJnzbmJwr
PGnVMSymmFizfE0rKxZBXpIzLQhdWCr7obYVGGKcTqPL51up/0vkepSB0CIlv6xEdzCIfuJtgBzU
IYKeK2MbFLbBET/riZn+aFWOSBXT7121nSKyHEx3LspLdli1+dqej+v2AfJYZl5tMVUOhZQyJqES
eIei3kvo0Vh6fxZDSU1oRx2cLJPnPiZ9S3ZI5c7mVVPgV+dewk7Pinn7oZiuX49FXysuoolZ8jQW
fQ/i44vB64LLTd26nKl/AT8D7oQ6wf73+Ng3Y/gg6YjHT6c+Z1X0++43tkLiK/3eF0tpRBkpxx2n
Q/KGPrXDI89UfQDwkEy9HJmd77Yz5iUCFPSdz5L2qXk6XyFtaBk31wj6zHH4hOSp2M0VRWYqrapc
ir4Cpke1pMxcgAtAGAbD7U7dS8p0lB7teakuNVQTeMM/NTxOGxydqwY1ROnSLvYiYzHVtjMjE3/4
etqF91QlaSAJjszvUO0P5wnC6RQGFEA2TyCfZ9uPNZVcB9QNzF9PHUlAa8mT1KmPRNwF2WDPcwNM
Hx35UVbrcBwf7tg68pYR8a/H/KoBXvatzvDwNI9KeyFBY1+DCUuH9vYQ2D2mlA2C8q1h4RZe0mk5
ACpqOd9BCNmiizhTMiYrCBz+/RWHKzZ84xfMBGuxHHM/X98yTSff2ATfoGmRJSPM1QZ6diIevhXp
Q62K/Cf+wq8UkYnsqQhU/pMwUzfXoz40gXFsPz+fDFJTuKDUCDgsyrzl1Q+quj8wt24h+dQmJKsT
E05++xXx4bBetvZKJgyn8BM7A0eR5WX8CGdOCwwwZzTKvytA6cfGaDX/yVo+KNEYw6H2hliqEKz/
xcuc3jAB5mntJD9pq2wF5dM4xGbihosdEIZiHURpxfn6GeI5TLqSjuYD0N0Aopb7gyC8o4mJlgrZ
gbjho3QjPJv4hgT0okuXu4JpkhOzPLV5DRzWsLo7q3TkLjQET4NYNeeQ+KB+tKgG6iXpaDW/t68C
QGdPFpIqbdFZAwP8xm8Z3ySxz4D09b1F3y+96OCKwZASNCvaMist9E6ANCzh6QS77ZQVayU10M/K
LuT6uT4ZZfMgauXEvynr5yXAdxkMOjrLglmYO6zCbz3zdH6zCSAXZzz9uauvQaZ8N89TKKx6ugjZ
Pav159/lMQuiJba+qdTcBJ6u/IltfZVJ++U74COgr8J3TFryJ3OklpbdN9H9sKKlbJjanZvlCf1M
dleKT2HOUU+LODQFJ+eU5lNlx96MaKHtEvdzkjZ9I7jOV5ts3cuK3ZElEKtpUywYbNCLyqZedvrv
q7Q4QySpjOi7zbF1qK9D2pl5787yEx4q2YppwzYA0uzV7SNbM30DyT8ye5EB+8pyxoM/A8PDunDG
WMmlIGsu33kB9Y7HXVrhSf2Rk2PTK8x/Qp3lPvOtadUpjAarfJ3TOOahDMXKIrO8snzexke0AvcQ
Z/hxa5wBT2FJUFMNmnOgzDQ9AtzDC+Xc3piVHBBD3vGMIplxxkqev/9GkbBJIhyPOtevwrC1LwHM
jQnW2dcWHXOtc0TJggR5BQcb0DQLuZxhVZuRqgO2J8uY/a6tuI1VDCUaWV2aXz92Y36e5ctfoxSu
k1UsRsBPF0BB1DmLwuHTx/Yd4YxSSzhmTlp6RX65aMZkU1MwL9jVcuqI+HAksD92P9NkRVoKQtGy
XtkFjwSB7o1tqTqHnjyrtWQfgQ/tUgINH1nhjLo0s3FOQEK90vzycIqdVr1spomf+sZ6hVDWD7/P
tRcKV+W+mCSZJx95EevWU4D5605Xv4+rKg5U9P0kJMNQIaErXWWvj2Oa2dehMszxxYxB5tRNC2ck
jXe4xg1Tt446waJPiTs/9x76jHVgOKYto3x5JNYSx/WVcib6tmW1ga3yvQ80JmNnBt+oWa8i/rYi
orxU9E0aC+Nqzpq6Tpsi76UiltjPh59QZ1tSfrYbDWmEFPbuxKTF6Rg74VyJItE4PVd4iFs4UW0+
0Yfdm3WnbsAwxgsD25W22tfwSfg9NRBrrHpPwPpxzJbGq/tfkAZZL0ml6qF2lED8uKHRiUiN+5Cb
jKhA4zLw/AscGCqeo5EHTYWK7WEmifWTcVS8EbdQntswdv5w0rmv41BbLqPvjqfc6wcaEnfzvhau
gLJYpOnJNk2iEun7IAR5Re7j69ehYbEAdQwzamhHPmiZGFoAZzay57Q+gtRE20/mw8no/ArPYW+X
/YPIByT1u/YdqubUXGJz/6I0ediDhKO6WZ7LO6/sai1ldVaOGH8vuUoPj4RMEXWgz/9ADBv8ZzY6
nfXmSM34KpsAJZIHDC2ruqd4h4cgfXhKwelAY88WD2A1tCK1pAEjVoh1Q5IS5XnZeaM3w8AslM0A
MrxmnXJ7P6qEZ0PFSaJ0g9N/P1mW6wPt35BHr0FedMoIu/6lbyEkI0EoBbMz3y+xITxc+d5ZLGw1
2YZcRK1bTgkLCF4lF140S4zcf6IdK1Zxm2Lq378KzWam8l8lblxF0BNM1PHyZuZw0Qo/gAT4eDFP
Qw2drj0xbsgXXESVYR2XrBGXhe/ejhQcoNCyljIpQL3uDiLKnY9QSHpPfxt3qtjcVN5vfNulSBTG
mb99+DjosiUgpZchfw22INTrCuAU1f8Do7v2Q5O+u+L0qaNuaZQO0yMPI94yVSXGuRbmTW17gsvx
TK0MDllmLE3/DNXfsZtjhl6KyNQEX8b/1GSrTBq4/4/h+ZTr7HI6QGsAGAGH1H1HildQIu8YCcpC
q/eYn0BSaOfGQozSqButxgjwGdGEAhLK/KPDi8O7rTner8DJQSwOyRj7bo9nxW/5RWQPIlLoybY6
QpaJohedx+MlC7Y0hU4wUa0O7myxCe50RigBSRT2+tCIosBsfO/L/GynN7F2izkTzcGf66XKOhAZ
0emyprSaed5Z/rsF+UXbD3OqWBd8fJbp/4hDtkQlpb+qkiW30eEK6lJuxOyDmWbOuOVKY6y/Zdfp
h2pVl+RrlSAo/Z9E9d2SLqDe1a0W+M7XlvTGqz8FRLv8BYRXt1yB2AyKo+zd2pQWhRgYr0NwvV7V
Bocl4aUr6Fd5I5uE/KBZAqDQIBtEaPC19ZtpAL2T9fgIrv5JcAyPej3VDia4TeBT9ArshmX/w9G4
vJowV3DHK9jGqRTHHvedug1eXLu8YZWCjxsSNoP/1GPkcnFxnJI3BiFzIt6Ytyn+bwJhTImnGs6H
ukk3wL3tG3yEfw6wmY5TuZ39K5pSCskGZhKn7maVsYZ3nu5PHE/OR+wBnez0h6rPDuvLimJPPUoO
67ayeDdiGP316+yCo9TicS5yXMWcjrQ13kICIDc3gK2lDMJn7eevKoMFOctzV52zS84NJycBddYw
FPzmnz9SbPnXMsUwVl2RFtHS5siwYgeUQRSNX9+/YfwAHUuth+PdfUPRSLiQbwLmtvIS3AvMShWA
qfgCH4A1BFFQGybd8f5zpCAYP/Eu6T/afPui86k5oIh2DuTvWf1Yk62OSmlRTZMlIUk6qZBzxjYG
S+vMgmVLYffWpGFSPBQ8I/AqPq1aK5VDQunUDw+APECl2CLrJt7/s+U5bj/ryGdNxuOBoB2U9hg1
f02DDiTLgL2prZ77wS8PY6Jd0xeAkiHfAGb385b7w36sh16VGiR0GgrhteNHGXzuzXh/jTq1ZLBn
3/bZe6rXdgTvQh3Iu3OgT5sIJKnIZ+3flnu3qGrnepFzAbrtizaIZDms37pTUYlTaXGXc6Xq0z6n
dOOURzyZG2Z+G0Dj0xM+6SUMIvth9/qwfh77D3s4ix1FnVYM77B6apwRGQu9xD7H3QMCNAq4JyNu
61X5sPCsc9QImSQk5NE1EhLizFcXhEvTZmL5/w7EUx3xjcoMWf3eq+DaNRxvRFpF5fmDceZqLYYt
Jk71I4gaqnyGhlvG0Ypu0Kh3mWCe5E681JE3/cV6PXeRRWcpV80JEDWRHviRhGJgWYM/fjokk8jl
4HRLPSfREsw8EOPiwfWHr43c7tIcWoR3R8MGMHi6PIF9wF25bxuD8EUFGrX7ZdAWSTU5iebHkxGR
r7t5FW4njn9VJaupu6+11xWTJr/uS7qqn38dC31jFAraoKR9Wl/r6P5jaY3X9Kk1fpPd/ZDu1Fht
jUjbcp1tcYuoaLrxszLzT0rCLtXE+T+OB8SzblWJldOCETKXhGRSLmagRRTjxMOqxuXHId08bKb/
V8uaE5i7/5OM0po61Av/+KkwnRbj/9L5DKnaP/XTAsolvv1IE+1C+kO9LmNxCFhgasiSsOGHb+sN
IXrpW+XgarrPmMb2T2kserYiPnE1MIt+dJmTbW/vvp2j/eEfTgECjA5p84flx8HohjqvBHAls7Y/
VDxY8wyWwDZtVqy1Cp96c3mGsxCKtTHC4g7muWp0sWl5HPhCwpz+Orlls3dqAtxOpB6GXzqFI2tx
rKKzxpYO87jizsuAzB/v3b48U6ElWGOHtmYqYhWNPg+BnxlGHYOXzSnv7K1xLITr2gJwiTWo4Oc9
ZfJ81jG8+6K5ajgL18YGhexEjsnp+Gj79K2frvXiSXPATU0cVmcehI92p8n17nXMfc8khhdkLhZv
1txhqVZYZN0BRz3pPjhBPV+qQWAuKkmZYiGoXEbIou+4U2EGkrNJ5FLF50WzZmhLVrEgG00QofIC
D8TAmf+EZnnfnbifwIXp8EDDnZBv3Iwgw64dZg16zwefVBKdJHRsX2LiO71zfeeOWKmjmyvtA8p4
wFr1Q3XjfGXXCfkgi18f2gYEvrXibD3y0VsRJMNIMZwPWUG2Kw0kFkOYfSi4XTrJQBSp1NnGD0j0
LhBECY9eK2EQiptK12e1AujFFSojEJFzMteJQUqzTufh/+h4giv4xOg3kiT9KPBcMGeGwWVzbhRr
F+k2CTuELJDgO539Ky1BSvtpDaZflFv6wQsDIp2WmJque681DCigHdRREQpO4uPWX6r7/UEM/1Yk
dCAel913xgQDYKXit6F1L/Fi6mc8CJfkRT5r4CIlENGCn5g53/BBDTxkZiMGZWRmpHblcR9UC5FO
3EfqmDXSrf6P+f5hhMhJOZLU/l4u1yQ/jG0zZxUNz0C7ZGBhs2Ztd2zFjrbxNzN+Vr9PqsS43YOY
fbKjokAJlRsjYxZv1xlhI9MKtZAvByrel9fn9rqsb6GUcHrgEfWLbSLctnOt25bpQN5HWlMK1sMJ
jpd602foMND3XFFbvFHb5cTtseKii0O6M6BZvdrAm1RPk07BI+50hF/fcTekKGGsYPcQ4QxY8Y7b
KQpeq9qUtp7reDe9DThU6hSOikw351JeZ8kA+8Ph1/GDigMqVPrhhB0KXQcx/ZVMVLDEkA5zxLAf
W1O3lbzXFprVEzgeawnDNfTh09zeJBEoWwr5MPHtxxdFp+PxJJtzPVp50nuQ3mElVVDVTydN0KC3
scZFoiyszF6+p5e52msImq2l6eSdh+GU5zbhW62g/WFg5ZKbwqNCk2X18zFzicq/sLwQYPfYQmAw
rhZA2sTWGXE1ht6OVTNXuxWeHZs+OVA8b0MkH31FwHvkCKz+Rn5XlhJDiluAUZsrQR7RK50Cx4N3
UZudTiBaBbHiT4jafxLufW2aZCBg5hbbz6pVj6ebi5sx1gLMnnBwWA/98B0dv3b2f/tOVXZN8Or3
kG8+nqwm2qdqSaLSUkQ0g2fy0ywDww1eotQQHC7xO8+rTDfNEVektULA3aybCyjqHufLDSa4ntlJ
F6Uh35cvRG7EMGxIGpBNRTSPP4i4kMpcg2ti4OQk8gatw+IMmUCcGTHQ+XYJf0S0ZZpfs5ig6cPv
Pl0gh+kS7wayPc5grO3ORol73gwcLbiC6wP7FFSm6pN4PJ2uQgK8YLni89MhEcOsXjcABCwWyG4y
FiaJDGbFmRTWd1Vnp6iooQAfif+ndnPUlNh1FhIzccNliguUs4xDPKT+zLuvti4eifwTIcQmSIyN
3AVFuoyN+E5ZH8khcAAB9W7ubCZHj7a00ZiNxfJe3uQyUaog6b3IomJPT/u8pspsbdRYRauItt6N
USxfghNpMSZ0WmQz6No6pdMY+g3RL8RE1RuuVaeGjh2HUiinahLtxnQhGZ2Un0uExrDtMKozCLlj
VQZUnT8J1+L46Xt7sykaqg/Pw3ghJUJ/7mU5Rk34evtOp7wAKr4w/wqIs2Z/OYZDUoZK9gZgpx78
m7nk6gglHroNs+3+Q8AvvM8/yr/NUtdXJqwvXFWgwnZZ8PJMS9mwv2/S0CwvoB1G4FQVKReWR+5j
7LS+kD3CNlsz41Ng9SlRq7Qw+RXWECaybbPXEDSymMCCeBO8dojmLRwPyqYuS6IhSp57YoWWVV9f
wOJR43YRQvJ26k40OEIyQ6374UWGYX6d7aQ19fZyBALbKwC25UQfMkgqhy7UjeaiYm2XvAm8JlT0
toZmvqLh0sY1t/fki9K5UIrAu2xCBtZv36lnZyqOptaPT3vWJP33U+k/xaDSEmWC5wjEP9sTcX9a
3a6Fa5xEDhTtBQtA5OnclIiuw7vK++1VvnB/JNYfERLUsj1K/i0pcN1J2vq7ML679zClBzVK6Nrx
+HhPEupEBW1WOOS4YFvqONXx84zhkLYmoeDkflZNVFeY0D1XtPWNRV0sUwayLhuAg6yTZdDDVY0t
e6kxwWEgLfQBPAvsesyLR9qiHy5vIl+9wVKgDqPgizjuWCLGhVGa5gdAv1MEtGhzn+zJmavxu010
+AVCo5hCFLNgS+ZJWBQA+bV8GqA4Qc0+qk+AglWIsEhtZssEljtY+Q+W/EB99ofUMGMzmRjJEhj6
kGn/ztLqMxRefARHs5zRdO4TArV9CjTffipWikhX3wY3qikmQa04Do48BYy6aMBd/XgZLhDJW8sm
BoZW5S7hn7ZbpOcPIQI6NucnP8Y+LppM46JVQ8zZZ7kLaIgNIpGD7GGuFZegUOwqSzkFv/eKyIqL
KmRauPAY3troZ0Kh5vYMUFsp1QkoIsj7IK5eBTp7VFghoIEKPaw6esAaGnT/alt3X8q3QCShhAlE
R18l4aWZ4u6IrQekVrkbmUJu1hdDr9SKvUhBvhkB53yjnm/yVZ2zAHebCF9LFRnpxb3C0xBP4jNs
T0X7JLWiSB/4xvTl3eAMLtT8MmEi0if6UYk5liiU2yXhjPEEMdrJyKzZNptz0+xv//PpfuUq2eMK
i7Lg9mMcwCi1Ofo13w64JbTLVPFb2uTJQ3/zw7VeKjyqDSiZAYb91afCT45Ykab6zuHMLDjTEMdV
+LQIAD6TIIxgB+LyV4Zu8og3n1yNQ9BkPmz3yVmGNaSpSjYZoLcTuLypA6+XP7Sfg+G+qJN2Bdwa
YWvwPViKkDBFJbaumIA79AkWcdfgVGuns41kSCbVhdItRv6N3aWtQv0/9HdIaTDbQrCYDC67GPMd
FNts1sAKCcMxd7BU8snLBaM7uP4gULMERXQBBTVKTBkvKu47VhtvdBOoQ0rxRSWHkSKTEHe8tUga
Nor5kTLo/R7PawsqNkWSauNzCKyEB/EzqYKUGcefD5tuakxtkcBMIn7q3a/NYaF9YVO2mlIvmK5k
P6RKPzUJNmScxxep8qTyMeYQ/N9QTELKCt1cBXBmIJny7OtUExGZOK2NbqMaopRkYTS9yoGSq8ro
XHOUy5kEWKTd/f4XBtT/LhEkd7YyvjCiCYsbGr6WP/16aN+QLmbrF9G8oipynn1+lGS2EnJhaAFP
nj+sZiO5MDa1QIltl2yXKuuO2Im0AuKowrORXtUwUqeEQkhCU6l2dogYojNHFr/fvONeabLGuMWj
6LdI1/uZodxH2ufMMv57Gazss2zqm8g2h1mWGKMYpQNCl3Zv8ZUkQMhOrGpXvJlG+wwzHmFxnY+h
PZffYD0BhiAFW7idLFLonG4SrGgMXV/MFP+vOfODJ/ENIBHPL031zuvt6bZpAgu7XdI/L+wTW/MF
bAhlPWfYtk3yJgWOkeQ17HZac4Nh7+c7zSnoBGuEG7LCxCESPV6YUTCjYxdDr4Myxu/4pDot1RxD
wUZFuD//HiW6dGhBneQ6+St2lWOIwqgiFRUA5+On6IG+COLtCjle3I+Ppo33+BvL4177xkEWoSI3
aKszDYaDvO47QLly1+e1wF3WAacD8DJM/UDwVS4/6c8FbD6d46bgJKjfl0iaHIEnORFMWzndnHIO
GtixZLtabgrjiS8VhCyyt4AWEuYR2NWVegQRnfoQmkBip/nFxdNUlLn6/ylR43iJQqgMJSnh3m3m
26i7UVWzezoBJRiHWx1DtB7EAOQPJv2ljRHKuNGZocqVBCg5R5SXFBMVk0WRHw8yknJmVErsDvRm
MrmnIndTCTwBhVgcKdCHJJZpXg6ci4ZM7/+3cr/lTZNPhfwUq2uC4SPFPxOZXDqQ+tBIbTd0gZkp
qDfliv/hhB9oGM72n0mfB5vmnYXMDyB9b3coGiFAzM888X5wf2FfKtZ/X+wjrHPrX8MU+dC46iMu
093XOQTgPI65zxUxcxRcXvw93LVZPY+VDgRnXXY36O7NFPrly8n4tjRsJ5nCMRYtoW4kyAAD5bua
Xe3B5vmM/rosgQe8hGuDreC4NpDs0ekelUMrgy/j85SbrpjDZYKFZxizDOvgigvC2kw0zuUCJ4Ts
0dFBrRyjnvQxYWeZrNc6UI3qozUZ1rbhAsFS5NOyG1xJxU5v7AReiB6SuwHLpR5pcMjyi7dFmHpP
+07BJq1u3vKQ8BloENuXpRjUsCa1ivNdboQjd2/6WLKBT+MwyBZVA8CBiM4ZpcSX+e1jMbALlfvS
oKTmhNkrvhAd7YaxlqimdRZPo0/N0bYpvAh89ChA7c4Obn4d81taM33V4K3AsTz1ZOExKhSlZhFe
BXM6rrGh2K9Sxs7rps713553NnVuvkeTqQo6n9VxttvkGBsowfTBrwLDRA5slWw1ifVyIQcLvemr
5XBeBhj/Hy/+78YUUN25xFJDfMYt0i9K818chcAhpNVpabGz+Ss2x4XSs/4UVvaNjp7FDX2sbc7I
6X0sptCV99z2S/gaR1BsU/7RZgJ+PNRyZJKbqITaOV79y4QDF9Sa0eFOqMLpm6mZIb4DxmNkrTFx
ilF4spksdLKbw0QgSUNABowb6+tNipWnkUafaGx0DubUUrxbRmRWPkq5GPTJGv1I8/bpyhFNx2Pi
K6LDkFPSr/DevCVa6qI8GGiKj7M8SUiMUPMw5FzI3NaZzS8h42lZ7D8V7ROWDvSJEjNLEBKuJX3M
UBD6iR1OwWDPVZBu8MLT0oiXom5wPFOCMW1qkvFzFcdt4Bm9C9+RP2CVqtLn5mkV03zmvVCFLmW6
KSaK4WC4NvUlK0S4yBgIgvjHoS5XHJWYmZhU8tnyoc0iftgK6qsnwgDDhP4h9bxsmjIp8OiPeiRV
Kprx+B2mkeSmFKM1uW7WZU3elvdy4SMgCzOgnyFrEQLP/R9dGEoLQSmQKYyyTDwpCC/iw0z6Gjbm
gHK082jr3jYuSoD/3AlHJxYdMf1b2BfZ/l0JbdIrrnyXZTjBBy87RGhmqp4Zl9U3glo+OS+Hc2yo
QkLIQRfdAl1dPZTOIBtgQuqgJ3hQROCylKfuIRy5UknXekVV/4OdbxcQdTStxgSY0PK8XV2VNUaf
3nuBoHedSyCK1euwgCPDYQiOZ+MrBq6myGYVS+Pg0TcNdfdonE5Ocb8UT428kEU0CmDns9BlowqM
0/cqKhW7tFXQG75EZZ5WOxosx3LIuUYEp8ad46NJXQvNvDRs32Cl3K8oN2mCUxzw8PJV3bY5yJ0Z
alZwHG09dj+cWMu2luKCh6MNzxev5vG3ejNqQHkZXhIH48ovCIhIQ/BN7wJe6sH2hpPsYjSe3C+3
ZfzmQnSLFp0yepxENl1X1ot2urM8YUJIMTGpvBwBDAVJQ1wN4c1WMWYMmWU9ws7TpcQi5bZqE13o
zlxzX1JiKhgYd6oMZy5Gs2gvB3ysVyEp+bFNOpC9bUt6Ucf9PMF9oxXzCKIP0F0Zz4FEUdllzcqK
WdqKz2N0tsBAKJTZ4/VGhTDZQsqoIF/J8cRyGWzMECsf3k2yZw598RUcJzFB3n+cumZgpSwvYgKp
IVK1Upve3hy0fAcoxx3HY5vIM4gJ5T723/fsYffLzG5WWK91OYWY0qzf6xaJ7ZtggxjL06D3jrZd
ekTVdfyKKc7OrIaxNRt+syfBQFgTtqS8Jvk20/rX1EtV7/ikynGklwMsSpJ+GXp2g13B9lJ/bBY1
OlQZNShsfYX4Xt2ETELcKgrUP/h36pDQAz4mSX5cpBDoF5EdJz8c3E75n1N9QORfGFXjTrVxgAXS
ZtXtw10inaqa3dIZx8Bjk7TQjlFvfEDf6kd209bVVTpwH6ndeSrtngzGVGjg7kH7Sa9N7MZGTaqu
HiTHxoPHbwKiqui/KOcbjLbnsyP6skWrYg4bT1kh9j+yfflTdQQkfNbCpZ9Eb3KRrr4XFjUtLO4t
TZhnhCwrShNq8AIaM1u3opfG1poLQ8hvapDX3WI3t07IiCv9YZOXLRnmu/9yqEApdKV3QKE3+r6S
RRuZRLD6pgGdLzxdx339WRY8vI0ykS5T99eK1vQaekaL3Jva8g+pTMCcLvAUoIM6n0lImQVbY06g
Y2z1WUWmw/y00UVBU8T6UZfjE3uknSU2pD8bxtRMwmW3FQ6dVZnMQhnVkknsdnvImSqQTlhFPxt4
3GAUfL4atplOaXMyhrOS2fw1MuYRcAqSznZnxrbN+jt5G4RA9YTv4xFIR0vRG+Dhlm0nKRJUi2X2
GJQxHAOPJkZ2UEe6k4Nj6snETFhbRUo95f6kjRJf40SipCx/fEVkx8MZOGAWoXHBndU9zVCMey1N
W6oOeB8N4T61dPAgU8YhbDdZxkEew9uCeHdaNacbm3otb8fFvMIGWzWx6qtNcLa1v/uVYLWASC1v
y+HXgXArJdT0Rcb/mMTba8w5oqnEYYBhc+aTmllNjIaDnDdlv5+dZOZ6nTKIDOXexQNIaq7NalCw
7p59xM7gyA25pa7+dAEEpBcOFsuBsh0U+9w1TH0HgORvIorBje6vYszL92hrxpNyCUFao1gnJQQN
cnNq6F0mGgZpzRbmRDRuzA2rsh6xeTW4joHgLXiBlMGBD+cciLYmXWD9ZzBeScJITsgdLEJ79zIC
hAG2fdXiXpQHHIJTskwxqOxLEf0Ua+QEiHU57p/kVKbOD6FMhcR1Y078ldih0AUbrLQ3O059V48w
bWurEIStD/gHTmhaMRxEPC2Mh2SpsoPCl3SHIu+5no9hlti8aWwESOwQOvmmnRDKM6PClWoqG8hq
noy0OGX40W3S8AranKxD6Z4WGUB79AEGRsB0P4gW4Mv/k0WRUYV2H5SiN6bqaeJWCNndqxj0XIqi
cqqzNQ4bPh6lyQAqoWTU3WGvnErug8oktSNVVIjO/zTjhEz547QcTmMGpnhWz76dSMZnzvYPEa6F
cMW/xVb/5ALB4BfJpSfbnf9XoouB+3sCr59wxRUDIZpUqN3bDq1QG2bQyY2BNmco1RHdrCpxaY8I
tKSggWnLw7bQX39HOkyZa57pZE1EoS1W+7QL1yZkPOuh7OS1JoEBhk7W0AEliB4kg7Q7CGid//7n
yRkuV/NMe+pQO9KKkjFhU+Vy/KEqY+IpotKCbfWJdromjm7CA0EU9FoMJYSr6wbY1c+NBvBTmhP4
Hij93w6++MCEK4tNOP0G5SLOqbRPWxS7Yw+w2paFW6VrE0F/BfMzBovA6lM4VkBkqcyp2qIKX0u2
Revm1DT8mbGIWFelvqBqcki0+moag6PawVHqeAp8BlpJ9EDzTUYowGUKPtqdNclM44x8R8vPvgx1
khYTpB3hruNL0SZRCA49u/57FHGr53T7xmeSVY4vGH/6vI46AQsOwhnXQLY856FHjT3wXYvgcB+r
dE0Ol06sWTw1E9FbZO+h+IHWB8HojyRcEko4NleZu9NqmmGA/yykQZu1nKqBueEAtZ/z5bqDz3EQ
lPVZ//UA79pF2MhIFp8cWp1c36zr6pCYX5IK1NbhdIgQH446ZBDejM0LryMJuS0LN9aaQMCEVSbx
UCI9A8CfsNm5lB392RtnoSdeC0XuqCOYE3ejVr6LdmS5kRNNBj/0qU+e9vIf7IXb39Lwz73q+WFT
LkcuSC5TfPrC2IrWGKZ9U0xQKuy/8TcrOTYbD821Mrp9Pi5zOGI5hVYLe8v/4ng7xAJ6zXKh7QAz
Zaksr5VjUf0nL/Uru9dNkxZXLgn+2USlc/aQh8uvT6JSolnUlyGzvgWVwWIkZuvnyd0oXZzXdckd
FrRoVnEbo4wjKtpSrBV8eQfqD7UB+GG6luZezdI3VdbESYhQTFfjCqx30/g8NHv0p0ZbITsPIIOW
mQLOvjdciEazlzcCysNr4n3+9vXUMU1P+3yIDfE/hViXDU5vEjdQcr7zc7Gdq2gMxiG0k5unoVDh
38lZnIwvqYb+WMKyszA2ErN9S6cKA+3n7M+8h6AqM4FNSBR3Aruq/qpluICkMbb9YxLyJQKGGSB4
2NahdiCJgmGRk34ldVLk/COH2pvvL+LWzkVwLQ9li8D2FGuLF8XyEsqOumB2L3Exqahdfr1JhjCM
nhuOQIbXGkEKjsK0DoI3izw+DMfUzgFTBb/MZCKGKnhh3Tva9pps045tnFCy4r7AbUgIvsm566/D
tbfraJnMOGpUOydBJwAGcYtQubcxL4tP9JYwdwLE0nvPfCxY+q98IMrpOJg9RF35Q5HAvAExv5WB
HKT+Nu2duCTN3DAta+godcyHPmeB4PP4PbTM6z4Xf5YJivehRABxwGYStCi8PZUJJSYZAiu7UW8w
KTtK3rCInbI8R/eiwENA3I46ENa7hqWoQoqDoMHL8zBk9p5W0bZ+NHmvX7KSZrPnKiCYbHde+kwG
mFFL+a6+mEdrmwbr9Dz0mbhiJGpmWnrap7IDlEsh9dD+PVuW5KJ4Cdiyd0q2i415XF3qUDNzvIbB
wzKqeH00CjIr7PILFDWTx2wmo20tIVF/Cu8AxfE6ZNiXCb3BktiT/rD/Y0mJyljZcahyvb4zT0g7
0HKfasLC5dxyI+x2k8Xd2xT3YLT+xFn3OFu47rTeLZ2XW4OMNm16Y1xdpgy8KWh3E6PZup8JbTmr
TA7coy1fDAZ7nal1arM9PHHHGgQxpySmS067bH1dooyjV03GvvmT86rCPvGiUfDdDJPiH81GpM44
KuP58LqqTvsA+qWdmwf1GSn5Befj0tzw6MRyn3rA8i/WI68J5C4NG9nlLsmBZZx6BxT3+7PQ+Z9N
wioH8GHzEBuEO9+HdAB/gq5IodC6ezMS+C0xDk34zLPJxK08dmyFkoNlnR+UxfPQysYoobVO8Tun
smVKaVpQ8zYSSZXGgZtAKVXG1FUZ6HzLVQKptStsg8dgvM4vCXY69EumsAKZ3Nrqn3ABEut03VkZ
GoaYhJvBcoJEBnS/CLcoXZC/J0sULwoZ6opixS74CJF9aBcec1vm6a6zPtD31KaH035lIjR10n/c
LJPmenAZui7+Yb7iQh6n1he2vr1SczZkCDlkredHCD3+PpPvuHQg+9R+yC9jvjxQS/2IQxoKbaAB
D44gVY4bRzetI3SiXRId8qBFyCTk5GsadtoxN2Fp8IMbtneAniDMJcPupgtionBL5Y+Jif9e65mH
LmYgTbKyVymmVgH9MFt8MzneMJ0C8kF1Ysvx1yeWmnr9Dvexhe9NHhP1vMGVln0GwjjXieSzv0tY
+RplwO/5MYgr/PafmrJFFYOaf8Yol1Qvq1TdspU+Z7gv/un7uJtgfN6mwIBuP1HUs/K5s0IuGj9x
MbybQ6OEZ5iFnqr/Zbcvtjt/65DI/k4XSEkOFn3lCG3SzQ/ZxZYFJp0tSx+YYGf/wPXo3msm9SXA
1qVH3F4KSUGXmALRuA1wYGYe3xfBq1MEsMAHkGFKU7K0Fd4niSQZaVjBzSgIN28eGfTH/3HjB5ZU
CjoVcQVusx4gIphUqQN6rB8AT8g3m2u2H+XNoKso//1XQDHIOV9eQdJ6Wp1xGBYACWDoyfzZerTj
AEIMjq7P/pcFUxySCLuVIMWcjCP9P2fGe34dDLdmNvs2vfjzgMmuF7YMVgoywpRTqmpZ1PmlXwf5
aSX5SV4wqxgtSUJ2NkoG4m23w3dvLMZ1BkuRdC5CX65hxFlXDe+LsmtfQuNJZSDVHqzEz1Ep2bxy
THKRD56wBK2f4wQmiW4PGOIjq/xMAPhyAMShxnjhQD2wu1Jo5MRaA5b1MT/PkcIAwMgQIPssWabq
2992bTQCNT7Jsx/BGLaQQ4gHw89e4g28LxrzN9kcwHn5vyNhU+9gaTIb6651pzAyl0uYzQxoA9R0
T9wFwm/MEb6S30O8ZLNpvxMiN6SEH8CxmewGR6ZmwZlD7H56oP8m/z+4UdR/P2vf9+Qzq+jmS8oN
h+z+fs6Xhaz3ZdA2bHTSoZ8uRD0UP+KVH85sDDI3FliOxje8YC60EpBCGKJwWAfU+xe+gXLY0v4c
8l2UdilOeo0+sonLGyEviW8glBIIlLH6Aa+YSpl//f0cpJ/pvbwpiIevsb/HTZovA3ZsPOFzQkxo
XetcTLWHHxxTAmZcoF9NwLwWjC7gDfJNepgDZ2F9gx+2KCi9kbxfkkw0aOzbUvXCLJL0JJAPq66H
pdgajR9Mm4gBALtH7BzvbiXAmDARrxTlr3BYG4ojtteQlkpRhskaY7gjit/nQZ+M8mvl6HTq4TjZ
7Sd7utWB0jNBZesBSUMxpXKP4FpsBOxtuCHp3sLJj5DgwbK5+rZkG47T9Nq3upN5pd47SWjPjeC3
IM0PpMDEj9S2A22y6BSRVrMyGaPfg4MsTs/ojKCbRUQCZyEsYWekEv+RaCpXc2gW0aqQYLuzAogl
RE5mU+K3J2U2s3dSZ1i4Ki/YW/FYe0hdSIie6Xjl8Vj368dlJ3U6tRjuxNCjEOEvbCwuYmmULW4z
NH79zPUz/b+LN6qrPExMqmD5JT4BV+poVledHowyh+sJlqt0iwAEw2Fw2F4FoKJBd7mJLKkuhruD
BW/1eqcOL+l1wNQVflFzU30THW5GhgHmQLvH9dfiXYRDJ2hpsbGisbQFGhmtz3I8wW47cSsPkWi1
+RlkToLsKQ4Fls7DfUDVJ5ca9phW/pI8NQb1VPYTYScJVVHDlrcGDBV0ZOHUV9prQPKlcomQwgH4
T8N8FZu6QmFQeJr3p+b6N4jrorm6/ETZA1RN7O/jvb8c9xKX2JCRUN1vcU+S5smo33qYDhrJ2k4Z
X2PReyBCVaHXdQc0TsUFrU7WsuuIoaKPRIq+eQKaXlZ10tkzklRKHqVvZ8kSFEX0DTvMkVED1d0H
zTp5eHbO+Lxd1n4OH5nvHFdGynRJdI5iCTxNn13MX4mPcsxQWAifgbTpeDea8vXvl4zJ0p7CnIHK
mujbs+nmQSQZr/FMpwdP86icETFuspNFVQSg8OswEY3UNjo16ylW9WGsd4E5pha3NwmUmTejHSZu
yZOdjjjD6xEYKkY2vG75AXJD25BSD+s2nCFmLHPYWAmEHV31ELrD1cMZT4Klrd0HFHZp8glbNGTY
oIDqdjc9E2WFXSj9cp94/voXmbkuRKE6xUnyAup+OIIRBsOab9JHw8y1AoX7Qo8nZRGMjI1oCa1F
0ffcWc9+ffCFlzzau1LgJXjzDTWpxtteszvZ2z8ogvuheJKy6wVLGU6MCXYmL5uPAcbe1afGqZ37
elbMyKQBQe2EPXFBM6niYtXRCqQBVHPjx81hS6a911lZmlukjH5neOBeft6ABdOdmhIaOl0Aprg5
L0tDWRnyYgTlI/2vh6X4A7R8OyS2Oi2RB+n1hnBSd4UtWP55tLTeqAhkJo03O3iIoA0yZWoNYhNt
G9DyT242rwQaYy+jxh75HEu1iwxjvZjq3jAwVlozjcJydLxmxmWqDzwmGn7gVmJsrG6QEAHX8GHm
IXYlmgxvefahprrUmiwfFakhR6GE896tDvPVcE5gFgZ5+eqEJMO3M/VSyMZOw0QUKPgcVVfBVWqC
tz08a6/Em20C1qIUQ9KPL1oLEEgPW7QNtfi3fMu192O+huxrlvGQykp50FOvH7e4PsD04Zsbo03R
33gfxZX4DO+WncBpo+zHUW8mKSwxWOJGbxn4IOh/Haq3ic1AlwmKACwRvU74yem7pn/Qt3PLEkAp
zQIKpCRxsPGDAH1OF/SiGa7jvQgKyV54SipOOk7vM/wwzbUdXD01lKeA0Qkf0x3+ih+t1ehoG2nU
1+uJpg9Qb58F/kf4vUHnuSFu9pcH/1bzbPgmnA0AzxR9jd6CWgSiK0gDbletpXtKbLxuczNAsFSb
uqtjzgdtUixJN8fQRokCJ/fX0ZrUOaKpb2/Bkt7ioqaXuN5j8/U6QcPZRp4knAZP8NXj8NSt1KjN
AkW4mHZdZ5LLcart1wh+/HWHxa+aaZ/oXz6utZUNbgRbt9ypWcryYAmUFpyUnIaWa60r3U9ADrYg
XnvGInnBQsI2Z3zyuhkP43CtBDDz1xfHKF1PMcx6FQptN0hB2QS39sC4z3Rnmer1sZMwPjRwZqUU
OoCRDerRTKctnuE46w9Z7d0b+bE9kR3sjh+hLa0TOb4ukm/XUveS5NJKnTuIa4mAHtnUQXOFpwwk
/HjkF+QuLsoLoaV4ne+ak0bO6TK8OvbAE7hREZDkv90caoyh4AIrzY617kCScpJOOD6NoKYCPLun
I0g2l04stUpKGGlv/jqn0YqPwmt9b1DTMqLgHB9AW2YKYqHQsHAQqOaAZ7lAva+Z/HO2UooFf9F5
PUojrmIhYTfM/OteN7nGMnl/pU05hUrpi0PhxRzrcotrSsEj2C8A4CYTz9+8e5GuStOZOM2KiZan
sxcx0SLwyaKVXBLk6j+KRFgEoOuBwbxMntDHGi5hcwqR+wwgErOWSc9bx/c2X7GpiNJlnrPPDsio
AGIf04eTUidRe6ZUUGtsdeJc2c5q8j40rE0USzqE+xNcDUjYAUP/tkK9qwlrlmZ/9/QnfXFVUFS4
oyUGYg6jyw7xImd2AM4dTVKHegQChKoKN9tVTq8eSmRNstH7cS9Ls9hPq9Jc+smgqi+RegON7Rij
r1ykjP2Xr2KBWoBftL9lUPQlRufvhJltqMExDA6YHf9rDtkvP2EB25UX/LjrbKrVAoHogGUttcsE
7q0Y1DTc3geDUfWNqYBcJ4jwvcRf/RZcAyDmVl8NUMAhevZEgsu2JkcFc9a1VmfhYe8YOqxxHqgM
0MGghsloW/4KEZi7ftooxZYJGpLxQskV99vvDUFgGtDgP229KgUGfZ4QYDQoNaP74bmPL511q92J
c/4keWPq7sdbeLFHeUOQbnNbBL4ZpDak178bWxIop0aBArMxkf2bCyZqCH2SsBY7bB+0jTWtbAm4
W0yP6BvUTHDLFQuY0iO3TtWBO6nmfZoITR/54OitukNPxXbPpebZPwH4/TWk6t8w96TKMGzwrZ3h
7CrzciXGnLhkA6TeQU6ift48H/4DQKCr2Vau0XeGxjhTi+6iVzmnDiXXe2E21P7FQCzLHTuDZSEH
6Xge5EDCzJ8DvEinu977CSLWpUlMyvv3e6FQIHftHzsFwRt2oSry+6fYHYH15RG760mmEyP2uQWZ
kGWUxf7qfHiuENui8VuK/GaMZjXO38iUYUrDHIauNXA2fQoI3v9+itchD7vvnyLPuYmHnNLZsEzk
2xrbK+nnj1jcWlaxJJNkICTzoxmN4bQLS6ZEElRD4cPdgVWJHzA5O1Zz3EY3o1onrER4/V941D4o
budVP3eYQmXe5MmcE9NpP3LtIwEWRCnzRJpcsT26w5zlisyjn6Kamepd0Pjf0p7/Cqg95VFANp7W
Moo+9X4kB8DoQsxIVLW8pU1AYZVrvm5MU6ngnqQ5X3g/l2mnmZ3t7Vr1YHRSEJb9MGNZk5A9+mrf
CWG+3rFzuUnl9oe4eUACo43ME7QxUvHa0ooYzvWSuURbG3OpntcB20hBvbUGOuwtBcm+wo4ROtH4
hp/12VKJ6voXJ0EQ/k+Fgv6EB7xChYB5HW2b4gUbT1Tu2uVhttq6rm01AxJo5Wrz/XWO4jcut+RT
CqhNiJeZ+aofO1nUQ862YBS8jmjkXngee791/rrYBfQl8CyzJtknxwxyyPdU3+5wwPSeseZS7Rb9
lDlkkdQV/ArHcoWLGhl/0d6Q+6SP6jvcGPqwQNDJXPWxfhcqV9LoFmub+wYMvz1ZChFz8uxzlynB
iAxY2FYZvmmnYKYiNJwspOFbStx6JwTIEI9YDZbRV3awPNiBo7ld1xrcOnHm5g9pCoU+xYXXIUQ8
4IZjqSvHbMvHqLeK9qAHsncquuEE+5Mj7GqNYM73vjTFh6lmY4K605iMLhmuAeLBHWZCJO84W4ug
vbpfGnf0gP/QYykYjhxK5jiCyxyKObvZBmo85F57fekdLnK5TUr2lesO37rLfzHzvGmieYQBkSQy
R4ohnlZApfQz4HapvyLwjMXZezKu0FxFA2NKBp9jdgRA+gVWiVXNczlzHYnMVeajrXFa5wE45B9p
+0DZgQxy4O84K/fyvMqqyN2x4nlB09wzSxKZIcAOR8J1e/vcs/zxyyOVkCJNDWN3tnrbLisJ6DQ7
lmbqgd2YCeDPLAh1otkdhZvPZlYRuf9aM6ermNcgiyOuIKypS0Y4oIYyhSUqCE8tbB4g+FNFWEzg
ZpFuw5/jP2YR/kUWWtoo7Ow56tTy4qbSTsqLM3tGmAy84CKqxWuxQHlhky3bFEQVJ2wZ3X2SQWt6
p455HPICyKDCbue0Hdp2sEyIWoHsgIl0zErhvViW9az3JF4xKNdntJI3cBREeuwrcyUsHAeFxZHe
pXxEBXqV1ttLzVs0RtLS5HwmIr6OMF+5YzExFSTYyds6pAMc/Id0gc/iYIKTOeUndVUW8pJHFGH4
fO5qTt7bcWg81aQHM6lkwbHsri/+OZpBszGaS1SI+BE/FGiwTJcxWue/IqPdMhZRgaCxmvxUKoMT
LaxmU1kfXXmPnaUxC/LazObLZXJo/pTRHJhSOKY/pqE2OJtKMgiDMe0CNnNnffGio9Kh7nOp0KUn
h5jZuWamrUfVHI2GVI7sK3Y7mkjHRo4mfQriB+wioDanEycIblp8LAEuAIDp8gvA0/CkVoJaWWK4
Seght5txjNyyFGREPR92Q1raliPwHH5WL55e1aZQLh8bTR2DGyGAh+4ItTt9mhZIfcV8y6S3PKCT
ZazqDOWkv+G/p4kw6twOlv8UURSuL9BnA8+nV9zODero04T8iu8fERVISE6TkvXDESQxI9tbGtNZ
ZgTlvps6vjOk9tNsckuQ4s3Pt9pI0xAfbhq22JGcXq7F12Yplc8fgHmGM4KJcFabQSL9Y5mm/RnT
Je70O/vobNKve7C/Ul2PQLlSMQUUM0LZTHV/SbJ7nTKEuryUg8V1kFFf4t0tmJ8x2+ziGPEld5Vb
0aGtotQ/upBfwpfeLM5aJM9YZ5FgnGHhcQZSPFUrH37Ig9D/RHJgLQmcFfaHPz8Eg66RVdBmwBuo
dpy1EWlofcGgmQkAz3zWus6b9Wfb+yfvdBmqhaYgVsvJKmvxGglJ2YuN0QtLUQiAdXTxgFyYxfdk
pEhK5LA6LmuV0ZsHD6K6TCP+tndk/iTMAeNGdDRqp0R7KGeyjBAmqfcJHyWI9hMdJNA9OtJsJah7
IfasxQT17S2sxLINQF6ip/v4LVcbOgycwfJYB/4ILp0nQ/byMp/sGY2JOVzwAiwH5iQ32HJnBJlx
fuyuqwCW44+6HBeLOcy8xBPq3JQO3QThi4Et9XmDCVovpJCXnrQ1+NYJRtu9KRC7DyrEzfv2BDTF
1GqqCp6LQIW7nyKiOd5vrTFhpz7ov37kw0B8H8TNNy5vR9B/CXcePrBFJpFi8JghCo/ZLqnraMM9
iUAqxeQI74piHgWhHiIo+b3Ib5QEzauVcAYc/uahUuvnWrdOoz5WMih8PnXPqe0I5ARWgsgyL0TI
QIWDz3bT9n5I54F9TvnbTeAnmsJA7rPz1XiHaFczmH849hw+arhufHhH69HS0S0d+RbpukSz4gQT
2uaisey1Itxe+dL/PQzV+DXtAOUD6JOn7iheFeyPqxNRA5xW5Y+7+UGarMWnFce1UQdu6byXP3cq
6Y4/jhtx2sw6b7CO1LPUm7PEWnpsdynKrTz/DVNXUV/6k618I+P4BSvRK5HxhUdDlWdxsWiHiYJq
YZCnySwTTZcMhdcnbqTv1al6XKFTeqcgPe/bJpART4JqL+o8YWTM/oNSpvxcD/Ta26udkbO1g0ya
mP8olQqEhp1mIqK02vcJxMqwHbfSato4zCldwWQnnqIGyxnSd5sDN0uYMWkKJAu2AcpIi+1d1sgs
oOjBFtc7uiviGMEuQGDuKIOQ32hoJpr9cn/H14ApKqJ5Llz8muttLgUMvAzXKoStUOM3xdDUBTj3
CdFTwLMpbPcc9NmPxY9C4uq+QCNL2Rr7AZxJynnm7pr94mcWozakvoAXzzrYsdxF4VEkLIIcWhnB
Tj7j4YNWbHZdNMw19QxXCTbMVCFhlJ5jM/nwuiTMD0zuWhieKNNkgVPvq5JfSJAJIYoT1AUGhmFS
HExDay+bYh2P4U3BQ8rWH3Z+z6XSvNyg3vFqPH+/TP+pcc/a7BSt/CW2Zgm3JMVRKUcOhQE86Acu
FV9Djx1R6EYwj30N72pozajImIVmCElKlRbEGnTDxviQUXhEYt32vOkeU7mlWBkZV31oGPdExJIO
B/Evswcg/KJACX7nhYvBL8LdiWeuNBnI65Yjrb0pcTdfkVQNCe49cGI3xBRS7ttAanIRc5F6Ab8d
DAAwQwahnv0belujMC/Q/vzjHzbj+NCvMn0cqHhW2VNK3cKP/jSx6l4IZXaSjcQL47tNwn/c/N6p
ILWs5rCPHZOAdWtatbgQm5Zrv4oMvMrmVddA4D8ZyXX4EmtlHkO7SXVBAgSnNXmkDbnHz4DShwNa
47B1Q4Ern4cl8mozxPxbykHh2kyzr9cPPpJZiPiINalJw457qo0QCZfjUZSZzpTBfDVIS0Arruzh
3QUszYfzsMprfuDkk91Dqd+7i3axJcX5rcYAcynAiqDMO3EOUEjpZv9on/qEUHnzI3GIvLa+JhoD
ECCHm9qGg4gf+wbVQkRF2dlf5MweOG9Z0o1li6VB8DIeusEC6Fqid2Jq4gdH7JgHGDr6qUw5CZqo
axjg9ENz7OSg1UM8OT7cCaUYnS3RY9j6igLn5LsTNYTZ5KvAYYiIPIqAe/VwBQ2w6jie+BCKUJB1
cX4Yy/fUGxHl2+ILG9fRqRUIuTjaHoayaxItygFcN/SuewC1TlAqD3HHlzijIctKbs0gqc+QrwTV
poHyi3p4tRUT072clYljctXN2ye0g6r/gNV/v6jDdU8CK9OJfKmOSMD9TsPZabPLOczQWGxZmhHo
KMkeGEuwEScrgHWCqtBZ12Ht6YSoGE5ttZX61L+dWkiMOOZ3Mue28uNH+N0uiATub6sXXfFNCrS/
JCduSsHgVHNTm1pd2CpevALfgeXIpI6ooMysZ8l7BreijyCWlynXSqF98QSE7QCaIus2zgfh/TJU
KPLhhCt5JuFxkPENeDfD6p38NG4La0xQfhaKjiF0UpzlRY4SFMtsWAvgrqttmdYOyOW+bWvZfC1G
y+0evI4UpsLeey9rXvaDJ2D9wEHxm1eu9XnZYxmqOSZrrotp2cMufNJnJqA8comvQH2g6AazNmR0
XJ+gb7EI7cd6tPPuIfyfpHk8EMLjCMV0v6rb2yZhSmU059C4S7VMGvG6WWpQ4pXKp6iBV9lz/wRm
M0pcdYFuGkhOZ4MIyU5jLvJo/z9nxxyec0U0UXsUckUjGBAoaRzLYKzVnJjfTyUWpzDSHokqSICa
FKq9hX+f6SN96X+gRSdeSaJdzkuC3w5n8C/6kFVGZTByU7LRTsehXAJaa/JwqfG0atbH3zpxKU8s
mjlFFVd3lO0zxNTE8MNm2h8KFZEpry+oLhSluGIe4ymyW+4wySzqq33UXYytjpnLXzbYnhXtX7qE
qvfLfXyOt6OxLmuDPM7xtqCQXkyEDEcPENddZsTxrQoPf3iqvENcwgg/wRE6f46t2PY7U2qeivgX
nPcAhkHzTNFfx//HdUzNw3g287wRwqUMFbT3pQ/I+8ZDb3o5+Bb79bS+3wJrXnvGeAYwj0rmmcEY
UNmH3CM+BaxFoQWUhGNFQdasmXQehF2zHOWm4OWKp0pxXIFdFzWpDKuHHtiTYBo2bz90g+ovLOdl
PN8DEK7SPG8agR86/QpAqMb3r9G3Nr96t5UhsX7NhJsF95ACJesuxPafpuec7Z6KpnCzMjlV01rd
nvltuurz7bCQ1Op/epCEMYIwPphI9OPvNfwbg3blU/I55jzSlCw1pY7iKsY7BWFPXgRJCrKkI92x
8wqReel0L0k76bFlC0qLq1u1ruF/oTIvJDfgKN1UJNLfrDCp3EmsfRLagHpu70vxrJMMuOjoik8t
Qh5h5q/AyEVj+UPPEOnFCKnoDWZPd/6pUNKv6XCnPpNJlEQg0kn2ihQg54qfppiVQF3lsoh33rZ6
0xEKoxrKG5TokI/vf4XETxI5+sNJJ/mwYoHQe1Fzy02OrzDzSUUPDqgANiVl7/v83Ol2UvVJckEs
xVIXuS/c5Do3C/nraf3PAJMW4M2td/yMNyOBdoQ+L5FcD/aapLxS9FqyrqSOBxDNJFAJeuWhMF0A
JllYMzQvlA3VdjWuqFt59cp6NCac+S6yomZCRCgnnD4WYXJ+/yaixgYqrdbNlQW1lFcTezrFrzWx
8e5JMWN0p5nvUhFLzOTGx9koTX5umaMGAYHqzdSo3NbHX5+3g29QeN+Uj+VVoScxdnwFDTvLBJ9B
be3jtvkdYNXe+vGoa+twkkBlZD0NzYxkOytWCs4I6O1kRxPI/ILxL5M8hMoJQbahgY4Vd2L+y6vl
SK7uKN5YwMxhwompg89lfKf3s7wJMc14b/Xu60C2sVApMAv9a5evk1SzszXM1jy3xENrfywdKhuu
PhYBxiX78zRuZ/YKyNNONvplnwpl/4ylvKqMB+EFJ9ppg3wFAM6aSwL4HLRdVd1C0l3BPidaSmAJ
OnDTE9HbR6Wd1mbvLyyu3eWAQZD7GTX9c4Tj+K24D7OT8h1q2BK1Fie1hKO2FLtDVsVvrzZCtMaa
hgQB9Y9mCYWNKClHhSM+0wZFciKVNciht36RMYK/y9oedllvJXM77b+azHphVh3ib5IpCoD+Vykq
744bIfHZTx/pNirjq+eGeJihy0vJt3MEL/GNpxLgAsxR07P+++MLGME4fqtsuIH8CHKMPZi4mzge
t9zx+jbSdh8VlUsIyqDptqRvhiZLoNp+JlVjzrEwIbLp5S0pGU1j2rHkd+RdJS6DC9tXgAWvf9N/
jLJik5MJsi6aaDAIOkLe1DiXcJxFOoerlscNU221j4I34MAN+qOKKaJbCEFeqjwUKqDY0HpVkkxV
wwvI5fek5ACnKtH9pyuCSUGW6Z5oSuqgOoG3ior5Zj7mmXUC0vs62qVXhqJhkJi6dDGpJYz2J8ou
SrdJvnEDeon4dwbwZ9PChlM6enZaRXDR6TrdBd892EqoWEYuKjvyiniCNZzv6P3ipMHfSluGquhc
hNa2Tw1ot/mI/+YfN/a4akv4osQwhxCbugV3FgMLPt0aq71dTYhj/f/QP/wOqC+d/hDUFiezCpK+
AAJKafuak8T6si3JE9xXgu/ymaRWDzwig+DI5fNmr01S4cyeD062l2zwMPF3Qq9Cc/Hyx5y+BSN7
QTwu6kKNyvEMcjlIzDc9PdvTKGo0Bqrl4i7JZl1s+pc56a1B6oVHUSsUOQMyRJVSXPZprjn9G4ge
zdElNs9oOPISR3dZ5NXhFTg51daBrvMlC+3nEc6S++dvuLcb40s2UVV1V0BR+QfcRFt6V2SR8lRl
QC763JWSGU1VMUHwJ6BG5x10VxUBn+NlV33ZPT/3C5IpS/95piGHd7Xj5xPi2lxQnCfyGgVzgc96
3rrPR0Fe3I/nqIgY7nycdSSFSqNQM32Yal8aGRfaqAEOS/xjDpskQesHGrTxSpNJhw12n/xGKwLD
rDtpvfFsKwKRlKpSN6FJDpWtyQxd6mOoY6H+jLXlbASP8PhNciFZh6b/NZLTDTdK4c3OYXX5sniO
1ZIofOTcqBlse/xfxLrbQF0gvWWtPP+Kyi6eGXJtshspbBgRbfkDUpljOo2UuB3LN+m9KOq+rzxS
oSo0MbD21dmYEhyJVT/10tOjR3Uyu+Bf9CATm1U37iHTbNJ7IAUqnRopzD2eOY7mU37P20AbG78v
D4Fb6FJqPg0n4fPdxdhMWJajKa9ashF/9+hrwVsWGL1lLi5poUovLQoAbcbJeNPmDTNdLrXKZaPs
FV0CuU7NM8J7QNdQ4/4rfuQYpCGUvEII9dIf6ZSV4GPqmB6kBmuWeLPwT0Rf4D/N3/mlZ0FevNR5
/23HAjA0eT6sRGxe3p5TJm911tdwqiyWpC8PCb9ugb5m9ucKBLU5myJzBMSsAwpA/+WqwkQFWqyk
LT840cEh4vj6mxbF6Qe6TOquUXBv22VAZLGZSwXAxz5dFfNB9RyC4oSWQgTD1/UYUNVs2uTIxYzx
YqShzfaEHoJOdQyrUIe8u0y0Cl2944y7CUKHy3P4vxCeIPxnCz/WPmwubwtlnMW+mke+hQBoUh+D
ER21znwwUBJ6VwUzl3+WOVqBEo+G7HeG5Q4an+qQYQXjHiblABjtbikzkPrE8RitVWkfUJdhqsEc
go67hcnpJ+ICwPl4ewHNdk6w3TLIoWXB6K0byYvqN4Sf0yRHYixpVUTxY2qDixBZCUtsluRRhgB/
NzL9tO2eGrvFSdYmD/pXXHQ9VSvcoOHDjoQ3X4QFoiXBQxZMbGxRzjTfMYBC9bUGe417Nc75jOur
CbgW8c9lKGs92saFbtb1sW5I7hTF4MzhziqDG22vI9WvslbsdDZ/FBfHo26M71IHYlzSFsmzLpLN
dgdrkqeybYn6o2+TT4tdXL9kREafHjDKhEXGNOrGpuCLt3n13QTTOtbRGanMsS00krjBsH2hiSJx
ziRakoAESEe6wS73UgZDfjdxo4u4+3wm/N7bEjj6LXBmc220cEebZO1Tk+1BONHd6qxxjlXRU4P9
xc1N7Vm+UqYUxFbnHQsEcC2b7cQteT9jcoc5AiNczs+wXZp58cTACLvkkdcKlLQoPKbzv1rBUwJV
l0Axp/g+WnE/j2eSyZ/cl/3LBdvHg2TTzv6QLyOYAzExEXW3Vft5ZxcMikkbJb4r2lzu/TkSEby6
sHAIm4GF4gKXt8fT/UOt8U++8330Q+ZB1U9CJb07NxjOE8VzIIpahkTsXC0huRZPnwRnXYUvr9/r
EEUbRgIUc8oc6a3qIaKDqPQp2/MhibB9xF5VI2UFo1vPfeavjZDM3Z+H8Z9wZGYoUnJEmjhapzUd
rwWpURjSnVzjUqBOf7ALMRxCap+uP51noFuKhNTWZqXBoM71IDWt8yWDIBmp6FcAURNg2flAumGR
xolKJ2fOCu9EEANiAr32t/5j8FSQW+ZyfVVLp5v8JQ8zRjXZ8tlEwjJ3t3XuAgDMX50bUbPTxlAx
o2K3PaXJzjFwDoaEl1qSfV2sKvFOMZGorFbTnIIciXs11PqOpYloT9KA8BveVy1GOufZUL/ReaTR
TrmErJfNrNNclTMXagGwLXW0Nh5DBpR5oesJjpfWCup7vG/OKmuR4C/b4Qbou0FXrm2oqs6f0/9I
rX/3mldpK33BfYDGwCuAjoe/iSVo7uTA6KDSbL8oJc+02XlE5I+QhsOTQlkO2OUnnWRird94YV0M
2KaysTgP/wsxtgHdSCqWhOQ7p9gOQPkX+MsMRNogHVWcarSsaQTjWOEVcP2dazOw+UyreMQA65xE
MGsd1S64IqWxcwHTfKnfiZweeXiDGILUPlp1gP2o1vXv2YBQ4WQI9+SxZtz5nIrLYyMEfqCiyceY
QR2C/xoT/f/WCoIy9kFljelxgCk8412eXHYwU1RKSfmOjNJARpUvsYgEYBJmJSj57pkJ6mjhcXaD
9ZkFiUtkYTOWxlWotVUq9nZLcQH5Ix2AmHAPY6X08daEGlr73HtrX2Wxix5MPR+ZQsQOya+pzN5F
liw4IxbtrS0C8EEzMGgQUrqv3fi14kZblBfhav9nouhUgVXwP/iPBlwY5gySRRkAU5vj+Rt/Tf3P
kim4nMfovPMHzX/I5QS1Au9Sgl+nn5rtsFuUkt2S9NU6sNnMJHW94EuYADAw23NM10IF4wYVFkeE
Fqz0TLjk8FNsxfFIeGG9yNQ1R51OGdHinaESNCqsbQli4yOJO4ls82J8S2lSQ7ibrHwNNvsXfZbK
D28/OsZvw9g9BiuldcQxJ/i+XWQPPTU+IOKf0wH30PuZcTBVAlJZ57QfpuTbBXk5ZVQ1kEorC6Bt
G4XJTFGaBxbcBbkXt5CtX39GGVNsKm12PT6ID/5MleeXgqIW/Wz7hlZ/8qH1uHqlS22Vq+GpYcDq
aFDtihPjc7NTdfmIOHQaobmDw7vos8MlcydGIN8d3KpA1L2qpolIKvaaw6q6PzYk/VqzESTUxl0U
Uuu9JTQRWiZEfxavcIuERYHSVfgzYZic3fLZocaBNCVON+aD8bnFy+IUwYi1GrZsb+SmvYl1K+3k
gcanro72kwFrelxsz7AdMCECfMeKEtQneHyHJodq7Or9C8hBAw4S6Y4gdgtlpfVFT4271xbhPBlb
oYven1PvOAiW+yURH32LwEqWwtAet6QXTRT+1h5PSkt7/aDE5KI5MaC3ZB/ZKxTG1qaDirNv9bn5
yM/Dyr/zeIm/0wjduaqmpwm1uXu5DdODB+xYRzL+wVwJUbyBBxIlrsMMFvf5HnqeGVF7Px7HFsYZ
/qn3Z18aceW0R1SR4z85aKnoQKEIiuj7GQgDZjFtt4AVO2ZFPENpDj23MRE2wkabovWDIUYvW/xc
ZmtyL2/6NvfFXCQFxyqogHsbHq5K629eHq7pdS6oumPgY2PMg1lxOi9Hia75xFOtYDYX1sY8qlUo
TffCd9tLbCUPEpBh3lC/evo4S9hn5Meslx3N7oR1zGm0tU6riguDTV8YmCz9BAf//PvfMqQdRQUv
GafYUw3lsTCI9NjO3jbgcC2E6AcQAMsBIsJPx0/khMau0rEVeU65Qqfa9zID/es6VSTx2zkeq9DU
CKeO1Po8MEPk9o3utvDj9RqS1QcsS4KljqoBP0ACBMgBDVgPA5YiPAdA6Iw02kQClkNOpLl9SyGm
DLTQghn9yURKunexNeGWu7zPKABK0fzeDmd9nsvcytfWaJOC0sgntKrNgrQzZ+KcHJaev7qVjh4o
ea9GauJLXlCfKqoYOmyl8zoGRU2lvWXhvu2np4zwPzbpKfjHKfWwEg0qXMGE9AAKIozBGofXPTwM
jJ6Y9ChJRSRs6YQaDrAb39zNepcAyHBmegjd842t5SaqsPQcbGsmSVuYTPbBFSNLAWw6PRmispj2
S+ZhdMOFiioX3xyxxhXyKygZelAIn6gGD6Z/TTzc7A78RrnyX7wbOYxFNow3vTTuSR90pRiRTa1a
8MEYsX452GCzQXUTwV1Qu7x5qEJZXU1SjKYyelt6OLov9l2fhCv03KiM28gev/93a9+Oy7lpnH2e
q0YwOEIo5VE7KFRnfCzLxvi72fu0AP+NTpWYx1RJ3NIJjSkRjFTHDmrUspmUlySX78+WF8f0Orxu
nVFGSv7FBGAyuCRqy4aOUfzaLV++y22uBCSynKqUHPJflow1mlTLpnqrLzytpm2v17HybTuOZvru
1K8ggPNGaP7L84N7JJi8ydZQrlYrFugngvgM2jmNuxEZizV45t9Vl0y2Mqhz2lvZCEez5fRCrnzT
lkrnxCt25JFJy2uz2TcEGlQ0ErgFkzsRyFrqcNXeLhFbq89VDaqgJPSn5sysDzo127FhKzBfBa4l
3zfBa4GS4GxadN0DEKrp8Gha38T21kWI8z+Y9sN2WG5ITEi5yPoUyQDv8ufh5/gWVwtyyxP7byPr
A1rmJf3WuR6yHNFfQLDdImrIzgvd+uCdp1cl/sreJ/rDlxXfbaBwMfv8jeo/c6swviMI7hwVE6WA
py54PNjUqphoU/gMp/N85Hmavp/TPEhUCks6uXJ5Xn/IiduBz951Wem8KPJCEpkYacXs7dHsFV9Z
a0yw+Gw/OqvBfZjpsF731e9yVx3YLpb13ATex7KqiN4duSTxodS4l6AiU/A1L28f0nDmqdVah+E1
AofYKn792ZVj8H7hKKweKljvXb+R+h325P2rCz1162mU1okyQ0pKa5cJ5vfFgB5CfBXKS8RK5S+V
EhrPAwp3mw//x3wCr7AOV1fl9M2KK4BnFdceAVI+F6Gg4Ujo+GS78gJSf/LjM0Xz1wbcKFRG9DLj
KP9E0NVZu4YQsxBprIdjVAkkh0cI4Tk8a1JCEdTH36syJFfoeqE6IJl5ntsnuaO1ZxUd2RicJsXB
eTbYpJMlg/AmnaD9O96Lqmlf/qEbH2hKuGX0yzaqroekCRKY4JaZYB9sVjjTLDiQGNkUcjtAM+Xv
J1Mlh0Y2XmmUbrlgB8uMlkY9bSphBJcWPepQKgm5jktwg3xDSNxf3cCicKbY/1sRlrObIUYAxZ9I
PVa5jGp7VA029eNrrzUAv+BDsT1EtY/oWIuZpQE5kByXEOi7eubyZdFoFNMdqhnrqHXg9oKVK1xQ
RbU8b8++8jaz1lr6KwLF44bU0Y0wssLgo+Hr1L3EnF2voOlq5E7Ol17BKfW5sCF5e7icbeM+Iook
NS87IGFSkQJyoP7YGkbZ5X/wTvxy25NPddKId7aQMAVuoxxtPHSYQTCvGnx8iEVZxvorx5vhvy9L
6HI0o5JPsBFuV0SvWvhNDR1FzJfeB++sERV1SFullyim+dN+9+wtRPq4cbngIDGQD8ykUsMl+tLu
sh6A24OFeOHZXxkTdl27JpCf+Ws9wocvgiYdBkiVbQothszLHmS4xmwutL+oxSxu9jX5vxZBJZqY
5+l9GSCVFczGxlkdWzJANc65qKziwJGu9BqT+qe+chJunagbkOP5Bjwi+uh6tAtzk/e8g827F7K0
RF9MZzDJydirjX+QBZT13ZyT9vfVT4Vzt/pvrN9tRJJV/B8SjHdpV+ns0Wz6oocYp1puS7jCcYHd
2GgE95CE40+KptuPcjYvcCk1ZZhLJ8Z+Hj6zZmJTkeZ/gKI/MltE1mi07kbYiTF6p1EC+ELQXK+Q
DUnraa09/QAH+RUU5WzaTrneaDcsU/c9LkYNoUvH7VszgWfi4L0s48jz/edeT/muYwB7Wn8mLeam
vYTpStmtMTLqpKcj6892FSIQrrDPEhnZ1hqWl3CYJpxtPIuPZg8sxaZa71EUBEFINCNiuuET+77Y
kkM6Q3Js+H/PY+Fid7gp7rrht1GIfcGDS25iUaqgIHgi1EK3HErmp6wcV9gE48lDi5YAUPAOcFO6
jJktH5lHCliXHp68jNbvjEq8EbZnKlDUhBKg9a/4hA56oCEhrBjoXUKeNOPsUU2AkbYws7rVw+1M
D0BeJn9dPsUz+PvbzpEvYzPjwx11NtLBG5oBAbYA71beqxpPQVenvpgZY3Zs5PjFcc6WghQZSup2
axtA6EIcHZ7u3sZ7P2jBKrnBoi3uH9eK+t9U4JHAZSju0k64/k1yPhcySaN+2MECCgccWZmoElgd
T2ABcjaIYyRr6SIh3foFnkJUb+1lsy5ayew5G/jcNEMxCEnGvybaxAtfcXmSIH0y3Pji2sWblvat
EVCpZM7ESzd/e50XHdbbq8VabXxSv1eMGE96en+hxBs6EnTklrbNLiBhN6ijGkssOWULO94+BkW+
setvxsbpbezgRlqv68K3OKmL7VJ9N1a1tezujzzfRP+R7q+RS9l1X8neYOBsFL5XK38peNNwmoKt
bKE6x0ba82MMlrnhc2rcxOT3oDOhyjAq+Ny/BJqczwXOdfTPPFJeA7xF1SQwDsr0B+3g8rKVEju3
5ldFEGC3gyj7TjZyNw+ia6jp6ata/Pl+GSbCResvg09q3Cg3V7BsUO2ZLVtYYTKwnhJJ05TB98v9
eBOeZNrjZEuCbvI0cfGmgJNFw1MjJaZPIzEAbtpiYVjCR2Y4FN9y/wHEH0Jdrpb8XcRJBePORpQ6
rfE+npl9DhVjfbHfzZZlU17B7gSbiqe3tZgm1jtQ8bAj+6uD1zLdUftL6atLZkyuLpF7QaDkdNBV
dKrNy/mXqshx6MBGlOZ7xIoFQNk3OHelycpN1TttsEyHTZ3CLV1oHpFlXWmg/qw3QQVA8v7IntX1
nHJYVyxqDTM6Qe4gI+CJJmcmkfoemSlcX0an+9zb7yyzkrfbeU1czf5BO2lzMJc2Ifot4vzijasW
lmMyafFS8iOrge84CAVqLSCRjITrtGbZx/jbi/m6thN5OEsMmn2NxqCUAjwvkKXtselDkpeoAzCy
k73pF6qdV+x+YCet1vsS5utyL3bpYfr4/0LCYCdL4ZZMPzNk1Lq+Ber75VHAjLjM55YMnh7I8/bU
xQnswxx4MvPNPyoZw3rVbh5qyeqzePXgWpdwUowfTw4u/ZA74seZ00fcxXjq3rN0picMZyUndF2A
0hIYfLLROrqjS9KLsYVUZjoz/plP8iqPWgcKgKQsYiBg4T7t1gxoMF71NE3Jq8YLdzerKvEwQcCG
/xhC82Cre36e9isdnKoTGXBVNQZBSMEyXMzKMZlw3EiVyrcIdhr90aQAyJTwSO6W9tbte6YVb1Yk
R4jaZ8NexJ4vzuPeoxVlDYY1fUP+0pEM8olYX19sKmfVkc7LP4KEYiCRCvofVoUsIL7hRQFmsE1v
SePlsN72wjVYatGdAIsWXqWcH56Y18w6iP/m9PmFwE5L+h1XyR89gvPjj8E92FO6IKgQYfQuOKCG
45+u1Xp3DiAFhoFgG8KqrqmxbkAngT74YQ4jvsYvUaoHwMefLsKkApsgIRzBXkqJR80gekGFR8Ol
a1Zq0FIP1c2xTmASc7rkiiqWnGBb5aSoT5FThMkyPHhKcRef80w60UPyFmdoengwjuw9Q/nght5j
Q7BZp/aqhV8ZbCkAXDKpRHi0n0oynz78awfdExSBvgHtHXadeF5/dFRXX0vnun1KZnNJ5FShS3dj
655/Hc0RmwsmkeVSB1K/H6oAgLtOgD/qRQpaafKj8c5JdsBzqOlbpU5rPTwABoU+4OHLbGdCzS0p
fBlU8Itq9U3YhWyoudm19Yk/U/9PhlDbT+pVuAFMuO2OT1Ov1Hx8yPm3WxcZl9JbhOcp77ESvtwb
qm3B95pZq6LihnScZwefPkkBL+u1mtQ4fpptuaOG23V3W8xlaQupTtVrA8hwZbRSTt3CKCu1Dfnp
YzwsZbC6ZEGvof+3Su4EArbk2NFbYd3AVRUIbsDx9C82BqQ87jIvOaSdXn+V8SSdrs9E/AN5q40P
Xw2VMvsgfStw8E/1i3Ha5MjklbWIb4lsFjsjIPFSEJQroEWBGPTJ3nPflU/SQTf4pcy46Zk7Jz3N
nq4rSepzP4yOkP4Eu0VproqfIdMqIdltWaEciOquplFWGGkwq1+TThbtKgzdpfc3OnA0cqmrgAI9
J3/1C2qMNgSEMyv4idIy6TAruwBBJ9iR1cW9KloSFsJ4noZqM6eCuf1KQ00/7qNUM3BRcvh4eUOk
fFP9Kwk7QbDvYGLfGKr5WIWKXA8oXVsBWyA13D3JnRxL0+siR2I7XKhG2c5TJvgHydTYbjRK7iMR
Dlyl6NurIfs4r7lUCU8DBgxiaKr6L+ciwdX7j2jQyivGUtHFiGMOFfvVWVhNy7mUDdLmfwQXo1hD
s6n65cdq3ljJXVrMTZACBdGRcSCkfbO2dIFygTKwkRl3a1AWCAlwan/w8w2xHaWUf0I5RfcSZI5Q
reLGP9rsVzj4Kj1fvSFgaZp6Os3UPNuFOkX3nl4sHIn0HrjeARpOkWtnHNTl/PcQPncvx0V8Z8Pj
7tfAKnJR1+zYYwp7AZObVugYjEmqtmtZbne8q795B5plR51zzuLxT3He7dPXpUmCgSmpamOwwCiS
nCtUtD8KzmtId/hea806eS3AUT5XB3nZoY4NBDn6Bq/zhTpAtFsXPfYWVnWBUISW49C1nPVKcDgq
RgW/EH8rV7Qc7sHnwXNjkUdzbrTZIess2wUlC+KMsNnntgFTN0eG1EpHActdteQS1D/mFgOEtGxp
oLrSDa4Z1KZo5PQjiFkXP+eUFhSs1AqbrFCDEs+3lCE6/+ap4Z+SGwVf10AZJoc42G3WCRXAWg4H
/Kdfe2FGD3sQVRAah3bqgCAB6YBdO2IUgX8eDwdcYSANz2UwXLo+fEBqJrYy8j9cFK541cfxze69
EwFX3r4Zl/LjLWwwPH74ScL9gZ+PDuVt9hQihpMvW5DiMNP67zWDFYaMK0Tz7hGFArcjAIr30cgV
Ey4lHpSVi2kpmE0crYaxWBqEiPU2wsXCnyT/Cpi9fzs5JGkRtlUWbdrS3CaKdsFuSFbh6mUKuVmP
17I/RTugVCiYlzfsB7v9d5sgm/eXtV8nB4z/ZF38jpZIw80RC3euzlrxQKV70G8ySGrVmRU8iZ7j
xAhCgGRF6dBd3PGduuNbUFMuDeaqJMwRb7kAgVqGVK2NFgIlrtwQZ1QguYb3OplNRJshA0t1fn6K
Qwv+F+jKALzTZQvYG+VWcybFsPJoEcMXkdG4FKr4Tk8x9Flj/maqBfPteTYkEBs/OI35jD26lOjb
VBnhjYTSnmsq3hDStYXBUvmoMd7ePiqOXPZIcKUABC2nu+x/zYWIosxeYTbltEnzeTk7KCzk38Vg
p8yHO47EYAiulZdw9BulIdyucgpX2VIE987ufnMEFdsfLMa/V5ec0ydYkL3gs0g0EiRIoxnKmN3f
bpAVlp9qHkSfWIwgjtmSIw2WgsqBYOmAZdriAtPWQhB1R7CaWH4v6epUjeMdlMqOIEGWEhoKfaDa
XqKHtNtHxTH6DZ0+7V1uP5e9q1TNkqlsjBztcScr/3w+xszbmwQcVojI2rd+7Ap+dg8W2jzclsf0
f9YVeYyIbfu1igxb6WInPOcVKY2FvapdwF5oW1CIhJLs8GF5eCmuPOleY+0mNEe1AEr89Nhhf+1J
y0eZgvmz91ZTRclaiXyq5MysoTO2EX/3wB59Wr9zSYu/lgGGxjuJQH43daekA3FZlwum1fBwq04X
wmjRrjwxzPeqKhhfhbKSXQc5KfgrnZoVZd9+Tw0n1DBvnNY+nIN0YgQ6bKIaSF9VJdQ6mGnvFW0m
xUSIfVEBrUfkLQIza/zXCPJL9Sj7Wd5AJXbxWm6Z6txz/HcCHuRlSFh9Tq6I4jQsNlvrPBMcmlFg
7hFxUH3J8AnFLnA84cxyNdUOhDObh3RWBFCwyEbRRxWOrRr5OGLLcc/5A6D/q2Bvo03o7CB6K3y2
B7YOVllWUVfkI4hv7bmv4k8sagJk0N3YIqZVehNLp5xq7Sh7ec6N4fjCF9oiSbigDJe1Ujrc4Ckm
ZPgCuO/QDGl8EsgWpeln8lL90gudKOtZkAYe1UDpRI3VAPqDQEl2BCAd9JvqjRG1mWtmXpu0PSoy
m8GfrKNtIEuDeukX1EH+1pyljuc68d8eeUfyFtpBsKmK2C6WsH4TEcTLuE6To+vBkDVAlhPrX1h4
46YPRQrk2HI/nwodyMxVeysSLnWlCOK2Q/kBtgtRNOmUHN3yjNatgHbE+/qSXgkSTUVOHpKbWiIZ
qX/gtNpX2hGCvgFKSMFhJsv9LlR9t3TKGimc1KBQpZuu636/ox0XQg3IMm6VZZSmUp1QknETCxdc
wgT0myPoo2i2Zq49zwE7BQx5bhVy9M0OyW7TXgsOamyQeGkNFMZJdWl+wyyb4nQFBYzlfZNgwxca
naScCgnm8l4GCzGT4c1zY8uLxbInnoqzm6vZqfMycp1kbHMWpoKznVzeKn2CwG1Aca7CYoEx540G
FZgdKxBigOqxW6J0ZTszgDL5AQLnk0NB0qTuE1txaWHd8os/CWcrAteXEt3VKQtKpelMqKJYu2PR
e8PC5jIOuDbHkvH5hSmg0U67tOW+Ddz6VSWDFtuz013AN/6WWWZNeHkomJ/Bjfhi5cVSAkB2cB8I
2X+dIdk3f6a5E6hvU5Ci6aCjmpa34Ma4M1cdjjSRmTepDvRah2NlTM3EjX9vRkaYrdg2GzPxi7Mw
PZNYrPLqQgQLP3WRbl6R75W99v3UfzNzIOY/RVERTC9JgZwUlhhHS9jd/5fPRHJ2ToD5LLVSi6rw
i9zbH++AmnerwGJrNCn3lXd7hRLAuXJYV3i2S9VEtQ+HwbaZfitpol1LPdSPJ3YERlvKv1kwCZpP
UqqTGJVkn3CDIhtDNy4AsHKIkA0Ai6nOyYZID1lg9e1dcTZsL0pEsHDrBJ0P6jTbtwerB0enUogZ
zFOoqa0/I3mDu1lKaha7S4XoqwMdK0G1zEIizCeqUzQn25oaaewOwsi9ojwISJJfQiONNIXYuTJH
pOrZbqDfR5plsY+ksnw8UPvOEqyClw0fhq/Iwm1jdVT8LaMPKr1u7t95c77qr43ldg/VktFd3VDk
0YEU9wjFaTSrV/cq+wnkk9GT85Jrc3cH15GqIHVRZx3+RoYVoXPtXR0P6cftIZZldZ/vQgT33KXt
T2M+5b5muL2pTtpkLE0Qp75dx2ZeD+b+vL9mn04gV74+TeUo0RbvuC9hBxPKpRr5Qn0/GJKFzjad
aOGBMGOLFEqSNBinl0gxMxc34TId8ISsYjxazcvjlPQPxg5n+Ym4sRhmPKsj5DpX/c8SIJd7tI3l
13JHTiJKFWQt2Vgi+JqSDzCwtLXgL8YWkUKpU1oOE+bKD5L8n4h5vMa1LrGLIneGDAhC/zjeAHdG
/nokB6XBrxM3y6t+GaU0RI1JwwKyfMuRAI2KVEM4T08/BJwH3uJnP80NKSZUxBN2ly49KUkPfOX9
VEdYM6Y1a4ieDL1tdB7GMkQ2y5NtON2qnRIb7iaKdLR57EL0KxYEIcCMhUuyCRvlzYpMqFP3LT3b
vkrXwjg6n807Gb0Z8Lk/AcU/J55blWkQr4IDxvV1aTIrJi8OjoujNGKzcw6iBGRNBgbMJ40MVAry
mvZ6ZrHxJ5+4BigahTozIAzvzDo18rl4bQ2NMRujM9Isg7DQwJkOZtgRarG38yu5YtTLsJoN4SsT
aYIoZJpCF7gTDU60g7mYZNM50YY4p8zYBhH6byoTou8Yu9j37/DCNk38fNXQ2HLWAvN9di4PBgRO
KSis5K8UMl3L+jWnTT0FuzwedBPfUYHINZTe3i4JG22hlSMsfJTSsuQk762LEQHJLAmmxn3LKdqk
aXDH6HyBKaeRZGYUkatH9LeCsAc+LdhbVnA4EVjxBruXjUVoPTogaXl7e6mC5twDs75/41Yek/28
8tZSoh5RKB0qkQrYry4JwSXzHEevY7FSlswepGfEblzMinTu0wRT6RK/R9MqiFD3QFMQdLHU//Ui
g06S/6691FNwSJlQlvrb3JmcDXBlqlb+98F3TpMz0RK9Ii8ejiJaMKDiluPtWOrA+odxQfM5U0/z
40+Nz9PAo1SXF/UBluouNOmFecTj0tW8SVx/4cCzr1L5Wp/ztpERGZn8qX5QYa1/AqPt7mQegxC3
aKng09ZqQj5Ubj/qDu9XsoJRANiQ3kYwH59qH9Pp1sNXu9migErWOv/yx9AI6zKpmQP/sThir/Hb
orquVaR6h5t4yB6DAY8Sy/ij40HwgCbBr0BgDT8mNIV2+1bKiOpqOkJyeSaPf5XihKTAsb2ESB1n
kKokUhnH/5RlJE0Ayk3TKHIJVgP4sGTf01sRf7pn1sNBnNtd/JA5A0uhBDJWR/LZQhYvjFeH/03f
Jh+uiIOmWh7Zx7nkDXZhUvA7q+5qxTH36lOyXu11HjUSH9fo1i5PL5hMvtVmO/PzqWphPpCq8eE/
KW3L5rLv7JdsuvaYRps2Me/CvG03plebN+oo/22ZQTtNTt3+NkosPLPxHvHPiPHyjPoB+MjCPyd+
MqXiVwINzT4cv8WC7ngFXVwjNdZRdlwQZnsknL5bTp26aeNVUJsRGPUZIn/jp7HChKzZUjyi6N/Q
IlK3+k5ISfS4h3jMM+G2ZMVDdlEZ4it9j4agYC48xMGdY8AVsVvbR0AnlkqVFfaA5J8VY0gB/b7r
FRFwkK2/GEVapyLrY7sMT686qbV7hRQHjO2Y6RSfCEO4Fd9AHe15Ne44KTf8cJsetm6uJNpIYyYZ
LZnNKdB1jKkzn+uCLrRnpmNzm0E4KUmmHWokuCf6wUwrVQNDStnmyFoqOj7W3mDG8LH7ivJY118L
pAz2g4ECbs8+/D/3WaHlhSz8DT4aU/oAKxGTpVBwaJIdQRTuhfTDupsSWqPxv/z3CpQeEgLS1rd+
zPRPYNDgBoSsc4KQ02OAX3RNsU98Lx9uaPnqF2LCPVnqqCUqSpgF3MCIpsAYEMUptMDKcfHeLbbI
C3kfUbXTmmawnDamkjJD3OTHlwQ+GFHyhzNqiNfSAPgnA/G4QOnBTNseWWWDrCGbgTu2/1Jehir0
fAZH93nPzrVWeez4BQ2ZrOvniSutIg8mCsOxEh/CmhWOwqDkVSRjDL1XslH9NFzck392RDGtcP6C
hd/iuVMtoxVrmWEDFn+nC8WdR3BllghAHz0SfRpiw5mcSnW/gLCzMm9UY0W7JMH8RlctwgPoM3gJ
d3bNToaKcMuetFD8F1Ftz6laLMylnp7U4olgxMTsejmHt+hdbsb8fIXwBVK4NORnBT2hffk8uzV5
kdCTYwMHfUwWklctofnTRqCwWp7x0Ti0ngOpRcCiHfWCCQppy1bGFFo2gBAc6hRLfEqK5335G3x1
PHnNtNaKjKPjLVeJGie7l/LaQCcDH6nQNL+0kTmYvHxSvkmOdbmnOeBfUOIq2XM3KZZvBz/XviWf
+h6M2T6NFxJHeSQc4z8TLALrWffBtR/CkYADu+1sB+pL2wXWPgbVWQoJAHKjilDsH2c4pQH8NWiV
n1mzseMtYB1Q6vM4OHqp47Cg3ij3YxlSeVcr0LGgdGamLVk6VkmWzIYu5kfoobiD4UwfuzfgZpdh
OYztwLCr0xHX3TtBox2XuOaZfqDR5Dp55gSHm/Jo7pfJNnsk6oYWpNf9Ri45TiZNxi9xvvK8S6Ba
RkLtHF0DnRNOeYbinJVdsHnmJCJiwSE3gFpdKChUO2SnKNooDWZyJLXa1pQ7POSsHwbWWqdn3xBY
tiCiA7yzmcEBuosMHa4e5vsI2LEsJ5lZTFjXC0Hj8V0vTVE6AurLsiSppG/AqkhxLBKpU7+7WVE6
m/vxRS2pdbxA7AslHnqrvNYyW4KhZL1wu9zwrQMhJ4XlLz+VQvMSGY1dHecDRVmBaAxuSUPuQhx4
RiF9VJg5Zg418Bi9lzVIY1tD+DInyGfuUv8Qh9Zj2yZiwdgeJfTGrWDliM1u6AAYvzhroOVjB++q
PE0eCJKIbxw2qvklunQGr3qvGT7wPxX92GLqGGqx5bEPu/2q69osasv2Cj9+92TJS4t5IFNtYV4X
ek8gjFI3Kkd/DmKHgBsbMIIlnnVqYKTlEFQqWmMANmYRADk5Cb2xONecA+J4ofzP5trUbxaPrrfC
DGdDheIEWZlzD9n1fcUxMdpD8mxn8NVSHXenBnaN1CSD+NjAqUyQyvHJLE/PtlebDBqspdZp9R6G
Jy3qIpDR6IJDiCR11cikWDJ8htlu7U9yjD4QM4Oj3VKaaHRMwHZ+ebJvgV1XnraVBrNpBRyVjcx3
a2k+casftdyep4IIQ3Ew8GAQ87i2c6kF/2OFEsa0KBcC/u45wLWx2KnEI7eFrR7nvv6XWC0t5daT
AdZc6SxNEyVi+Ui/FDy7IzhyuNUpb2DoDm8jdZW3FUmmiyPVk7HjGiCxmDJPzCaWvm6TuuT/ii2m
h7A54yvU2mHVQhT6/e6JK/JFWHNuRhzoyu4J6vouKZiZt7k347Pef7fmnzUW1V9/oKDrihFwpgml
BmIN/fBuR3O+xn1fzV9oF7aOR5v7/qgTleJUxriYMXu4GoQjXyo5QZjjU4wjqjiKaaHrdwp+ffXW
V6sgTb67kDQoWycfkL8k/yqtYdDgnfFPyzik7XwVZ3mEI5Uj9ZjNTxHpn6i05lVQmyCsrqLK0rXE
U+bzlcjlzXPCOqEg/UiPjz52B7qGbS0HA/3CqeIMwkIo1rdpgvcpQ8O0CxZnP9e741DGU4NpLbH+
CxzC8XMZXhunHI0ru4lWN2tdCDTvlB+Io8uM9P463SRNf5M2B5p1X845HBgDdzejP8TdMPxrlCYp
zYaDD9dS/31qFRV9UHlixUoeWKW0G2OJKZT1Eoezcb9BcNyaCsJ8bepitttIS09YCIKVue8jYFy3
E+0lVTRcJHNtSiJ+IWAwna2zQLKlFZr3qSRn172/WJCoWcVI3t+xOh/kCZx/I/g7rDDKV1PymRza
8f4KpHYkqyRL2yAE7bcStxGK1GhfsHOJf0RAvkUj3p8XdP8G4VHPpTd0tWJD/cHDrFpe1BEpsOOm
WhpoSjT0AT78uT7PGLZW6vV0S9vbSid4WGd9y62gwwqXZW0jCiRUOlOeJ275fomOL9KhSK9laa6L
sToIAUt940wk1Ua1yf+WyO00rUGmEL5bfnBxJJzn2XfKz9vHKs6cNoD0FBMPUH5HLvgLzd6U3Lw1
qlq8mg3araVPz/YwUk/KFyaS8JOd6Wyc6XE6+7wAFUTdLvtSceSUwRCT3aehq+IiRamYYwiW1iZZ
XKZMkDu1rTlB4YKKmMMlvTwmlvmoj2pHjXj/bHBfdoXozDBGTe3dFyqsuqWKbr6D1icq9Qh2y6/V
5kuSebEzRxPXHa/XhlHXkyo2jBj0Zhtqf3VsXBAAs3htlHHpUT5J6v25rORYAeBa6ZJ/NtUr+NJI
Bbn4TIY3PIqoYmiWG01VUHtK75qT7kPPzXjUjntAv2X6o5Hw4UQzCpxxa6GzNibSMxfYbQW6VP1E
Ld3+AotLFz9u7Pvk9oQauhoxkGmmGOioyeNaeZjpDlMQgxrP8p3jMgr9PVvtHwWZP29GyIFph9Kl
Tq3GWZiHLqW8A0Bvhnu41ew6/3aq0+ni7yKHl3l4vJnimtJqxLPQVuZcpPYs+uTPpUOjCvZ/BoU2
3zxDLpcnx7pnvfu8kN4M5hkHNodnYSSjJkQk97sxJOS/UdgC4xCgUhUG2qbFNiD05o+aUtVJoX4T
AGiIgPt8lOfHjpzF28NF0OFIFhzB2BgmE2gqUp/QtAlzooz9KNvD6DFatklFVY6LfF3H+nF6Kjca
pxjC2pEqRBXMZS5GDV06NnaxDjGYKnVIl5fKuySGa/yuT+CmDkDmIVLXO1iz50S3rgR1wLNyLyTP
y1YBcEqw4RwQ3ci/bQ+VYzcpI25rdtwTiuEiig+EKzy4//dgW1sAuCOQwc5pSmLpEEdjWKEYVK2p
uD1pN3M2UdjwsqX7bQCVG6Gvp77pTTuuhPAIlum1P7uKzFTlK9Kk/tVxnnZE9VWn1SYW3TSlGW+W
9H+NS390T9/j1o5QSR8O8WVN3gUQhxqHrv332ae4CfcB8UcaU5Wgo1TEQZiiZjpSjtB4GvgzTNLH
4CU56eHwGqfmPfmJlanPsJfreehwhClVFG2VsGjulMW8p/wEyBM8j+BoDB8/ifVKqA6GBuOs+hAP
mJgnMjuQex7jLCfhtJucV2aFYe4//kMfvU9TsAR6L+RXtvcGx40+ttgYkLdvLFM89NsJjfMPzZls
jxS2MRxwi0MjekCPcwRZ45Xv03wfpObIC5Ddu4UMRUQK3G+mFhD6waZzoRM4hWUot7NDPu8do0mt
EYpEeroP50qz6QEQc+TMXKMphOPFjh7O/VU2BYAXfn3HNtJidP0eAZbNPY1GCS7JFNrwQwFBylu5
88LJgTvW5zKwPtFObQJ17nS812rniWSK0GdQazSi6PIdqvMPjVZ0TAVtnjZnUmnNPP4RcKyykg8x
+L0OsOHqkBjDnpuDhE7tbj/DgXPy0HDcoRxXN5i8fawqjo84+AQ6yJZMN6jhox7YB3U0An4/8PMo
M4sRJtSguCSUPBMKDi4gb0Aw2Tc8YFf9+32SWrJEaKOmlH7mYgclXNullk4uamdHFqC6V82bCm3Y
KUxTCAtzxW2rxpaIIpRn4vLMc2ik96xL8xEx3CDeJ4iKFSiZlBzvSCKEdMG0gyhq7ArtXcvZaWfa
IsFOL2g7pQslz12632BIGEFMVhRAw3odVKYkn3Ptv9nRC23rM2OakBrJK9xfeexCjG7tXlnO7vbG
o3KSaaedqwqPL/PPV0/si29R0w4L2rK0uildtYgfCiUtzIZMwt9G/dMjheNoiZCmDUTWW/B0spdr
HCrXjd4nOd3/O18pOQdSjahU53AR68EU0kfS0iVUmMDEkaNVWKrwd/elvdzdixNO2aJwzFUS+swl
axWiM48AvMeEzWdNF2hmEl79xwxBprH8yZYapRyf8hIMP7S/zrEHsqkV+jRTWQ+o29wkPHFFY8F9
qgJPZWSGmvFs08Q46WGB50VzhRZ64alRVxhjs5m/lje+SFYNEzpnIBcQbNdbRkoiipGXMwa5mnp/
hfy7816pzQ029uVGI7h0zPq/FDQSaqSnT1tO90IU6zOoefsFvslnBLl+x9MeFwcSYr+GKFtMNaX7
rLXjOYzFu5RZ8FB8xfekNxyNCECj0wuU3PZiEn6eNdMapZ/fXcOguSBYoLhksX7EGzPGw9A3FilJ
3AfvSnZ380tUE5CYiITs+xMZn1VOoBweV85QML9c2BwrecX6MlH4xmeg8yrFTzq1uTrJewsD6E0P
VMg0Z0DdiTnh3UJWT/S3ZceEWl6voqYjSI9QCm5gLgsq/HOiVcafYiIzfYNkz9sfCj9fA256T2UO
/zAIVQqORR0qs6RweYo4SuBBDOkLCrOeXTpWxN0IgVCQJtAL7EzgUgCR7JvNwydc20jPSYFb3SAT
4JN/l3KSml6sH62KQoImTOCLR2bKhJ4DOHvwPrtfJkwjdm39/QGVKypr9nH9dHr6aAszQFTimi3z
K/V1H9d8r0Y5GJtSm+DdaYlqgCbsl1DYglPRaEsoOqHRpu6qBLFH3PBrfR3zG/nzVpBiUoyoRG2n
p3KWopBho8fOsgLPrmGZxVYCWjhe3zK2CaDh5wFAuQgf2sGVPzSYUInIRgtjyh4XL8XOQLruGWiQ
jqHupi3qQl4NgPhRJ43kmkIwcl8egY/FUV/R8xVkStYqd6vLd5OmWXx4pPFId1CgdUFoPGvS0ecH
VPTsgESiJckkShc1onS4Mai+iDfwrV9tzu8gH1U76LnwZxKMTGKIdX8fJDXhHmr7VIn10I1IDwMD
xipE4ySQVyWbFfABy+RQWUozS9cyQHP0MFPEn4dxByea8yXQebm0e5ySf3rJbei8I1ouNkd+rK+5
N1ndrhK7It/wl1s9VdODi4qq+2s+dySt/DQhL+PGykWnUrrsQX/t8ChCR1J7gTai0zLBpsEYM4UF
jNcl3i+3bryYBqyMPDV3EIBCfQMChDOK8gioyyMRuApP7lW2P0QeK3PLTKkjjLcAUz9+DHJkrE4u
fV1Z3f4JI7Eo8nCA4UrJ6pO0pWy+IZ2tVrr7c3SMO2VT2/D/OD3kJG3YRF8ffWyqWQVS0sD5bOX1
9LjNhPNx2kOgIyVseg1b/Ik4sEyT8/S1DVEawTm5X9uK67p8zW0s8ZFRaefHW/n7SpK41lZuAq+d
A7NnVUBgw5kb1rE4umabVCguCDJ1g4nuB8LMWeXjvc/F/ZaGPR03uqUr8o21qC49YVwGgoFJGVAB
Jiecs15cc68ssAV9V+roZ55L290QhYhHCCXI4jtXXAVtJA3vznrCu7wkZ3Z1jah0l9LOFrR466Gw
TGlnvFEW6QeK4XCPHoTW0KxpZep3l6Qqw24DEYcpXQcj3DpHwIWqOL4LFXOM4wjXfuTbg83Zbuls
jE46SoIb6ja5gngdzc82735X5cDEszCNYFmhNgXRV39wDIWnIRkkDT42ns1g/dhtKDha+RfaHC0y
hb3/PJf8Dnu7VaEwIWpC4XxicmKlk1iqvId0u9YVJeMTWPaI9Z2ItVU0d1DBLK8mhHHr0xR77TTu
1RehPaCWahB6jtEOBGN5X6+r6dwOykwFVrFU8xhNeV9A6NSJuozk9vlM5ZK9ZzGdbboh1c3GJGMU
QmyHVPqnXBG34ksKzobiNr2x/3mbTms8G0wsAz0oqk+N7cxXE4DC3Qw6GB1gz7TQSUA7+Jif57TP
ctVncwVP98atruvh7HJxbuspC7XSaNgnh3nB3FiAlDBp86m24gphTiejfOTzIAtA9c6JDeL/5QwQ
IlZL6FL+zPSEB0mRv/r+wbu3/7MoIOHh9jcrylfhAIWTXU0dxoRCWOsRX2UEXAYhuvgBwvSz819o
ACbu/9ghQiG1lveE+UaUL4z13qYyvwdHzCMjD4ncp5d4Q6jJYfEwHQsbzcKZZ/s1Y7UBvrCwtI6L
gblGZcedee/U5Axr15hPyMklIbW6acI4gx2a707RdCS+TRLvSDRErXpgjU2Po8NZOMMLIO2WNVWQ
TJjq09l34T73y+iBKyFsLZN5MTVIDLG4Kcg5juMh+QaYnBouMkeUeJBChldi6gs3hjeEpUSG39cr
ePxOQjBPjVBjdjzLGrbVi5DvsIDVSZpADBd1QTDx7On9glXnlkrzTlB7QBdKEFyImB/aofdyjy2i
KeQKJRAiQ6Kwqf3LL7SkyTA91a+xnd2Gn42+rhCDvTNh6qJSra6TyFtoXp/Nt8r2784WFevTD1J+
v6At16oAUCimqKzzEQjaGl/zZ7ucKB47LEmEwrH8EVLSFte/s2jSu/ZLB7JXnOGfAgFw98VKC2oN
6hp18ZdoihIVHSmPCQCCAOZrC3kU/yau6tKtEBcV40LlS4HNspAh1P1Ai76rp76/aT0BcIDtt/bk
w9NQxFpbV60XW9wurR3yZLPaSlNWrT0n8OzXuvodDVfAsNrxXEuGQIF/qfk87CeHb3DzLKwt4S2l
u/PEr7yoSf8qZ8XZ+t9AgbXmmBecJH6ujPJ4RM1pxFYrNlGuJr2JPG9lE8QnhiSA9kAfzVSjO37j
hlRDXbXvFCa9+LdZTDCrguh3xQuydRZELAseIM0uRjfgomHGZbmSFbGcq1ozyT9O69g61VTHKovh
g7Qiw3W39CNk/fsYHJzEBofluzROG27b/PiF9Q/Ozp8VZvlfyqXnA7U6UrXe6Y1mvsOvktJq5HKQ
g+R0YHEMofEURrosrsqdhJnO35jekYol2yuaiYclBzOotozs274+z/RCPtGDeyLPeYp9EKaJTH3B
yKpDBDGAumzzahwDj211BR20K/oSE30flIKcRPvAz5qCCelsWdT1EJm2f4vtDg/wlyqV+5IvJTGZ
sSbiXTLJEXYld0XhwmwAqGOCK4YFcEfW49Q4GxACHGT4V4BPhZs22C/auvZTpZlbvwwV+iyU+6gV
obAKhOn8NYsgh9LzCrddnFTzJjmERHar3hPieZHOFVWag4IJaFDl79Kzim3kEm10bLEOD6DhxMjM
7qWFcSecCAFb+ZZM2enWz9owlzcpmCKfnWGvTBbpBySXs7yIQU/9Lf8tLCDqJQPEhCHsCLowiSZO
Di/M4j+haLfmHO2MtfAECq0/3SLNrHGna4pcQMm95MmLtYDg6BtOopTRRAAsF9u8fBbqbrXQX4xT
dY1MJ5AYTqJBnn8IzqGSOqh3LZNqctbfmxSwSYGwpOLhetB3WxocgQ4+Xkul4BTgBGI23KQ0lpQD
yY/bk+lwFYZfRmxdxgXYMDHrfgluWWhKOLlFh5cm/CTzUCYQesNPGlyj2qVg8vqKwhHhpHaQSg7B
DQ3pbtM6Gv6gilTJojsk4COkXgaiTFCmAZ2+tUmR/g1ownaWr0gCVS45TgyPtLKbSIpF7XqTRVv6
+o3T2zWP7cEYlvOkbLgs2MI8DadVPmYr+3A28wjMXABiRgzbcIsIik3RtjsIVeOY7JsPtSfwxOtZ
e3DrhYryHBC+Az5ANVrfMxR6qbJWoDSk6W/9tvjZck0/VTTcGdqrcyllQ06Njf5eAsr2waJSGTkC
hXvmLv1mShX39MoCcuv/oHYkD2QkOCQPn39Ae854FePcs/ToTsmEGTJw7MueQToqrGWc4mpWzcPn
pYK3oq71Wy+S95cIee4N8u6SPs+ePa5cwG81VDll6hO0//TU+1kVBwP1wY1lD+Rqftp5nqTWgPoG
zgEDJ3JNa9w4tvJ87/ayvZznv45UE2zDeeCp74cz050RLYZG8ZdH9XSYK22EssGviPLUXv5TDSye
rHE+RTuSqSHve/fdzOHn6Qc2mxq+i1/3XKoH2S+rk5VaV3C72XVtpr9yDQ8+jejCRwyMPVyMQswZ
d649ivZBQdMw7CSt9L8FHTKbCRW7kgz36ed7P9JqY7M6zs6Xa/FfS4wuhoBsFOWpotRg7cgu8igq
uW8l0TZlXhL7XFO8QxalikbexPVc0C53+WY+KBkkW4zsw6tyyzi3SPUjSji7voyxX7awepGfXHXK
XtplbwRGiTAbsPC0sWEPBWvvWDMh1ZgXE2LOw0V38KMj66UeTvGT0YOcIVwpWSh7jzWXv4tVUBOJ
1FZiGx9MhfZQqZrYgNv6uH70aF/DVX5X/3+DTjS6XGaJeEDPO+oOzpa5AxfZsbIF/9CQiKF+nS8P
rxPuOPHxIGFW5lcgykxqwdxTMIh+1NLW6/DV2eB6nIGuqE7dmq9waZpPV0iuEPQfrUQ47gUBb1VK
hd+LqlIhveSFRdfG0j9sGQjufZ5L5KYEHzd4t0es2BaWRd7OSikXEszPERyJLI5/SDraRsKybtmo
shKeTP8aSj4uy8+fyAeuVdtRBLe+K5jLuLNAQnOwiIWOJ/8zLnsifZiiElXFNsFTcalYPKZBU9l3
l6TQxf5tCCLrfbQcWQjGmQllPJW1yql7AvV5od/51M62ZUDAXnHgKMdKrsR4JgmwcbjP/zsQE5FC
p1Se4sQsWYDHSgLWK/Eeoyt/KezXuBR7xyWMljvkxfWTkhKinnNwtqaT/u8UzoizsjTl0ojJTJOf
R77veys4KGTBY0DbVFTxKC9wzZ2F7SDa4M9P4JQWanSo15JkPe6Y0bg9lXFz08CBlnT5FGebXhiV
bDlmKZGms43k5kYq4aKTsse5VVhwLC8Py5RkJI9nL7e62XmiNvMBZPpTzqFVjZBGshmujdRDAi/w
2OafYLWDCe9dAKzn+8dvVB3lAcBy8tNK1BWejRbBUPpTLDfWmYOnX6Vnqzzg2I0XySod5W8T7VGw
up0IoScRKZGXKpxmvaMzj6OAFIvILH6LQcVRNvpogxJl261Eo8p8ddKUl5ZW4NIPqNAtDeWjwS0d
2TF8fA/0kWChqaey+bt91XsBNDGCVnuYv8zYh0uE57viemsUModVhleclSSF9cFL0jrZYr8+wEWL
oCvgz0jCcDWE1tqMbsnya+w8oOnVINvJax6xEmWfE4vcDFjVuNPWeonNuudxLmWKbHupY5zvZEjy
fgKG8YTckX/O1tV/2MTHpJ1/FZ5+HBftZJCU/JUBiH0IS+HGs4Zd6AxXZ04tTfFWDpgANnbL2ICf
S2LSz+yaW894Ii4mN4x41eNLt18lbKUx8j/KM7LL4bPTuBtoxRqaS/WBlcUs8BAljhUDQtsEiH6E
zyCUXeliF2UvHf/K1z9C8uqtsEKI3JOFRhFmGupzJH4mukVV1Mpavvjs94z9xiVzuc8hVdURl6sb
84AgnG8IU320A0olZiSHDxqG/q9Svwsu7YHPXGdrMbigrZ9A5AxYItD8KlgSIA52jKMbIYT2j4fz
7z2INV/gsZpdktnRPAR9fLmxQ2ro4M6dLW5h0gCZHZ6Ao1xk93/sSA2LKNKAoscJlAVt0iJDPxdR
f7iaMcK12WufWGm5+QnaA1iK4EvoFShCwXx1evM/n66/MT4QSZKymUJy12VDCY+jQ0dUFFIOVwrg
BEySHLby4HT+VAtNiI9aWJxULm/y3xhX3u/jwbVsYj4HI0riGTo6Fj048VLddSClncHSItEUxXCM
zvrIN/vZsPkRNeRrI/S2G6AzTCWdx8ulA+SlhV782b+U/kVdD+OAgQtnTK8bDi265IIHD4dXUAqj
fbMFDF1EoKjLeGW6XOER02/KsXVqPTaFrfSk5FWY7ekOOKPz4jOPnkqKSQ+9BCRviX+w6v3Zu/Ke
mh9v2OwtSygX3DnLOmpLsSsnzGADkLEvE+GT3No+nbLYj7sXurv3TkhsVBVEg2BD4KhU/aynDP/l
lYKcW7m6Ob1Vs9u4Irrqsf5iP/ScrjeUBrI7VIi62zLGWGb56/6ItJnh3yCfUGEg8AcPXrv9Tf7t
/TIwT6VboD0/Mc5/6biOkJfMBEpz+0nY8ZRpE6pmK1mNj7bcLjSWCnvMgtQAQ74XZdnNNBtKX64N
/5FnSEbbk3eL+RqHVCmKKDsWpN41ACXSEyp0eFy88jZRoW30hJmEmH0aNmkWq+GksjdTqFln3U8M
gcMnjl0Vyo24Dl10RnMPC1NjkkzP9+sDv1rbSYDmEAlW7r1l222Km/etVtGqyBIStenSYxoz9DBT
nSdU3u12spYmQSX5U7Sc5fMeiz7YTvNRca8CF03DaFGtUe7U/krMOFHdSUnfT4g+lD1d829VcT6s
1nZgqXMFpFLyXNVOg9INi9zTLK6hXq4Yt9o6n2Cq1USNtMZ+eIYC0Vcip0FAu84Vp8nTlwM8/oM4
artmnHK1fq+uFBmHdZeOlRbqZD7HrfL0acYIhDd2WyUFYaDFRivqLmtUkFQY6oM94mD6QHXKP7yn
6ryQuREMEgym2KWySGhcyRjUhINAG5XygSAkCh9ImZmVdKvLTavjUJrZVJo4Qa8CUjrxIzZaUOpX
9+pJFGm/fgOIYTyYzp49gNJbSGG1/XgscIS6CvthjSjaIJ6z9y03UHVzgRgSF7l0XHm20u9S+Csf
5pb5FpPjaM2fc+HAGABahWiGFmuYRn9PmK3I0mcgNam8mZMGhzU04wz58FSML252GbX4U1xop0dC
4hbS94HsJpbEy2c2nEXcwyI5uKvV6AeecI/THvqVrApZvNNW6vrdfqxckqhKAURrH+zu0UfX4Bf3
X/oBe4ODsI2JhzY08U11Ekm/N/1UBU9w8SqeIQi8tHkbg3E15ui5nNWV7IlQf9uwVGS2W+r0CsO5
pJHuXIH3dsXE7SgbpkymNc7p8zZ5Pz5OH49MTIiU0DhWKz7+/qMxdjRzqhZ2nVrl0xZ6r8gBneqM
4rC8cqOy4ObiXofYmfKTN1SUAhErnoXD6IO+jMjKJT8IPKR+L/L2ZGDhQ6hSV8gfM7J7vPLKRPXd
H4/d2Z9Br2aNfVhclH+ohIg9c1YiJP9ZCsyG/Uih6StIazlw22iNbM8ClWC5nahqiScXM1yys49P
12NdpYQvD/ytNWrWnsW2G5c/kVfYVFBi341unDJsCg2q90rSEUbYHHhKAa+kluszBnCqx4HsicXH
fn9QE41Boo04it4qO3S9VsSJn89daRak2GHfWZH7Cwjm3dYzRGbtCTow5TLT+mGYK06+3ybDCBiZ
L6WL21QTtmkvbRN5WSOKqkDJzrQXmWn6ZJXhSGE4HxkeNQLq9uEiOpS/g6Kz5FlskwENzCaZlY4s
YIZ3Z5XRPOgUfm8Pb1JQYqEeRX+1rJDZEnc3+p+STNBIWEp7C2w2aZMDOVGqCV60xBBLTUd8Ryw/
lUqt1Gt/vMUz4ngsKqGPYUd1gLreIedDFAjSjzDSTZD8U9VslweZsBsYvpou5qDDEryh5uQ1OS8z
CEOHNBSBYfpeEuKXcMSEk7S4yVmfHfRquvnJh9io/ZTnp9Xkrhsk3h2Jsfqe6KflTFpMArv4bQ8t
qe9c4sshIZxWke0m3XkaTBjEOkToBN7GqDaLD6+Cjg0oH0AQM6LZL8yrSviDiJYkOGnNR6b2vkZF
pDDQ4GEw7B6ONTYgrwaSmKg9Pa7m4xTOi69bim2Bbs+3XA1EWkpFQm240GIJjBSWpVsIrru6zP9l
vPCKfa5RKqqhcj1ltMJLL9iAiVZif1W9vnDpqypE2w0+J9xFNY72wa1X8QU4oZy9DOvkOK/s8cE2
Tg5ikxiOlywwZ07YMiPq1j5Xxlevbrg9AAB0esDj7+MIXnsaZnQpfZjTtHDg17fw0CwQa58D4HuX
SQnP3KdaaxgcdBTsusezV3gbKtADXkVu10JCLs60rWTKAFp9UhtZeSt5C8xVdfSXLawWBSLaRf64
fFNO7qPJ9bvCxAu8Sz7K3KjVRaV2CJc3ZuNQv6quusXYxdQ8vYkLDGyXo8wf20ukZTBioXRemebw
8EodJ7KqlGAen/pf2ttQXhdkPPqu07M35PXCBk3PNd1LO6rO0OIn8mF7Z7c6roJpk7L1DnI15deM
8j2cC+7P9znmyUr7fx2T1xRA+QdEVB7mJa0V54QybHYArn+4rROCydGYMB+jSdhMDdRNTjahoCdg
Sr68YbAZ7G9+1g8WCXHlPegz362U4PKBWZAnL8889GpDPNO83AEE0x3nsDoEvtmAn6L8eIO8GGS6
Eb7vfcMjJF6h14dmDOFF90T4zv5ccZOz888MUIHlQtyqopkS1UJw92Swk3WGbFKlbwLf56+vvYXy
lfJwbFOiXvfp0jMl4zSa1U+BXv7jgD5HdvkZGnngnm46v2tSl7+BA4c4RSxF4pfjsVlPjHvBtWSW
7cJTvqUzfzVrDQQI4ronCGdgfAgTshrQBjharmAUwD0pyKFgqdKiWpUsrya76bL3cTq7Z6bnP5gd
JhvFhwcz2cqGE+rnjquVtCIWnJtADfX9JxN7uUC3G3z8+bX26DruWPC4k7jylIN9OvUDpE7rwfEK
U7MvVY0nNrDMQAii+dhoFfhq6WyAh7ws1uDA8yL7hZRTKeUT0AnfvBkXSwIeHn294o2SPtAE76Hy
IHX8pfr+2UeEUwZYMu8zKZPtnxsXMZuoXbU69ZQcbZRSHIV2rP5jxeHcaU0nrsF/EjYs113X4aXw
sLEVPMgu0At/RjiMkzdSgtK5+zU3DXmGN9bXP0cAKbrmiUVB6N0DJzHlzCqnxSveLd2Uq+me00mI
2pHSPsmJ4nTFOSYaSdEfdfxHph/6M9Xvp7tRX1kXIcyrzaSs8YVArKBLn/AD5bnyrombz0wZtHbt
FK1tjnr6VJS6XcQI4suOZSXmnavT5nScLO6ssmkhy6pE0Hd64n3dE46jb7gvobuS5aL9lgb+qRAA
ZRJzT9zOW+L76P2TPxo1Dbo8Sf54nygDoR+3FiyElDlgeUPlguw2A7HiUOhNnfLpgJ2cwGFrngvA
GRdp0IMODAwOdzPiRbIscnfB8fGtI2HKFvZDhMVaW0Xfh1lAzSqyYYgp6bc0o9e2aCG2w3+iRbL6
PGv+DNFopTlpA2+JGnfvAlXpVQtc0Yc5hrHy6DlWOfG4GC2D5tbWfhvmnk7ivm9cQuj83shEdMov
tiO3VVn/jknleYnFAGZrznBp8V3kZicJBnp9AuQ9ELp+NEcjxvVx+d63PFHk4pRucnWNaZ+afIhw
s1ULs84lOLzLNA5RcN0TCk8UVK3k5Ae4IsloA4ibml6VCA3cJ3HALvEqnSQ219iLKWmUpT9q42fY
PMRttE88zGSi2nSkEkJUkJ+XUdJzdxCbTx1Jz4e1yPbhtIzl/1bD7hHHHcai9sdJPGif9mGiHqmW
qoB4X3ZkJBYWp0Re6DeZZRpZ3kdXaX3gVR7ROmTyI+Cc09bU6YhFa8AjctWQKkBQ/wUrkXmajHUM
t4fQP3g37bk22/nlDVbjB0DbLpY/9Z2cy2a23Pca9aFJ3AZyZ8uCeahMoqMJXuDOOurQbXbiOoz/
HE47Qtzl2fFD0fyjHIoxYqmkM61YhkurooXTUR4mvat754r4+JIeH6ea/R3ldlBhr9nnHATKCFZD
nEsIIIYFZ3gjpDBd55zZ5oXUbItKIdoVau+2br04YBNuA90c3UmG19FWpnJY8JbPpf6vo1JL4U69
tUWURbVvm7/DxRqHD9BMfFOPMGzitbU2lVIPKTv/Bmg2OZRGG4szC9ITQHXRHRgKgDhwsG9HTuEu
Hki8ect4b7Pm0pAEDm5r1b+nDJQGfNx0BR2jogXiJzNyPpphDFpCWUyY6z7qpWydHB8oZAhKqiBa
bTEBMNXTnVefZqHsrwwRTThahjPl+j6ZDemdmOPjeJWoSeV3IKQd4Y9X5lg040LCNAJYfsAMNpMD
f71I2Gwk6djvPIgvz3gXCXz/PCG3Spi3e9f8Lhg0UtA9eKGfYZI0n7fdolZFgPJzS2UJba/CuOrK
Eii9RnEBgeLYOdmF8pS35TqcqsM/NvqjgukCRNuAe7fpIiD+2Yal2zf7+HqqkjIIYKEY6+UW03Sc
RvmIQDHyAro+290E1WfjabyUKpCrwjnS13c39uejVxfqmFEh1P83Ux1EljVLZlQyf99Ne+ebrQnc
yqsNMpg2tliUvXi8wysXLW04NzKkNYXL2p4xdAvNqSoWH9hnedQ6sgPpcWNOmByhsOvlSg8e/MGv
sfXsV3bBqZ0sWKP8RyPPwiOJrD5Y9Qpcwysn70wNYcKxGk7EQNvWi1CO7WarNlMfG/qeJdEpTT6l
XxJBNC3p16N90BZW0vj1clW6e8QRLV2rh6hKGiqVhtyfUZ4Usqm2ypzdLf5Vibnz2qeP9lZl9y1U
QBq2pbsJbsdZNVi4nx/pkwqSQszmbLsD19CD1T6Ebq767FZg60yY42HhjbNFzw9wKb6aGMU/9Nng
GApnD7BjTURci0yn0ak9FPjOs3FV1ZTl00E0XGRiis/bzvly7csMasVsDOd8BmzlsxYTMvhH2XLe
ySlpa0DLCTXyLajQJnwU0eiPD8A/9LH+6tBYCQ/ggM3F1tJvDKMuvgd6KOIu8ec1aFYebNLSmSIz
mSVauvCJavIgg1zAW1Hdf/u8dj2OOEnF5G5zziXvJ5TugpyNqmgtUnFUrmfax7ehQLcxcect0BI2
m08htAa7dqfTFRnRmzbOADfbyKcpXZoxQZx6Mrt1jtv9FbMMHm9yd5kPJIiqVSKo1XExCacDGKM2
fEQExvUDzTry9cKoQaeP9sW3iaoZBLKd078VotCfIoI6iGJZ2K9G7pHdlPNUnU/QwI3adsfDJc1c
SKI3wTo+uWzSq5Wktdpg0fsu2uGssfh2VYZ3fWMgJqomSOHZUdtktBWX9F89rJxcVPZEJKyO+EAO
77KTN86PalugBh74VOXviaYs/U5OMyNyez48s2+OXWDIYVkMPVvxadgVzWHMQQXgDje3GKnPi6y/
egVkJ7rS+VEMwNMkulu3dyDsOjTF/9MSHXN6Qvzao3Q7ZIo51kXQw/T2RKXd44UvsSRImu0WnHEp
oXtfSVC3TQEByAzDBIsB1lbVAGEV+feoSDmYS0sdfB+cJQepl8VOD/dK+S7q969VmrGHndoXF065
kI4q35HY4snFEYcYWs4a7GNNCPUpW4av5zz7z5KiGrHSheNQ8KwSKaRGCIg9LXFVC0M2iYC7XoKB
wTZR/FQlXSuqZqg3njA1xUblDOYDkYwE7LnYSDkqNCfXk9xqj9aF/62d/gkiTtP59S4zU1vlRVKI
eAdQ46MNlHNZWvB3HRv1ezZwvXxZWSVWActLXIxRyyEQfk+bMjzjuZaM42LtwkJc9J99xfJ0g4rn
61OmphjCyYsr6PiM49mp/yQuQzQXkgpgkcpNdB/CjN4xJYi91cWoYZMu3UCv6t7g+oGaqe+67ElP
MBKcPys3f/++K0qX82JFfV+PA6DqdXgrdpl7kbCrXQgFG80yA/hBEp4n99JwnIhl8wqH1PKixQBg
7aePhPiNpyRUzC8WhPP4N2AhPPgoEpplU9Hbs5qdtJ546dis4fIJrNcBNVRRuWSMKUJYxkQ+OmOq
sZUOvzgHwgygGW4Bz/gqrk54XTuvqN8yrezLgp00bYxt2ZmDwr3l+Bf90jVQU1W2EqRFywEemEVg
AloUxoCJGpKffHwPwLS8w6kJhFter/b7KN3VeLH1shPhe0wYez7yLVlykGPSEqleFTZ+XU7Iyp8S
ZIiN9kJ6tvYXDMmtB1+LMdUl96xP5yXUno/U1AoFPoZ/faIw3ys0Ckk9crpvMk+5OP4JEwNnVtqx
cR8DMcELh9+C8pee7hnUTp9FglHKbSNYO9Nw9mYQKvmt3EQwK3BSM+yYQN/OgTT9JUxtBifC7Ag8
G2uGwMpEiFz+NyE/t4HizHfLMHCtGOQU3ZEBgVJslGyuwg5jg5zFL+XWakQgTWM03BnGHnlFtnDO
TfiW3z7Tp25N198WoOOFmY4tECzkyBlSyy3TO1pdkRwPypW8FZmOrFNDa1zXVSzGpAX61nt7DOO7
yhMBcsm3YboQ4E0XMHOQdFkc6uXUnzD4CzeFQ4eiu0ci4fN2fCNnsTXvQb3VROutq4zTO4O0t0Ik
7y3eXgtunOK0rXcsb2ZEFWJo2M8+Z2MTgmxXvEPxGVUhxgfh15ggXz9QgRC4N6GO4Z7Cag2zEF7P
9uL0yhevEKEzbcqlbhpNICHbZSVj4QbmttKgknw2joVV+qvNFkGlU7MoSuyk8E5z9t+nhV77DTzL
O23Oz8S/M6GL7LJRBAYzP6kaJi4uo6qGIGb8u2+bko8A1l1gBGLf5Ypivmqo3dDcmz9Wtz9Po/JH
7PcXrxBCzprPcIlVmtrMaqq4z0b++xDOZ6yctvjl+8ywG5XNiGPSwBORUmVM/2ftmOayUM41fcX8
4WA69332dJHwr/wEJvAF2jrK3Lw4fSqVgatgO2RB8TEz99eQXUZAtMo/o/marefbxzglVVs4d+wh
vXzoIp8u+iUZ5wKciycdWeZ+cAfbnICJh1N1/NiiS7zPmbWx9V9rhM3PLBOTLBRrvUOCPg1PGHGP
+uq9F1HgG+3Sn0mTwvBnJrWvUatOyFlke1YTSPRnbemTGP+5NcDFbLJzva1FyX77EVpn3OVls9YG
apPnV1fmmrMhRJ2HzFT+U6UHqCkYaMsrs/iNSjaN6jFkWRfCAJA0yjOSV9rtV0WWrckEby3fp3fS
g/rFLDuqHMiy4bfXwQ8z/5bWdR0D4H9mZp95ocQuoqkfizHH0AZ1hlU/ZhiSaKFyNKL5gEEIfv4S
J/Ogc0CMU/9dRbUrLB1I/9FMtzmDO2I3IXM8ITPEJaxpCnSIAQkWpE8MuTunOw+ieh6fytqxHrtp
UZTXt55VwUR+9l1mZaxxYY0TzxUrJVMqUD86vm3QTZBTyJeTNFfz3V+UllepTBmLZoQ0tyadFW9s
g2muKiKQOBEqpeuwM7yZ6M5BhDOnmfrowpGKJsx0qC8XK7Hxsr+NQj00pfScI9moQ4lG8ICDoDOq
ij3ng4bnoXGQmd4slqXsVlq2wrGaoxyRXDzWweGCYI0+HZb+xp+xk9o3owfpfIZhxcrxESKZEi4l
QA16Qdxljm+rR1+OWWguqZPPCsxL0puzPoFNP+HcrG95Bea4wFyi7CPTsNgGQksTV3YWbmsl/W1K
LigyFbhDaM5c3Iw06jidECvRJepzrGWEUQe0ujAYDEiHGuyrYEel+1+cf6EK2Ccq7hRnADkR+OCO
CWnbOdMHwFzf5i1D+fR2uWnq95QDH99z/y4O+eBn0CEPg6rQ7q1qKI8K30t0cfpyNb1weB0oFiRv
86vnF9RTWPuAZf4RcN2NH+ttidctAXlr22fKL9gy+/PHDWjLFpT4HZC5MwPNI9Qpipk+jyjBMGRW
lTjYq+KhVDUQyPLA+unnsoFOVpG+Yu80+OiX/CH//DFrLKxyktTLgSwPk3V3m0nAUNejPUsEUFYd
gqGMM/hN7v70QpvtHWtSvfjn1QuhAyYNwUvwt5Uq1R+q5vciCwSEv3l5NQu/LnZlpodIQgglVQaT
r6AsXNBxeZ1h7D+hPKmQqOfExv8a170aoETvfwFfMBcPxGCEP5hfIj0GrpodDyTA57VPVcVbavuL
ILtgzSpdkR2AXxjP2gwTeOfvLCOqZn2yVv6qQXd1YY7nlWYkBxd2iwcgXIniNa3+sM0iFqYD6r9n
c+oPAv8YwgSbbSStPTScVPsCRNY1B6Gm60OTsf4pssl95cLx+o2MialTaUMH9RUpIAu2RUYLx4BU
35nJpRdx66H9p8v7t1HbkqdSrILZg7qHVlBxo/R/ijU3RKBBSnvzHOln+NkUnlwEsGc8+mCmk86v
DUhW9ISQ+UnUdy3pbcVl4mACU9gPCcWyXm23gv3e5mMrJ6XhULQp+w6FhsqRmHI1vUyYtPzY6826
N+C0YP70Fz7mdtXg1an/o+KQioN8Z+l+/oyy0nf/VqJFDnm7V1cYjXPrBJs0mMPAb9YgGok3z5V8
P9eJOY1RAZ609yaTX2qC7qkKBhltc8GPsSToxyQZjPNmQGEYu5SZnpAPViQmgHVXwYpf5paZUv12
bCF2JjYHEBwTxRHlQaFdh2o2adem7cphbg0v/1eyEsHso46XtfWJYGo6JG0Gxz8Rp/fHqsm/mFqI
F37yLgU7rnW3zC/WkU6EmTk1KciqpTlY2Z2Bi4kjZPDlNDdiJkAZvyXYRMjkcE6xLEqbnG2QNYTl
WA1q9VuMpI2v+/3U1YaoSZcmmn0nhMiwrWcCfrutbcSP9ueNZ2ZRFSag92TekXSEyfDXx0le/sm9
bL7n33sAwFr3r6Ycr4cQ1p8EuOryhdz3pIR3cg+sdTSfNG9mOy4R5PSl8FZ5iwtDILlDiWVTqHLG
j6wb5rcboo7boZNOToHj773U82P6IAfcOf3oVlMxR+eU4IOZy5fte2eO9IIzUjNdBiHZjvADasB0
3nMUP+lcASo7kOzP46CFFU6Jrc+DMq2Up5EW88mCOgN8t47yxhdKUbazMXiqlZMlgxIgPVMgqmWs
+es8+xl9i9hpENRG9bQ4cIWX7gL8hUlinxXXquL222vt/iDTCQB1vdtlvQr+gyGYwAmBewJXEaWc
EB2XjGbvI5ONsdZ/XYPWgROblkFb1e8R6k4VIKL8A3hUEPVtKxa+VDUrqPzTbxTpr3LHJxlREA7t
QYkmmM7AyYGAZhDaJRVcU//WndoKLlsnbTaqYbbJ3c7CyxExxiFcgOHegvUgK4xNnGXMoCd/I52E
fbmhyv1WSCRShcAokMSmeqNDowYJFQnHij770i80B7OygEXfmK3lFSD2PrZiAaZBgAHfJXvhzsuM
ZKfpxzvKAF9q5Qq+FoubWo6oyWzXXFEX1wcPJjkBjgVcdFtl13+nY/VLcm7bMGUumroHa5nIr1VL
3WlVszvR3pkiXt2uEK3jE5dFRZQKuc6k7iHr/8XKTjeq9f3LFl6/dvMn8SaoiMVtL/7YZtQJ/ccW
hq9JPJmAIL3zWeBRiAqubPKwsJljJ8CkS0Zyr41eyaKXKLLK45K0r8rsmZRGuMxLTCcjCI7J175L
/8JaVrR2aX1mZAgWNPHpP/j6ETBNl+QhI+UgL1YA4x2soM75z9Cw4Q/Jko1ndAoac9gZyeVrzmF4
ha3TEy/7WCmnQUwP+qImGpYP7YihdXMJIneTa/2KpxiG+C1jeweTmCt9llQpU1wVF4y+jPL9mnZW
llMhrRfJLT6N/uoFnyt3ZIuKPCSgxlbsCpd5phWk6sV9L06stMp1YOVMER3wYQRseDjhhkswcyNn
hnUjfeHsTPqL5kImSc82kvMMoq082/0KF0Pzc+du4WLld+iUHKWHz2cSNyoHf/TX5f2ZXkVBjvnE
OF/9l+UXhbpvABQbIkSadhSZf4c+U6nBab6Un0yYW5RSxipw5zGw28+nmjQoZA6bmXp1tUTRZRsK
uwffMENFd11Gsm/ZGCmDgBAG+qYHXa5mhZzBbbfJ/IyrU6fM4IYSRGMB7ua0Pjb7L+l/FVG/Kuf3
6f4FOs/rIgu/65g24ydWUA0UAkJarsA1XqmvFy9SWnYYKlcUyAWOHavz/QSZIPTeOoBFRyap9siX
F5V8/Y5gh41t8zRaRrrgnC7fzzYE0fmmjMrXCySUR4prsS9eAq33IBF3gVj5SXNbta4zmBUfIOpT
p8MxDO6FhbVQRYO8eB2BoaVPMeibqbKpO77n9jb5decNEH2sP2opodq8bZidvyVnlvOztAWMYcYy
RZ5/LGJpYBKz8WAJGBu6IJf2GBS7/AH+3Lc//bHKI/FXjFCs3gGPyHe0O1WvestegGlUy8eN0T/j
RI53V6q6bBPrGG4K5dW5aWQtO9qc22hlq4Fv7Rda52PKJG6ETfDyaiY1C4hFbYIa2PmxlbLxaYAL
ddBBAjly4NCumu7uWDtXy3Wl4xKuh4WUKCHoDK1PxFAGIU+/jYAyYg6p5krC06czyNQYnrO3GrE7
LzsH6KagGmqHFCOm1CX+Kvsf/Xz+WM0Yj4jcLmV3p7H4kSrEEs9DupQeDPo5jxVqIH6k5BtT8cOy
JHsNfTZgQUOAMjPWbiqjDrH0wSNDTWlp/tdPj3LYhbi76WyC0NCQUfkZsJdJKdNF7AWKelKpQgYN
n0pB80kMXPpm4ov2YtekS3nMfvyhK/qLUOCLp8iFXYGs2PM8nG8jKCcY49guNK+9o33Yd3izxYs9
KB0z5wX2uaYvmNeMWIYl9JexPh22KaoeMHdf612/fxb0OLQta4fAcaNd2eD81eK/KfFKZRzReOMt
5SSDKT372SzI8qppzMZCo85CTtDsnpiY+WPWEkGVWzOszW755+XUZTJWnfZP2ogWwrKYo1ctGag4
Bv/CrOsmROYAJ4ifGbLLt/tuP4Ok0J/MiEBLIygJt/c3XAXyWET2EcDGF0+vwQuHUtbP5IdgD5CG
i3h3RelnInSw1PNf8B7t+hS98qeOQV+LbyDxL+o1n0D6aXrw3ntqis7ZRQX47Hn0ywy9u8i/smcQ
OhaLh2kVO1++0dQDDuCqS+pa4396vv9LTtMARpgzTbFOJ85lo2xhtciVizWEK2WhVUGh+U8MWbRB
Enj1jsqkIy4NduNhW6RKUzx80149D+1ThdkDi6HdBEIKNVakdTkbxrORfR28PQfSinf1wIiIRp3Q
T5WpvUqK+8eG58104iGn43EaVKR1s/V3HDac0JjKQ0tV3XNg4Bm817BuHrPzmfIsHxtbfdZ46cSw
PT4MtYISNVI14C0ro0Hpg+Fcgb0apw2mPJyeatz9Pnd7JusaEjMuIQ0YHqIDNtm6YQ3SYb2iKsc0
MVZflaVn/vOHMePsmzdkXgJ6QtuUCOHiuQ3s/nzJTUYbphI0QzmXIxYW32sRfpVa5UYAfkrpk+sO
yZhUAlSP562EgBgOeb/qBSMyU7DN8l/dTzdT9y3VWN+KzOHJf/JoK7TVDFz/VbZwQRucTAu7OPs/
kHSdrNoIXlitykBA2QNnbhKUpfNlzbBOL2OPpctuTaCSPfIeQ8qSCM63QgcRCBMgNmk66r4zHBmg
4G4OLYzf7r/pL9s8Pl1Nf4rXNMXVobBl3ylCPdznTNjqEkGsN41cA55r0DxzrLS7lHvaqOFsLQh+
Jq/mLX3fKrl+CEXCGULUA+iOWCSFSGUtA3UY86zqyOsnNoZXatESpz14gpBmOFJ98/RTqQb6SZ/Q
AmWF2jUfTf1ITg4x0yu02gSTbOs2iAEGEiuaxvGl9217wIH/u+eYxTE9dxshIfza2UhMM/5AW6OS
tnraw8lVisbGa5gHtLOOYAINN+BLaWRJzuBsc6+RRmUK5FXQKhNQBiJCSCwuk3R+Y463lASuliCC
0vI+hXoRNNN5KaThKK88aO4e8yZ5+2428TOB86y3XsjykmZMdcnBT0xINOG68bLgsXKRu5L7RpO9
x+OTptxDBUrYz1U/Wp3CcmZkxjfNK48wyt15rrYGcHeWMu/4LRKraThvnoD3eGOwAPtNSJtxyoD0
FcwZb9c6IpAiLuvV2ASDMNEfuELO7Ut4efS1jm2cLZWzrSvUyIYZAYyI8aYCG5fdRZA41f96L7dS
O6obNedCKdy61QAQMgohSgz7LcbFPqQzvQ1ZAkOdgLQpQQpmup3aIYAl5GSyu70Uwab36HQdtI61
hi4/jAkyH0Mo3ZhSaCKcpVFm7flOaBc0nZQrD2u+aNKGKU0AUeRW+INyjbHUVrPn3g80OaGNsbKL
g574fG3J1fpBApBQwaDm7navYchnGNjoMGV8dcoQzi1Bo+/9Fwbq+ASirBW9C09/DNGjlU6/QSGo
4P+aLtQ0GOrPdNo+414zgSHTKiEqwC7kb0KW+k20UjJBLtGo2LK+zmmGe7/EA0Do67yPc3zeWNlr
pWce0YG+HLWcodiYKIaqpZvS+VyuNZsCeWo40VTps7/ltghff4/mgHUrtMPWP0pPu+BgM2eAYM24
b8fc+RLGXNPKl3RRKlpedc20UpEDc4CCZlDjB0IWfY+dBvzgN0uUlqkpANOfHfuADrQt5Kid8TXD
60OWgCCKcl3y9V8J4q27XWy5LHbkzn7cgtWjySdYnSr7hm7UZPbKEaI9zdJu4ieQoRNOKB9P4E70
gsm4RmnA203EhrpsPJLYlxEsUjcy8qQQVpfXntwMqae8Exe9eW69wPk1qoUX5rPhcziHUQpg+pYV
95gwfzwjHCP3/72nBEG0DOoQIEmTaiUm9ZqFiiqs4XYDSR9cGh4rTPAoyypbvy3jMk9iALEsdUCX
LwXgK9DM004V1GXQlUt76XSIaTWWd17ONB7n5D1lFWNMoFhApegYtdM/VzOd4NkcUx4UGIUB6Arz
IzaKlotSq1FNop0LGG/YhNImh7bZtyLVG/nWAueusNUd5bvRDujDqNOFJyyxhoq39XcRmSpdycP8
M4Kyv2rYur0Pj9qV2gdsClaGPIdvUTqjeV1j2K/BjtjOV3+O9vaSJccZJptxjjHh4pp0QFkxF8Ux
nSezqtEKV4YvOlAfjL9hlsiY3V96Lf6xfudxFVj3rnzDklp5/aDoDQIeCG3SPShm4M+cz1BcslS9
8mO4Bv3AW9Q3S7KH/eKaN5r8sNUHTuChjaVRP4k+/4xRdffx8KgLdLOixVww50cStGMscpYqIS6f
9s8Hq5dsrhNAP16+Lywr+0lxfJGxy3bbOcUKzDOMAAQid7RXAqNnChsfiTJsHNQIRKkNqjMx8gpq
h8lBPyR6CbjLqk53S5PIyUtfh4GfE71SDRllXm4FLl3z40dKurkZV9hpS2cKSXFPtxRKBexjlhVR
JnYV/9t8HlE2tVQNonzyzKPHUZ59xvwOMukdfVoMFMgExEDRrZAEeH+vA4f34uFRp7EH1vyZE1n+
RFxGJIyi290vW2aLL5aYaz174lwl4ELvhDV36gqVqa9DVhX3FOkK3dFsqCzt4yKjmMbDQgZwHLZk
jIpLjzIgVCMSdIvCwR/JGKpjU45TkR/hyica3okyvDvBNs1xQtYuZlVHU5xevUOyrhwJY39cP6NV
13KD21MAev4PeuDAmdBH32mmqjByQpkN0dP0xAjJBh41FNjSRIJ3qfMI+1fq9Qqr8ybjmGL6xRoI
Iybkscxt/YAYTsiHJ7ZXrLkbpp1rla2hhvoOKO/ogOTrvQg1JcoUEb0qAn7MQyLDiGzWVuhi34Nz
oDfbDYgl55zTSECFZQhxrFrZ3QnUD3UgGpB/ltg4H8oJe00RUrwbe3p8J+IkiIbnc2cT17vo6QRf
2/6jEfmQlVLae3TptDpW4qyS129RGVhV9Y0Si9NpgyRqJkDm3NwDGBJWfk1jhAQGqyITmrYA0GAS
p3APxzkgttMGjrfucvvEizgwEgRCD3VHiCAk3BtKltWjfQBp0lGAITrbigSZCelJwcZnhlihfjsL
zfBCIoQLxTWu/EPZbWbzKjrikJw9kC5zfqMuJs4pg5cXxjjNTafegy79NXvzq7i4FqD8VcbkBenI
OS9AGpUPdoD9vCN24CXnj4ULZxP/8Cb+OXqa6Y3WvdKD6PwVPuY8YKV19p4GlleW0n3/cFiVE6P1
PG6semo2X7UgX4UgPbVCk2Q2t1Y9fx163wHs+bO157PC59y13Xjhnm7yx60i+n5qJUmYNT2EKKST
Gy1N7pvk2+rll/3+jUGaQCKaa4KChUp1+Aw0cusrnVMo9wypeKbZ1Aqvc7AcMJp0+7XBWRNlDvfA
OYWTymuLOPiLsm6p+VZpkH47ZC6SOsWU56Y/Kb6Q+nfkVMG/ddvgmmPprT//ePgqGyNTnWqS10Qe
pAtr2p+rwaIGx4h9JvizSIfm/nlpXNcl57T+IWOOoumBXL1RaXDrL2PNpk2aVQ6jv7x9q3qOPZnI
VtOoxXyIHXOMhWA9DGYqi4yPHw+ey72ln/IfFDRgbH2mCk5FOmTYP4KfdarOSYZH4CMci/vNk/Fp
//fJ+IinOFTr19MfBm+SiAW5DEk/a2kE1Fuf7XPcxxbmt0HqqdRQQDdTRVMcytItSnck4UkZjL/D
MFQEzMAj9a4lZLJVKTbuEFWR1T75zdVXpc3sVQDk0+6Bv48ciz/D8DfSt1yytylzy4SW4WCzqILI
U4EFdSgrUnyfCiNOKud1KThcdnR4lOcyrKXbDet6gzadnXMEvB9Xpz6bNIa8VkttzhkPo3wQ0kBG
qabPqqlg/2/EEd9be2zLFEAxdkC6SkhJuwSDvo2osm81n2Vg8bqDBW+G566JMBHxKXp1wFY/Mwof
oS0MTpf0WZ9xNR/pEu0/29Foe2LFFDhojruCCIAjecAKcvRR5fPxKzW6/Vy5IOOe3tqjl3tjWYyW
KiwKo8q6OP/UQUNl94jYjIffzYQUXLatsssCgsKrACOc55E/R+4I0qXRK8Z91fMOB9ykjS9FSKn9
D59KdN5kTAtsMtb8yNXRt1x0IEl1D1O30wYfJ491cvQIXnJjDpUmyr6bMMXOZattL6HlsnpkkGPe
OczCFOGdyklvT/qD4ujuuqG2n+zVtC+FqQFF2dxNBz2xlDrmWaZ1x2F9VUa4ur6tesCujfXt1EBE
8AC8i4H+k900OHMq5Y2uFrWGR7pFo1RH0fe999DZkUofCO+QRANs1pJSdT6J/qtN3x7uXi/JyIXs
WVx9f/H8EaSjuwKq32XnJDis0Bq4lyw24GDkYfP0VUlPYb4hGfS/AyhUT8UiV/lmuWGYwegl81hL
+Wa3quW70+UAK5VOCrsasYkukKucgNSgEX0s9ytXSzMvpD5Gq8p7iWzkM7OHZkvk27sqtPsxHVXb
upW5i0bYRlreHwumPxBMFbYSXuaUovgvZlPXIm80iD1NtqOcj2fi/bsgl9OmDutJOSFbGZESXDG3
N8HhlfYA+m7riVghkyXmXTvS10VhoTq1O8DCq25ZyFthByxSK9wFQ9GPaH1N1eifgW4n8ad6oExW
y8sCTuLYFoEHrB0Ui+lLFy4KkR6tlynm1fQzg0NmJbrjEehIRNQBS5Y0cw7UMQfDTHB77aQITgD6
mvpnmiDwQxfOeskDtubfcqJOrh/PA0JOc2W/TdlnHr7xmI59woEaDTyvwksbUxNo46OAyGF99AXK
Ac9WsL4Z1YpJdA03YSPxnYfp6xxIRgmZ05YQDf4YTttqqJnEZEV0oi3PYdSDX/RqANBesuHD8khJ
YZnvyGwmGyOZxe/3C7cu3wquPJyj6KzH/dF1qn7ZsFnwvAk2mOGaHFYqTWMIt9lLuticn2CmaSEm
8pYjPRCnJ6ukddb4vzOITeFd50+/OKGq7tOaDh7gFpgqbaMjACjyTEGSsYMkAC34nujb1AL1U+sS
xU20f4TVrLeA1TK3VpHlAu5qwP6tV5oBkh0Jm7quQWzjjr4HXhFADe52p2rfSEqYyti/qtWyWX3c
vWNxG4HwezBOJ19AWdvRl5PuYpikLiC6q3HvKrGnh/UtUxukjDxZQm7NTdq9TCF/eWJ15cjY0ew2
s+Ltm6VSJZ4tRgcv8zaIp8BtUw3W/vcR1jpGpDW1Uz52BajRKllXMsCc547SszYsmEsifS44nd/z
qFdGVqf65/CTdvL2irURnMnascBDVVK/NRS/c1uVgzf5M036IGIFGsYItKQpumnHIejdjOTaKsAJ
vL0Ilg6jeq+xhk4GAgl9zMUjrY5rWb93aw2PjwkEg/f33dvICixUoLmwuPzYuxW1I55ljb6BQFmx
dR03sPpRT0sboMTkp7sESpDycAS1/Gk0yXBpFRjjErWev3BspKHjw8bpsncdOQ84Q3/y7fH9t5mu
dK9Oeod5iGKeDUD8I6Tryzs0HBDa2mYiN6iBKAX3QkEBLUZuEXY+uZXveSSsGaVNCaCfnX9fWY9i
eryixRtD4e00OThXD/B6yIKPRuX7WW9TynUAemdkdz9dr+oKjMtYdcvzAKCi7QOCLy3MmTkiA/Fi
8caCPKn1sy9um5eof//aVqAoWie/ozpzquBI4sTSm8fGVm8nb+jngCQuBmfNOGDm3z0leNAg12X7
s6ztRKYmmFL2mB2LOwGcZkGM2e4pIr3oZLrsgdx/2FfzllfrAwKKGAkcN2zogkB/EU3qilQhuWwe
phcQQJAvmF0LIGbfz/tmqKqWxqnqR/OZERA/Oz0hzK9WOw7ArNcGIjpuqbct+/aYup++7Xt6y6kz
Jf/aFtjKq2ukTytr0fvz7MpsC4Q2rbb7ctSV4UOr5KEppPJOrVpvt42brMUIdbLmBoCNTeg7508L
U1S/eUiRVbuD5HYn3bOpVZkepPrfJV2KxgI2A5L93vVjjinBn1yOjdGrln3/PYVxzr3R6novbm5q
MUV+GT98xrrobC4cevCbRGhRJlLWyR1k93RcFOtlQ4jIiixzJyO341OAS9pNWIDhDBmlWOsjEgYG
tQ0hxTHyi3KFIVJGda09nevtu0Gnd56qWUSr+1Ib5fvd+Mvf1gbVNGUeJaTNJP9FjsW72ezvgTwl
k52O/dg3SZJyGJYWSPnurzDVrRxX2v/H00kUeX/KHSNOgNIRnxrEZy0neAEZQ1qaHA6qKjixkImC
J06GKCuV4Q4/KDgZIC1asRYC59HYdjc+qod2r48h6S5wyJ9ca0BNHsz4QRQRzU3uhYqybv3/70IA
VfBt2Mgy97N2/I84Mm4Fv7zq5kluwi1yTSTY4/ClwRMnaiZd7zD1TYZ6gjbeffWvXqcmofQ4H2m5
8yZe1BLoKLu20bDKE8/WwPd/86ByS/BfF4agFSZ12bHN+NSVzqf85ha+sOv95SlajfV7htMQqgCb
5esjWtzxaSLZtPmlxaEgcMXXu2Kw0ilbe+sbT4XQEYgI2yVuegs3Xtbz3yDMoyFueC2ms2Yu/1fa
olYeUk1eY9+dA1lMwNUKs7W1i1K4Ts1JzwXhuZx2P6jlvDh/CZOvlLFGUa8W/kkKkX10azGd/y73
fp2RE9o0j9Fimgk/teuY/EGFIwMBNarBDhQb7/I9mD0Vr8W6HON1Np3j5HzJ+Hynko41+s6a1sy5
G2OE+M5zPyOKzjG1LHb9u9lNJF6U+WT02HjfMGDXJpTWtuZ2qej3uc2pxQ3IxqCBLXCYJLsXMdbV
yWvJxvEj9iyEkcOGVtJZ8Wog6FKoQ7jnPgtCYnna6BDjtmmcn/fmUtdpqH9qXoS8Tgq4v+pSfTKB
4ClEoMRkNt5mU9xNbJ6aWrAztKDvkUq9BxjzMUl3VSICEC6SrAAbJBVEPzw2Uavlj6mSalhBkvOQ
C7xU3hzp6wOTqxNErbX0jTQugO6qOhf5MFuttMYbSha59yUUlErrSvKjSks36Kpl0pBqUzP1jLh8
DAspj897Ahjz2zOJ0+c/Gqn5OuTLWl4Ty3jIG0WXkqrjxPW9mXjeCKUSxv1uSFruZdByeI3PgsPN
2DPz8uqUo839xG6/+CtoLQtVBh7yhQOcIJUi9RRrK6w4KpVjH2Dw3JYy3OTrvm8CHNM7ZHc8heqy
VM5drUCTabHDFQrd9mMfB/KaFIw2klCBh/I5WUP4rKXQcvZnD43DAujr8vjupxWBbPNENWU/z3YT
u1XTjqxM0HuUUMy2b7blax+vnwTx9aV5sFwFyhjZNtCuUbxtDvjlq5VwiJaqzh2bUgOxTdGWM4jH
ryawP45hcvhl7e1h9ze8m153Nxay+pcwSwWGYDNgR/SLDUuRbyypi9zbQBC09ssvCBZKRrFjNUeR
PtT1xUA5mgFedxCvbUPOEtvsDdGNLSDa2r9vFCKCchqjK42BDRBxmkLPkSGsnX/uJhyx5Q5eVoui
kd19m3ua0895jpy18ktu/jwYGSdO5uf1MpGaZtooHx0Qw+S+NgpciIf/6dE5wiaIq/d62KjLCPTw
IP7ubVVldV2Q4OTG7bLjb7jUFZ0Flbr6xXx5ut5HtYIUA3w5jerjiYLlPrENRVc/xXibTuV7wg6t
eh8jykfETyhq1aW1g4miLS2D7ud4L+Tmz8nrte/ASjAROJ9X4mLRDeFmTCxxipBkJupWQumiPY7X
MnS3cU3UL9um8drtTXE6XYQANz/CfU1fqiVDQD1KPXVAhzP/7ljc5126Nmp30kpSzRBYPMTYGxRP
rpqsLTkxDZGGESdIw7YcOfn++f8haFETCmRyRIosqbs8aF0C1VRtl8QEn5NBXsv2v812APIRYXOf
FmdZGQVUUVzsq5PONZm0pXmK9dftTi32+KI/ffH1VtuHCYI171CW3RvhvoyF1v8PxQVop1MUncD6
PSZvoQP4JReyKY+tv7AInMk1DUQQgv/RKMGezKt1Ujee6zEwjncpLPyGYo7wPjcniAJyBDVcjpJ3
hnsv+5a9Tg7KAmdmSsJ87cuoD5NROcrwIRv4N+z6KaUj8YQm1H8MUJ4LvaNfW2jMhcoxTECJHRpb
FCp7ingAb8gac5GRs+5/srncsJnPOR70+8JNJ7sNpcaE5KxuUgOmWwMpeeknXIgLHeNBGcrloeGi
rq6l4DXRGmijQbmSMVi75m+d3rS528VogUGl0Ddos8/3r6GmODGLSv+7jyGtbM7Ow8JamqjMuPVn
OOKtitxxZlw+OrobK/RQHXaa2Wv3EhbEHJJdauWAPzo6G7896dZ+Q/LRFExau4A+5PZXDrYiwN+x
xc/HjbEtdFqzx9r4Oe2mX7meNEuiO661gDd+SjblXRD7pbtjfLZ/A/i2U34qC6NR54cn7DyvO2pA
ojmYcekBjsyp4+cBvXsqqdxXYEBWOUQbxXOqnisixcrTfvY2xoYkiNnD9dNR7mC+1TL2HRra0QsI
o03FjMgsp98KKhYsW4lN0ks4rtd5QrqHxTO2ZRb+h/pIUs2SgErJzUlJyyOAuyGE3yTvPQJDXZO+
dzEajdJ8TK8C8JQh4mb48j4hbchQ6DyyEogXTtsvREvuSxGbMxmMaM/oZhfX8bJgelHmamrytss5
B7vn6KN4pcv/Pkvqj1k1JLnhFHLH4i0r/PLoWgHSrrkUKy2A4bAWIKBbRUJ6TBqjxuf6eFqAuWqE
rhm8z3pwd6GLcXd4yZueboUCxbkssyqvYuC9ClrUFse1FdRSDa6Beund8n7JP4J+R2n2SquSTcGw
XyZrsdHFQpMGX91/n+3GlbwaN6jP2kXAw/QBHRgJ03jB3NmyuAK6EJHWhQ2kWX2c4mNXT6YlzP/U
cuWZUuTca5Qht8fUM2XV4jEKuBHYyuJHD/ttEKdzyl7JPhymVNcKztVMuEp2ySZD0lxbkOya95aU
eTir2sqNWvHQgLk7UQYTCyDgjl0EHTtht4SmGRMiW/bDHMm1cBkHc/2iL3s18z2G5Vlw54kKuO8z
iZKKGhte63yo9OiAoayP4uDj3UT/LX84kD4yprFmIMwm3T+3nZv9Hfkq+8GMWSFnktiT3jqE4018
KYzlSeJEj3vZfoUz3X1UQRabsDo3z8t3vdMVnU53/Sd1Fw10cchsIdAIrjggcAzCTp/ri1VaQYtW
MGsoEBNmppQ/cwU+9R0AdcXB9nB6QnFHO5E4mrRx2HdPJn9BgO5XZCulTj9HTQuVuGM4tYNKk+Dw
cE6cd+Q/KnYdSrVklcCldmegOinMci8tRUynmj9WwFJhYFc4a4VP3LAH/3o6vddmpyeLPbV3yQ1K
kIEAbzl8PTsGgrp//rIAHh7XVOAMAcd9QJswOHiooi5RdJ5KTNQSXRkrymdWYVPHxyoWs+jtvSEF
XY0UHX6msWacHp+uIWHjtgwlb9spCvauV+TW2FJqLhiwA1n6zj0FviiyjCzg/ZCV+y0Tdg+01uC6
L04XFoTA6b8ZGgiYD6lz5d01ymtANuJDvY0PsihfIWQ3fjoGvTEbBpZI5HgJwKSH7iq1zVTiN4M6
XhbYiHeB6mfNNJ9SpHXqLA+uFp03yrMa0stdYIk5uKZ5Em9DupTozhqgDwYuit4J2t15TDZiNtiU
zXkXglqffhzba+zZk/BI20+ByJ4IUBjCMWRPuy+zOKimStAdeKV7QYbAPuPDpjfO2cpe3Am6+KK8
DA+2VsA8TowWsvzimrQSjNHtj0CUk2P/i839ImoUEwifi7pHFDVZZvOjPpyy00GvVNH9eRUifkTc
B+dOWIQgJFW69WsxEzKpwI9oc01MRsx+GGemNOaYNXS8K5O4yKZ39s4sB7Qy8LnvGA6CbrMMMne3
ou351Sxxx6M3hmXYPRmK2ZIxagLo6bMJ799foYIgtn4P2nxvmBe9oqKDUHQ58HLC1qpUgjXpHtVm
dl64/NkN/ELSkgGdKl30MXUNVP9BcfUgEPGB61JSiG9zQKjRkUymVar86+Disiq5IwYb/l6a2AlK
dgwpdgGYI4iKFwVWLggkwjhu20XSR4YElpN+9ohhtBoQFWVR4cT3lIkW+qlHVGS5uEIASXZcS+xs
Pyrkl+7y38iPpHW/g6EG7uMCAfH1C2vZnD0IzFoZn4Xt0KljsuGght8dYKvkYOXwFGuZkjTuS9DL
A15W0/KlrlpJQs9C0+avZk48asRZXjO1DmQH2GmkdNpqvKAy5JcYmA7EV5EIdxOgAuib7vXswyxy
mH7RH6Tt3i4l4c6w5mcrPMaGWPHVb0uvI8HwOUQZ/MQCg0jZrnEsOCVSTaBOIC1Go4mzlITo0eAS
OP2DxMzreMqjJNGcWGkJ9lNmgyMgI+6AYubgBtxpNPyIabBbTAzcOZ8SfXjXfiaRndeGr9NMroWw
Z+aVeQDGtmteDv8IgqeA19793IQQW6WynT+NgU1jQF8a7oqMZVZ+77wC4PaHH9fSeGdaanFZARuw
zV+6kqcqft8QlfBFN4021LuC1U2WME5LxTlwA6mN7mtd3wzLS74tOaFXdaNZiaD7OtrXrwlDn6Uq
lA4/Ib2us/U67t66SPY/89QrxPmcshdBl888xgb/dFMwCSomjcQ0hFDTWaiqa2dW2DMYknwH0ZYE
oyjDRg6ZRQA+SHpfG2SR7gyPnNJO7/EfiB+sDD5/GPkNsdDJltlXkV/CPs+6ZceNwGhw6daFsf2n
MXIqSQ851PPw4qgt9iuLrCozVU4iUV4TK/rfWlMi//0VoYJk1KD1PKnE2IT/H5cASJV+/nijl90b
N0ECBu9ghWGLy5owNCUhbazBNp2ouy69EP7yrazXuwk1XU4m7zTHDt1VOaMXkFU9B9tqKBWrXaYu
xfoX0wjdAVEXYbOllLzJblzTUo6hlLUUeEMBoNn9mRaNN4oHUXKiXLAwS6EZixBuCU3tshGhkIWC
uKNX7oyFCSrOX7Odm3mjG0BX1dr3ORG1/o8pBY3fcZSjwWfONXhiRvFcZOFNWK+2MfbaXg8lu8dI
hP3tSgniv4troy3KWtUFb74kDtmhfK8v3//Zg167G/s1HWKz1EpbNnIYDONBas5RZ5ScOqARfomz
BJcdRuXFJSpME0MfuAw3w5nz01SXy7m/ngu36AYeXSCZesIrzR2DD7yOXweReDXq1d3q64Nrjxwz
+kVPIJ+AUd1bRTAkwT3V8FIsuGimefSEwDKDih/rHkuy/EoOiWd5NUyrJuQKW1pyMgk8iHI6IiIt
vniKLLxrmFSyD+gpxz5WTM7Xa80kDkXiakWq1OUZmg0RT5vxnYJGwVUJkj5UoKg/B9pg0hGA7Rwo
fbR4B/7uC4AYWWcHaQ7FyPGk0LyT4v7YUdmFcJkim7fP+/ymwUeet+QC52jA6frfP3ZqckoOCPSk
BPOLK54WXKtTUjqUoB/V0khlglU3PqKCYmmIejDdoaSSBCiNaO46DlDnnxWTTuhBPsGm+D+5Onu4
li0LzV+kPTjuDg9pY+chFWVA3D2rm9nmpxq7i2Pi+z/fPMnRYXj4YJO4byUDOMvn/CK6ILUghcQD
VQCu8/pz/gEdjLatJYYPzbXUoE8BzVaMgfjmcJNPMSr2eDDT/Yv2aj+ugj78+9ApEzuMn8+kLcDP
FkHTre13aZHrBUL2XiiO1DTuUvv5RWy0vhGTVbgZlYULTpcIBbwGQ2m0V2oUuL6C2RrKaG0TXG2M
2Zk3dNA/IlQUA/0QZIA87yJva/vpS18Aabd+vqEAcFDn8kdtdENNhXEweSkzA8/mJE3RwknzBpM7
eQjrxHBE4LgSGGTsbPVyhz8UYMtnB7sKTnKFs8k1NgwSvzWW5FAjrwClXLZFYqBXI+acqt3hR7+N
+Je4f6nsitwLk3YsDORzGNLS7pJDGBc00DtBEOiZQxF/rqXt8viCjvYHOxvLlleuWm+wU5Gx4oeJ
Kp13vFrUrpdFjmF0HZEZPJR4JJ2/csc+YLDIYVBVS265xEvwacg0QPZL790C54ig4mhXa5kqULew
NrYqDLF2gBFjBTh+Yxjli+0UbPo00ao/lxTrC9DvHBGRfMI4r8cTAhTUd7y+yu0pZTFv9TRekbhd
WWsJJszG/kL8X2Sw6SCaMDeztrsA77ijiIbsJSgpOrFuR3GrKYQo+UT3NZPrIzGN+XCVZb8mf4zo
yxRPHXRei4Ap0ErK7xPBejok59C/hy6gyWiR7As7CxWIaa4Y98My1eMpPFuQnKWR5ZqAeOJb8QNL
tbLGDPAFglVJPkRym/QtJvJwWv98oPRqcoqG5jl1r+CGVPp4VAxnBXktBIQLOlizAOm3OnTE/wG9
xVgXZRdahh3MeIgLCaI6baV8mGppRung5w8s8ROxFVvu+Kx1Z7bCWpmGxbcg+iz06CZbWYcKnGzq
ubOqe0DlqHl2oX8mGiEUI3S+ueLELQM8HlFEj2kUEzWEgDIniTp83368RXGHmkvARKnckKI8Vkri
xD/fWfI/3lR0aMKYg0QaeR6w3h0fgC1KO6yijHFjOk+I+ttMwSKBVFNPZVqfcO4j9ch54E95STEX
F7oGhyIdsTc2TG0XdaOTbWr/VEfzDqPv9BFxl4vGTOBgKnAyAAewHgP/3jqzZngacNCusyT9W8Fj
lsSPJAskiwNhzPSa/oz4oVI79JtNu64N5sIr93o0+U+vG3vV9rVRf9Gv5LHyh/c4qZrQD17zjKuc
LWBMdoPa/pCuH0VPRmJ75xbKFVsU4K7EWvfd4hFYhpakLPqyJwePLUKAVwQdU2aM9kh6Rw+EHvr5
S3eej/DO55/BM6ixOSQS+PrbQ9SRAWH0AQ5iIRhmKKx8BAkg6pfhvmlAbZ8pSFvoCguwTidkyRs3
Gu13Q2gBBNNjwnicFTjWdIPxzVYUgJFTMgqTwsHuW+MalLtvJBmpmoRkHQnxNgnHfC7b7isFkUUr
+x15xylvvROTmdlbymAKsw6hl3yJ96BOsQUWD4xzbQ5kiCo81YQti2KJI2z7dlMH5oOvg5eMA0zD
Hd/iZfCTPif4CgscTUDpFncXPzWIcZ+FDYBSP4bn554FKbf9fo6mbFkwE20ecb4oWAgFXRluiHHx
/8EOquJ7JARCyEa4HCdMCNuTnsrvrhqA9gtXy2GIyVvz5NbEjCXV/5PFueFxfKVDfkM8hLDT1Eiz
4kH5IlXZQK3U70RoaraTz3kXhvaH4SJNDOY/+STh9sTzyKIDifV9DYLuwec3G8quiGg0o6aGZQeq
etjmCHIsLMtWu8pHxM/B6kY7jYCBCR06CaGzywBFtmUJrI5teH7bae58FmQMN9nJfZfRoDYjYXNh
mTyQ2S1hhpqjiwpOSAv8xm+YFpVbTl8yNFOUm8uYekwMUv7iY49tyEqngJJ3jt5cEcPLW95eY+WJ
s1eccUx6zKqQhPEc7OLNTfuCrn4r+QCCxofMfgLhIHyHo5q72dCcP65Mif3kzIcwYB8nIsamQOPC
WTCnvjTDfYt7031jBlvCvokbnQxJCtlBeJMB0NgULCjNDTM0AQJSp7fCSpSHwXCB/Kea/uao4tdT
TE35i842w1LMDGm4dcarJbH33iH6SAzzhf5wdRfkwu5/q8XeDlxX0fe75oZ6Ziriw+Dw6i9Ve0i8
Y09beeGl/sTCRlHVaXGFU2mAGql3pcAVnqi7MTG9vkE2fbBb91EAR7xD43l4340i6tqeoAFTXK54
tRn8sdXMFwCbFW0VrOgdfNUL2M5De3rikLthYwwNMMvEf++WKzqifT4101Z9kTK9qlsMUZHrecJi
tDS0f0LG/0pEjd8BWrUM9M21STYEPV/0d3XkCPcC480QdFqceoNlSzkNcPV361C9ejPxlIQ+vSyA
Kj4suWeEevA5zi7qv90T3EtRhn/+ZCa9mM+BFWFHo+hNOaxHLQsmg7/q6T0GLRk/aJoL29JVR2zl
O0s3RWx+4+zV0Bpy8y15nRA0d+OTt1ZeeWXl11uwgS6BREJY1B3m/VF1vP9RkuLfnVjtul1+fEvF
R+u9ovW0KfisNyU+E8kyUU6nPzvTeEDWs0OH2FL52QazGGyQdz+DHrGuh9zKBHIc1giz7/13AEFw
/o/X7tutcVaR5WTk6naBSHwJWa9gXBcXLPaA7qcM2J5ozx6surD9DCCcOb8WybLURYtcOW5fvU89
oxlw+d6sIuobqICFBTuu6QRcu2vsFbG2T0CRXIh76ben8QYW0Y/l91PB/92BoAKs7oZB3JOb3BGX
JYKnSngMGsCMFY8oIflwpJGgM3/b9A3iXRpowC8jrZSBBLa1AH0LyUCDc6+uga3eHbzlUITp9kMD
u0D0iagMVsEpfO+dQP0kiE/msUCr75/YzgNUEEEfusHRx0V55i9GtSY8LqcecUxTb6ITpy3ZLoHi
17eOIcoTADB+6kqGyLXvu29ruYdq+RE2Hh562W44UILxv8Xqncig8RuGgVVI5zK9CxaIYLRKJKTO
VUYHUnfl5204dIx84kWtZPOmA1mpw2PZK9A6NLq2wXCp6NWZKQFbzbBkROyrbspbytLb5u75JNHt
1l4SALdz3V+Yxkhj1U4XptlCmgUJG7m2eH4Y0bq/KRXM+oj2OKz33pX6xv6XmSH64mi6AWj6X2VF
ZNOw+KoDlUAu9VBh++blGxavfOmeJWIjwK+V17N9KO0xHGSplFhT9NHy7u9iOJ/Qxr0xefl+kMnI
R9ik9C2OApY+nn5huW8HM3IMgwqwl1BIMVxEy+anTLRA1Uu95e0yZOAENoiZtpsU4IHiOsxhHitU
GkGZH/k8C+SzEng1wOyScpUp1+GqGkIFlEodyJdvgwIEPwkp0ZVH/e/7noGj1r6HpToOu4xbte3Y
TQMSqZNN3q7QYeYnyGAR+7XDgwd8HTsbDaFUzAjUs/18lrbqpylNpdqQlbSDq+r0kM6VpZIAHQs4
W5eYAfBZ+0H26an8bHklFI/jJ/42qWQbJZ/gIk4ir1ikzw8BrZ9ouJCILC5KfSo+6Cl3/I3RnNvP
roDyLKTMcSIx+KI/gDGTlYptpr2gNjRs9CozXYHafLLisV4+o53c0UqIEZKF4gwp60ZU7oBJvV2+
T05prbIRoFNCFcIcstCpSfG3pkpHQOuCO6saaytpD0Le6yfbiKYvkpTDWUruL1jp1lOrzY6+ukTm
pKdQJ7hMJ/hgsh+xUsdUh+e8TjLaj3J4aK8JY+ix1DWLLCck0pcqQXn9TDmrG5irwMuSVhk90UBd
iu3zrOpz7n0mEmcKD9wha1kyZvYC9k/Nl4/xDk2LMkRbn3foDM7unoFQxrLq5kpC9Yoydi31N9tV
j+dxQf6RmrGXEatpp5ihfWs+cnR5mnwZzQDq8Ims08qlOGSG/AmMo8mNKdiMmTa9u+sMCjXpqpoq
JdPeOdvi3fGmLjwsIYL9iMaA3ohWYsF2IU5Lq5fG3FaWaJG1AmgZHtmR0BsRV8dw70MNyaZW8oDj
XNw0yiPRwshtBW8L3Csn82oaRSlSViAaZBkVH3C8k/vHGfr6NQwcbzue5pORfjokTNa6soUsPIwu
lCAzUE9exLKUi64JdnAHguAuhWfrY8gwngjg7PCUjDtEoN8zbQeRXc/CagI5YpCFTlE5tdNQ0eau
cuk8E/Ry+j8oreYOKf1STqHcmxY+LleGTo4DpNpjyrPTmFqD86eAjIxOisdCt61SJEGOq/xLjMg0
4NN7zXiRV62kcJkrUIOyWp1zexuomMv+hR0o9+T2u2oJxwuYJOm6IbYWGujXAx1TwuhSqq2GCJ4z
zbqsX7CWiCmSL9rSByLrhwAUXqH2/efqHymWC4+ZRVSGhl4Zk0siebW5Maar4fvUN+2IzN1Wan98
NDwcroYOtgQYTlaR5fshu39WPDYFkGKhRK6ubSNzZrX59so+2+VmCW0TRtnn6SUYFwGYC9W9PllH
ZZedV8t2lzM+SXzE2mfaxt16TU8+gszrT/RsZXSdt1h68p5XMwB+XZtpijVv5PJTogZM52iKAR0S
LvE+ukPrH2IspK7fvu/YSRj96Rx747srJTvfWaCvGCLHTdzaDG6BT5dYIebxTuzTMFNNJ+UFAiYa
m8RRc3BU/s4SXaAoBhH1BL5Hl4iGzWHN+0/Svx/ioSOthzHxMXHgrnyWKvZhGme9Had75ARbMqj0
wwmBFow0FsJg9EbmeyQ3/Uj84mqVyhSCn0cjE1xdFqnxiLomwVvyxJ0GrHAIsgxBihiwC3sMjGL+
z+gQ1b46/Co/99CTrpVSGKp36iV7aOCTjH7SLpYddyT4RR3VSNUXmXWhezq1DOcXZ6jFqViA8j7W
T2bfSCXUvG71xjn/J7EoCIm5VOfiZ/mVXscJDJBtWj3xTTsj08VvaQvPSdOlYOgIpVm6ZKeC7JsI
W7fCoy0FTu8tAhmO9nDb3zOLtFk93V8wk0XhZ3LbbrO2M5d5oZuwruYjj0oobQ5DzEzxsb6yhvfN
h+tfO6vq9Qg1MXzduCuPgMo2GbtdD1s3jdrFMQNGmd5NVH6Z9D3m9+hGQx4Fda1xLadEq80XUdbo
4+MvOS8PEWrZDEIcPB22Q1Y2FUPBgn+BkPdJqGzbQrujxpkTWDgcVlKGo/g3JnBIK1PfATiYGuqO
HwzSjhcv5sXbEf1SEqrW+XTnMNM3wM+XIi7sqGId9hqTKSQ+iVEqF2J3KpSSwBCcGoqlMw0mJCh7
Hzjg9s4RYAvgfvMQBQtpLjh2Gtj8si7c+bJrw0e3tG1giF7ovvLzbXMRls5H1jPjua6egR6nRcdJ
RsFDCmoJ52/rBYElNq2R7dhwl7woA3cMhVBqKHX+FqeVWmwin5xlkx1v+f/o6gSrMimxCALhnyT5
4FsO4rpGXg+In0TDFodr0RkVxTerWr7G3LMzHoq1AwWL7Srl1FwIE+tKljiDpRy8cvDiXI2/2Zy2
4D3lPi69+z0MM9bP5GeNPzOw7/qUkvVs+VwVmlSkV/2kXiSIXAvP623dpCoF/ZDwwOcXuIJRAT75
WzHLshOtFHwxG2jC/CkSLI439Pi0YUtnJHNzv1hPXPro3cPPvHlu0wfHSx/DnPDPCzVN3WmmuxTX
iEgF5o6qQt13VHVseiJVR6t3qL8sycgcFLQgeoP6RDIXLXnYcFCk60GOJP9cBzhJ3IAooNruC7Lp
7zCjg9lYcJ4PyWGBMCo9rjsrENS/JLpOXzFpb2agnSgKH8s5qnVCHy5TNOndp27BnE7Vqyx2C5+n
LuOX18RUm6INrBy1ZIueGbo7H0zTiBANf9uqcAKgHkZQAHhnrxeAsQ1oYWgwNmyulnXpALv5w/OR
parccahdQGJzhZ9QMbijnDrTEcI/IipQWDvsTJ/QWHqztHEpsYByn/mTJBcbm5En1uHmv/SByhIJ
TsRMG2+ijx3WPSZZlFEaqi9U+p1S+vpEJCH+ko1YkfZywDqSXVbsQGe807slLXtkbzBD7TMl6SUp
pT+qlM3aYlXhxgad31Aobwq05OFwKNmKlOQ7mJk78Yl/6tHI8JI+u31td7KiD+E9dfmVioLh3tqE
FDor4EGaEUaET3uoLxmn3X1bvVT/X29gaH+NPJOuG76qTOnea485jikLshMMGv7SdW0UvmfG+Bl9
Zc5sHaSi/azca7+Wtl3S0+VrHKH703kZc9HQSETipae66P+bthkWw+dtVa+TZvXYBvTf4aUBFUrL
GwXCRykC356+1QnxUwowl67M7QzklZ0UlfX3X1tXBZ/NjYHZYCZLqRCxbgx/fZRWsjjwe1e8cqqF
gOTnu0isxLVIbsYxQdYIBCtEc4kA9ItE2/BUH7fcjcQOMhdgUUB7GgxH74VrUA/QsC9nIyLIxart
ZkJ+WVME+W52kEA08r/FdFStE+NcnGOkMJHIQH1WYDq7IPzPXSkhkIF7hNiWRg2KmU6l1mp9Wrpl
VT61vEW7QIyb8i1AxAJNXFwBIIH5QNv1FWEzMOg3gjWMJvApjBCChgA8s+zZ7IDhjUp0rjsz86eW
48GQDtqtfTK4A4Regp3QuyCTFd9M4krdWuytW047JjiFwPudkbI5DFj7KsWkaq/Pp0w+DYIsi/cI
X937gpYhxF6k3VEWnQSdLlNQbO2TwX7Ux1KqqLdznz+h7xvMaJjd7Regnhk8tqg3P0sNeHCXQ6rN
ELswLSQuKD7LkltFH8sePn/9ETeJ5RWPBZ71lcKg/c7SHmJzPBZz32h3zLrL0P+bB0wP5Jkf3pEh
ejLvQXCitpyfGYJcPxNGWUljukufmc6kVyyzwwtrWZRkRC0lPXPPFBaf8vwGVJO1zaWTtrMIVVUn
FV+pEUlBW7hYMirgYEznqOCsRgosgO2IdyZNLI6h4dQaxmSFMp0nHDU5X3fpywydHYds9OWnXvuQ
+rx4s/MjXRIHYk5lLgbr8A0lgf2jtbKInOJ9LoZg1RwDJyeNC+puwWyp8cYU2pJq3O2Kfbu++umQ
be5SaD4g5itYWoDBNTr6l6+6RtummkQwRpl6MnbUB9UuILMH4h0brLf8q5IXwFRqCmGOcj+xmaIz
JeOi8ITmQwesmVND7/TYvsOYQl/ZXRXNm7spHVZrcU2Q7AV53n20fp3WiHJ5lO6hwHIjHsFpviAY
53G9aU+nupdo+ROpoFw+0eycnKjW/wN5w68saggU9PRaH+OWwJkPzYQOdoWcHVi4qh53Dqg9g61K
KxHHzfBLgNyy/twnpufs4sHa2TGJ7xpJT4yeFFBLYkLCUs6QbpEznnm87DHKle4eSLKR7MejsCL1
Mcstf6iTygyNyjRGCDimJPiJdAyNGEG3VWYZv2vRJ+0dF861PFQjM0knhJ1u4Ck92Jh6L5dBfLUK
8bulgTJ0E49c1mqWP/kiJ4dSGFhaYEEqqmBKOoXgLIbyoUl66Yt3oOAjzhN/wkRhUGMUnEaqT9Cv
YS4e9Dg6EQZHPpv6im0PK4eZ6GgGS6seZzF7u8rhNOBs6+qAgsYwz8sqpy6aO92p6YHHYrt8vlyV
2bwlUPMSF3SXnsVpMDJctrphzEKfUUvh7ybk+cPbn3Eusn/ohOPDVRsf9biPTcXXXYz69xR9BARY
et/YcE9cU3sbPKouDkT8l05zl+zI7sfpk26JYTacEbNxFocysxRF/6/PThglRZYZ8Z1cp3IwHLXb
aRTjf+01BFP8ddNev/jrwNz6nbBO7VKGE933CbA6vbadz15O+eUCfzVsZs8I40myrhVQ+pgs0+et
y7RGMr+5WkyuVCAl7E02rJ7p3Uwm3qBaEoRgF+pA7AyE4YHlRQ8x6+hZVouDgFUkfE/nVhjjBrqg
MCL0TyiQnXIyxGPxq7qnm5fUzpTKBMGk2w5ScvPHY00K9B4I/1SsuQTyTdeSjQVbMBRsg5Xgj7aO
ak+csHZd8dmMHjgJRL65KjQuALtiZDlSP9Rq/gT/fpPb0W0asrp2vTWavLrfprouc666+rQ9GmVv
FRVuQ2X+iaB5Q2ZLPhJI959r2EPc9LJ2ex3BhFBud0r1pbJFX8syxw6XVV/eiPfA+kB4SqOI46v7
bO2eSH6JcyF61bW9MRJBOpdUnh2Q9MECPoQ+oVlxbYKdHn2bnBfyvjeaJqrf8neYA+XNO6fZo5oG
suLxn2F1K/nRc9WByWLLwKn7t0Np4+1cH2jyQ3zGCll3mnvOYnxCW4wAV+CRmM51/HS8X510YcNO
mKJyJxHW1ixy/ZrwKN8zmcfHZJv3cCqTk6RTMqWx+Glh8yMg0VpR1ArZEbKxanpmJHAR3eAgAGxf
um9WWgjoa0f0Wq3Pbo2WjmI/glyQBfubeMGotb4q8mdK1umlvmlpQKCh0lOI3omQWK68+inuDk7z
6056DRYSzU5t2TSV+gFAUc2/nWdkceqk4QtkuDnrPPBHAZO600ibheDmkHw0b2XKmKYpzvsK1tPu
MNLwViZ3PbLdXU8LQynDXoWbUWAw0ma6F9+e6eSacXMWmzWoUSGTm4s9qyL8pwXTc4RWs5FU9RFX
TAYG4ce3+zW/p3kr8M0tSewWRIrWDqsO0r/7RRRIX19buTF9xbg72NnD08aVW3X89hDN4jcQSEE0
yrvK27n53QJedqSq7dqClCskHLvvZ+05owHsw7qNxICqg8JUOmIx0suQzJU6kkA/bG8qvkl2J4Ny
2Pg35+ayxg6HHwdLmovLkLjZGALdVi/T0YoL9Kc3rHP9WkriR2oL6PpMqWloJAeo2uG8CSTreGp1
sI57UEyynIJZJuFXrqnY2nEHpqJvxRC0DVVb+4qIM6Ekr/CjjLFjZZh0j0EkkLWc6LOURSK95YQC
dQgUuWAacmovK6f61xQCanzRicFuS5c7bfhL0KZAIbJP8uvpDLFPBQihk7gizKFc/RpZcJExWYyq
CLzIw50AFUvdTuSpXFlnsuLPiuT0rt6hueBakzD9WYBGxxqbBDDBIj4bWb4vs86yae0Q8EWRF8bZ
NkMFb5VjUin8iia0dcoxPc8n+3XVk5hZaMny5u2O/Y46bxkY+JJnfkiQ3VJWpSTkG4a7yKEDn649
BEadxTIXo5vmd7HsR4T0N1hUAlK2uP4Y2T/4LIgZC/zm9hoYpb/ZQAbD4fpT2VOlFwli5E8NRdF0
1mIoPznOQC0o9O9bIO9QieqnI+mvYs4bu/IogUMjbjBynLdNAQkVYXg9kf3XHAyI89y+ZVgEFt4Q
6fLRvlra0gS0f1wekkdw7Nvc0aoi3pGAFnPDUCGhclf5IR+9xcDJW9x17WDMs4ufM4w3BI6lRjYf
16mkRJ192ad+Km3ZAIllDJAOoWe8/SrdBe8wttaRe5fkIk31qPGad9ji+IQL0BdKKhd5bskWceoh
ZDv7p5yqRCy4In7CRlGyg1U/bP2+daPVxsxQy8mtdi3yinuIDJaMHf2wHax6B+MH8JLGm9NRvuIT
zqKvJDYwQmOKo+RwOnMNKM0TmH2KaHfMPv1Jcvfgmu7LNY4MLADvBG97iOCcbeHy4GgC6372QbnR
V7N6o0uDuzGRjE/bAWaDDViOQsH7y6JYWkpmuTlXk/XCD+ZTPcgB/FfZmnxqQZ9Sifzm8BWECHgQ
l8mUwyPla4/GLwt51T7DGJB3cqWYo6xXeb9t42AxXhZaQR2NzCwQxpPx316HuoHLXPZq22JpNI9l
5Chg+r/ZeuSQJ0WnTuLu+/6IdublU8lgEtjcBcTPeNkirEBerpfEjxEyLsmQype2LzR/3COOs1KO
w0xqi0b9AZnVlzM31QRSFpY+/EULxX9suV0Aws0srEg0koWmJKSr9+Hq22rSYKPYGS9VyT/uMGLD
4N0eHgyyjkts0BOfDAzLBiNB5ToMH8UCnLfFJHFezseKHbXcL8p7E8Xa04Mjc0cHJLPOcNrddxR3
KkpersegHSaiZ9D0PL5qyT1yofaRwbw8iUM2rW7azTLlV0dMYzvhrLZmNG6dnc6j7qNQnTf5yKXd
Z+MPRhPXM6zz+Cp2jAbIW36Bth7DJt1ZZdwcI+KAcrbPRt0Qejd6O1mDtN0ZOJ175sAQpNOjD1eD
Kl/D5lLRUtJmJ2pA3ZWaJ4MwByOnTZLaABIZOffHGBGdCGuSPNZJmJHYJCDlbhd6eOw5QFaJmPIz
eyEZ2OrIj9RSq69ZVLLUoBj7P8nhuKlHSOTE+N3pPSgPE1RQdjnt58a6ghO+66GCJzL/R8uO47L2
FmrUHWONC+4hQOMMu9iDZqG+BpIM6SUumFQEp9LmG4cLOD4UouLSMgOdyQrqVc4owDmrbiUzA5jm
D/ey+91OavfCAqvBj7xy1585fLyAN12uEiclZTWngebSOuxx3yWSF2oDGYDDmAJCQi8YIAfnWBR+
W9oVpsRzQ3fM6hRxVPBzGtDTsQ8eajjc69zVQeRRYdExKjbkv/3ViRuroGQ00oDfJ89LK0hX4WQ+
qtL+s7Tc0PR33y0Wsly+UyGpsqGNGAG+AtJAp+YD6JSp8bhiUJzfn/0jX7eJiAA0vmJgMZGV9bWh
YTs1kgAa8LK1+2nYlncqtB9no8QW04TM8XIMtCCd/9/tICCQSQMsvCGJTN9ha5EWrAkoBQ/q/UHE
HBoUrPUvSGZLtl50lKj0gsAa6JVBcVv9xkdNWDYEcsNJ/92ImiJ6f220aE0e0SIvsyAj4DMMGTBh
Rs35S0e2LYcW50EGIEj0SlBwld6rdUeYRcXWn0eJA8d/QfdM5bxNRdDnxB3TbURo1FQJqQlEp34+
0gHToEr3CmU5xEh6rj+ZkqDnwDUAiXT4bJSJ7wcwN7oUHTxIAxbMOTlefyHKQcFBgh1Kjz7U+FTu
+nNSYzwhu0Xt9K9BAlLeVItuGMH7x1kHUCeeOxFSqvqmQ1YT4aFW29OZR7ukdcmA+ggX+9425LKc
ACf546asfMnhAOaPwMelQn5t5rkGjgxDHCUkkv+L3BklvvYppxYjCGFOikHsGUuIwsWMBEaQ2czI
h9HqjHPb/Q1H1IGZFgw/iTU434Iowjk/bUP57DazAuLG1HLesZMdlv55j8HobB0G11tsejAIXJZA
FdjtlSRu1wNMEQkn/NFU8Drt0rhp53CNaDof4tQSDwBro6wbfcDpKNml6xFniweE473OBca5DtXS
fihke48r+fy/mnsEGr/TVAYkO9FKYbiFM6Wh0jDAW5TKStGQqj1ceb0S7wY6D71XsKCpAuTxHSJN
5NmEnD01tNPIn85H2vjFzZpszsNQtcfP+zFrXxPfNbK1m7/NMnJpB6e7W4eP9RwbES/Mp6WXOvYR
IlylUX27Taws6yW0ltkyVjpq3EKpqrEzDw61EXMM7Zdg7/TVR0gzUprfkN3+6ei8ILO/1tPtE0I5
EU6mqgCxWYJR9tGx4ZkLgoLcR2+mIkw71XdhsmmviItQGz2jY4DcDqhpE4SJDGHegO2YeptHx0w/
dht+RfwjMxxZjRnw5pc74zFF1UEPTFBpmB+xdP9Xn+26n0sFCW/GOp0agpLTbhiG0GP/RvK9YH7k
D3cTqHhDrfxVmzZvKozE38phRrOqUd+z4thFA0Jy/N02WS1JCRRnihGQ6nivj7+jPenRVU5dCDmF
VroiI/qPTCO4QBic0N0U8HxCMR+XVWq5Tawi8s0nh6Uc5YinbHuEJk+VCe6gpHEny7NdMy47Hwfu
fpzlSMogbwcDuDASINV0QlnQGk5FR7SNBZttZM6M69XeFei5a8h8NpAvjjOWEc+5P2f8sXKCAWU/
/zo8enPu0ujAFrxpcakPDfzpsdi7k+1K84JMxz94etAWTw/2JYMcVmGwnqr+ccFiipq5rtwrKfAH
+Lsn04wW3TyNTtbZQ0WNsj32XHKt7zqxCA3FmalW3pGz29ldIsudBBXB6vGse7siq/5uezLEMgpX
OHMSm5Pzy1KIPvyPYL2D3rdUxliwmJGjGcakKPY1a0jGTSSYLhnBAPWTxHlpwI7vyiUIt+CcCdyL
6oDxu87jWbSFULPrG6fMYcKhMvx8BHIWVrhvh5CiJruDcfDGkyukEjnFqfYvlqjUVwCTFb9j5UAL
/3qhLh97mBou313yQQDO8XrQadLfY/amUCZjj+Ze4HSD4TIc4L87u9hUqGDalWGgD8GysCdPthBp
25jvl8XYBxjFg7vcPlvn6To8sQvFf6hKe+hUeeE9BR4oQYwufIVmVb1lMx1epHB3gILranbR/oCT
JWOothM9u/iR13FN9Tjtr9zR/L57m94SkFoUn1BFP7SNWoPbE2tgwUo2GX3iyfYtJEH7qa7CN5ex
kLgqbRA3+ppgX9FunPSW9giYjLDtgQ/nqBbg8snvZkphs0wlC993USz8VsNQ6nUGHtxYfM88rSbC
q+7bKIpMaTVc82rTv7dJWeRbmTYQJy080Ejmki+sUHAScIa4/wfamcpJuKpGOIFqVKXZ6rp7d4Yk
mQ5kn/k6+/lgs3FDkRM9eJp1OfnHE7234NAPuT85yW1/d7BpMHNetM5bw0rYe3bW1RsT8ygnV+Am
7ARruk53oXu321JB2Mqb6wUfakX+bMhAiKMq0X++WnCcTmyzAFaz2lT1QH/9ium6oxXCpN5ntN7Q
LT5mLEgaJiBE3S2EztTvNcjjZx+uuT3ON+izFh5u+bHiWnIC/l5APYVhvU0nDbfr3tXRyK3U94xq
SMF2JtKcpKNBfE0AEOz/1K5UtKRn4PNguNWFR2aK4sxPPbukI6afSCFmYEGikVieqLqZkY4g3mzM
mm74Bli3wcaFqiMu9ZKmybAAJa2rkhzdvwfsHnYjwHfPuV1hXt5ZHtHJ0G46QvGGTgnoth6bRF7f
ebmc2GQ8jnetioErQmGkwTiMeCEBxAWFgi9ji69XjmXowySlbLUBSKaR6mlLoS4D5ODSYSjDKpTz
jxlwsqdns5cgzNTuXZxLo/t8rGo0Zjs6HyWcQpi0kAZbN7m2DjC9kKlj3XXEeRZHduJTzOPuQmtZ
KzkbWwajQJFWjh9/9UBW8LsBfJFyhdoBl9n4OyoBYEOWLQJuTzYlIndKg8OR27t9AWNSo92qnrmB
XJMYNInuOLkcOOiNm/tFef/L21HIKIcqqQB/xPH8S52dXUXQQm7UueTLAjkHN6dKwxl1nuLU32hr
eKVE30drb0z2AP9IWC2OCuU412RfI29JC42myLD+CIoWi++JflcQ0wBc3CF7ss2J3VpxH+zFVjR+
pUsFFKZS3FxBKpSODyUCl0OmJSWUPfCPw3VWLXEAlq1FMv30ibgXnOrhDAlkl6yI5BW8jxdQP1R4
VoXwfD0krVlCp4I5YY9enZ4CM1nsCjk0DI7Kng2gftzmP6kd0Cl7U2vPaMMNavTqQxj/PWb6HgUg
bbqgCUhnA8Uyd9ifYAbUn1Ck13uzyipIGkoBJ382eV0k0kVDF0medKH9Uqqe6oZwCU/ABcRut1Ty
Zo+c9XoX3QlWt6/kEbQ3YimFVyu85a/CGiIKZEli8kI8f2pxMa7O2S9QLsdDADEzUU7czt0R9Axb
aPaU60FhYDupZ0WZebiJYCupeWX6BAkEFlGKTUphdBLO3Lik1uPoUUJdCmkMNgJ5Q2xod+KWC31F
2dZLEnarDnXaGUHhO004gFIwvfrxvoLwTMOWbafCVnVKxiCDKsFDFshw4ZQbyrQPwjt0Su6idZ0d
UM5duIxnFscR1fNzHtoMHI7+gjG44lhohmYFx5qxA33TURPqTg5/zxP8zI9XBiwvNQ3R3w0ml/He
OK7tbz41TUDyoGkva66YNzDNuywxbutjqOm2OLBTt1ElXdyPO0FTZKF22pwHoz2O6YbxowAUSfMY
JZA/AIViNK1gK8FHdfCjPIFkitemIpv13741rgQlOwwHD+eaS+CIt/aj4jeJ89UeKmbWhvepwJ39
bozSXAIprx+YGQBIQ+8jtydQSbt8o2L8N2I7R84umkDkAsFsdB8lkDZs6eA3GI5URv/bq1G7sH6J
psmwd039nmz29E45eLMJsAmWKJwUYZWm6+MjY3gcSCtrfsbgetSmmMtF6irpnoljHGX6oYS+XN8I
E3wMz4JpVUbnGyrjAT8TxFdBhaUr+TocF2hamA29VFZa94fQCM+yt5Ht831xYUvkvnrp5o6UeEPc
Z2vSSiY8R59AuCG2fmYrNCWtibGO1GL2bVElWZmq7tbZqv7O/dHmkyFIRwjRK9wzUYEr8NuYsntk
yq+2SE50LN7z7Pi4ukFcXtUPXk9fSOsU4TboH/q+TjO5PEFtmEmyrKI+kccpG0/lsU9C3v1Xp2FN
BlSUW3eEhTY8IuokzxCOWI5z6YLbN4m9DrW/m+Nfq1Jeos9Hb7PLFoVIi3QWDH/BAyOs8RSzwzdN
Wu1EWEJky4cT1gQd73DwDH9lGpSJu42GMOxoKCEP14wgJc2Wo53TVKHR5FKUqDzTDwGZq4VOYLgy
8c4LhxD1i0J6W4GU/vU26wNnKH+a1E+0IHMHNe8j6a1lEuhq0AR/Sj/qI766+RIyfBl8DNf86sFW
IWhRKkyKRRg0idp89OuueiVYy81dO9hwke9vG7IArKuWbLaytOb5ptW/kSkPibCxsZbe9m3lsFC5
JUyy77Fr4oKdRZOvL7V9i55BnvW25bW/yfCc+HwahRx/TZ6wtM4ZLERE8mRBgp9rZUshE2NwMehx
Mczj/agmrQPtg1aQ2QyAXL2u0nFj+z9bYVrAQ+VYxkoxRw8K79InBJ2pmk9XNNjeYqIG3IegH7oT
o6DlUPt5KX+v9NeDfuyNjZ92BqZmGASBY8YDMdYfMN9ZIR3upSkuzVAeTZln2w0AK97ArIPCf4Ln
WnbWg1Kaf53+hSLB+B9KmCZ7dPbAJ1uEGycBbP0dGD6Z80YVirbiwhoA4HnkxtutUOtxIstCruYC
Vy1QUeWR737OMkevT7O70S/Sv9a5kSD8ibG29Ge5zEOWHILwImuhMf1YMV56JusthMLGsfqyiq6z
dosY5+AXYeIReSK7zxsZsPhXzGoNy0hb2Nb0JyKI+ufMeJ/iI00UAl3B6xdcWPc6RPtQJAZUNOcc
nMRvnhcOnbvV1iKqFZ1SL4fUDmuogI7J3+SYUlKqfOk0RujEJCyrRLEK/2ciGoG823p3hwUTJjTJ
tn7VsqFc71ydj0+2ouLk4V8NOQT7k3xLWbf9oyJJHnetLZLLk/qcxE3SZTGB3hlZjAfoabh1kopK
afPZaEyaL8epMCP8vimyJEAAFk5yxKtZ5k6fCjwnr0QoyijW9XLkXAyet9eEpmXCukjLo1mtn6rY
VXW2yP4ESNeG2g9gdxCypODZGPctr6xujDC3FOTQURzdPV0rQd8jHUNib96PwppdbfgITtsXoq5O
0CuMO7BrpWGHt05+jCTjHjlXl5tKHGRYC6u3vfcoQ1axKIYvw3V54DTyz9eNqYOUfGO2byjY80cL
GtBUvC5qTXe7Y8kQ68TjPsZzOEjzdcS38zu/JWSVfx5503w3jQRx2mglBGAvjmbG9IhlBEnxoKv8
o21SaQDqM8BZn5dDOMX+q5ta4d5b1zI+1We/leNSHLzNYIdfqUV++djyj5qZd8u95nZbc4MRQOF/
G8sjqt+8pwjkpz9FmTWvrM82+TenXocInNxFF69W2nOxrvVEghA8SoMm9I9SrrQL/T21w900oLRb
888+V9JIU3kXoZbnBEt8XjnhpzN965jbQg+yezKsHlDn28VimfjQIwEX+sUEq8N9D2NA0ukQBv/B
H9c7QO+XCqpZFrDQMOtLMPnbHN6muoQmw4muvr1zJRmPgozY4k2MzOPSXhtdjveOLZZ8mqW6uQi7
jjbOC4lDThol6Es9G2oIctWKyVHE0IdGppzt6sAvjv6m3xaWMUoslZ4IYMMx9qR7ynq+GTWM52vb
d46buTiAaJd7v/APey3ERhePGQuPpwBnGyqpgn8E6WIPRbhMDVagIP3UM7KX9eYSm7ndF72tk46h
wZtEVDrVsdutPvv8x/M4JJHjz5/GQUdS0pmu7fjaERbOaYzCEIcrpq8cmLpGt6/UIg2OOrCiboZz
GDu4PcnhiZfN58UMFXCzXr8x9VHEvCX095Ou1X9ka/7cFl8T7TKabWIaQMMc5XS5R5htfopbW/hF
T2KJru20NkjweUxqd9JXfsVPXX4poHmjosIQTzq+AfDqySlQdoAElvqcjLP38xU2lxlWnXY0ZRyz
ozfwtLsgt2r20b/HPdng5Ev8fBS2O2BeenUWqnGjf9dSZVYA/pIh6xnJaHg7ZYVebv5zw0iRm7yZ
n4VUarStb49Jb8spcZRtDM6HxYbr+d8yiUuX2O6i+hdbRp4VDyr2GRtmpsig37pIe4SDtroyN4gu
ZYSl4gmfgo6LxLN5kJjcSl9cocwacJL+/szgnpIixHUy1PnuYSISDnyCDLAlMUxa6sSnYyp3oWST
U/IHYkK+n/nfjig6XSfMLapAHq7dDulVMFruYVbx1f8BDUjPUFkjTEiH9ib9u5+oImqlHQmbSxxt
fFwQj1kPab7AmcYAMO8Cjvei3P6eySqzLhAp1ByTyr7apy/OCOWg9bcOswBuJl334A1tqWenZwpQ
9kEwmifL+ePPSByecUp6B1F1D6YPH6+QBmlfMCllk1xz9MHEDHZHeo4TGsNRTqc47xlFXXFgC0/c
PgQKB7XSIdD4kqx5pmTj6q1ZbnsABJTwJmhgVgni8OjlLV64v5QKRRKaefGca5+0cOheQMuZAzf6
NYO0V8YhCY0qHC6yEiqjL1Uur5pLlBiEIoFyeEpETqd2ZiWWVLjR5XldscIcG+bHoX9RE7mSrxxx
xr8e8OM9UY7Bds0NzKa3Dg/i4JfS/GrmC4qCDhEd+Re+6ysygqCVi5yLBvcgvOXQCbJUHLo63HXh
ziI9H3hMev8yMsBc9kN7V8pJVVBGMTy815UnSW2DK/hrUkhcRiburyn18/ZY1L7lcHUUTKJnjArw
TZ4yjMdhBMKXdk1HfZ99QLX4zPmEDGmwvApBg5dmbInt0Eqdu+ykfNQq2dbnkkjJjsaexlRucyBL
QcOVI+bLpzzjgKr+Ip9oshaZR7RaDVySlYfX6SKb+Al99kKSfmocrlgprJTrXbxUFe90aJ1P4sD+
1cklHjQD1etpfkLSLDSE+fVWCfW2x+J+afVCWhvUGM6m7sOzppVCwatsvXyFrJ0VWFpA1z68YbHI
9TRYHvYotDk/rhmGwU6H0OlMNLq8/MVk04tv41OswwXiRRS5vKAZRQrPS17mH9FXFotcJmCH0tyT
kaRw/xWCi466b6jLy9RfLZa/ed3lepN77aX7tEFfbFoC02YUHDUxdcDlQeGypbB2EeLq2baEr+2k
NrrkcBBIaFCCo0mXKHuYVk4kSTJrKBB4eUmPccunyoDsEpw4OkMFp+eXmxtxQ2vROfOieWUwLVS8
HUDqTtl+bTegU159aqN6OHN8N3HCVxMcV8dMhUQTjbi86FhttSE726psEDZh3tHGc2w6INL5XciN
gmozh+229FfTbPlsOzjTJ9JdUYjPVVzILV5ePyYVy3X6GnyCMgN2+0t+JUlwOwAa/QW9O/p8Th4l
Ylmbv01rqyME8l97RRd/a6NWeY/XsRauhd67lDDS7yra7XnoWJ39crWjsJ8zE12P3OWRLp7dPP7W
enc2r9FQ0TjRouxi+9iC3FoyVe5cqeIqpZWNcRT/ul8CkXah/gKjnkN4F5y/AYpkAu5XwRRWcDHL
pJ1dpfsLkESxBq8pd71/yC4ZVJFobAJ0EmO4b+913JScuUIXkDgJGCYLPAd11xVh5RzOGmBsnODK
2nWzCAsd3pCDMaxtajboq52HUR4Imjlk2eMBjo8dMdhdSt1PBRe/XUen3a5CS5BuPinYvK5K7TLi
AbdgLeeQMHt8bSh4HUy7pCisdbuW7htB9oM/xX3cBVEgUxpd7uS/Ym/ZBa4x/XanoYbxgBw5YsyO
fX0gWLShbnoTZiWgtn84+XSVPcO7ByjO5AoH+KfGAvcA4l5qgvOQZUXoiJSARXauNuKCbXMQRS6l
TUTicRpVSaK7eoxsdsp5SqwFR3Wn0imd9lyqonJC3B8Ok5eWftonBKMulP4VBQMhudZ6DzPtqR3p
Y+6Ntxgnkvj/Zf/fMWtJJ3t8Q+hHW4fU299ahZ7c57qwxllz6dtB1FacsCfbbbkwGWRbQ2s2HD2R
EtkgUtszcRC/PiiaX4Y/8KzpnSL92tJ9EFHJ8YR+0ovEk/825McKetDNafZEBSenz/AFOy4GLFLn
DZxcYb8n/7UsM4NRgAD2w8b6AwELnD4SBsC+J51Rc7Q9+a+56HqzETU1xs+X2JFlUjz2TjYHCp7v
PkFyO11WMAIeFQihL+v3aJtGC+JVuDFD4PZYSvC/iDnGS/dnmhKVg40u079xFGb2uNLhD1jXz+am
SkG4AcFZMXJEKQ0rEK5xER3F67KtL5rCyp08XOY9/+ftXu5Eebw2FUw4NB42eJNuT6v1EqS+DZEm
fwKaqsFQin8pJmrDNOl2JrJbAZtmfb/WlT4OhVX5BEA4CBonhNDjyUok1uZ1O6yMJuGj8wpt9Pis
kaWBIQ6z+k7zlER5X6FL1OO8rIcfjrvWiluP5b8rm1ZX9rw/Qr6N1dFr2OaAH75diJfwTvk3pe9F
spduBrr+5Lj0lLR8uELSSinLHtExXXQgHdHNUJMG2iSU6Dhv9abd3oyXl3eSF5VF+OINLul46Q1m
cVNfi6LsUezY5m3IVM/aID9f/SZnc+XMHg1P6BqYImJqassLlfn1vhwmaXmrKVrulpvxOuLfDD+M
hn51FmdJsPv18Q3UDkv+InyklADMSv7OTozOQUJTTMPDXkf5PNvcwij+9wpeYm5nlE3dbV9jsu3c
VJulpKd6NyoSWrYzDKxSlEXvgfvy6/u8PDBxBjGtcbFeXu4gZYBlK1o4uAw1lEHpB4YlYvX9TgH1
VOG2d82Gn8gx2ezZR8M/5BuVfaolfbwak+pDndAZpqzKswk0CuML7PBJroO8pSO8Y633PZSd2Ttz
2/dScFaRLlCPssDiEqDaVQxNMGUmNfW/IIOCYC6e3pC1mUgSMQ1viJ5o3vjP0DDoPlNG9mZGh2yt
UnCBvx0XRuue6k4at5BzEVyxyZSBfmeBGRpa4CaqGnLEjtX3Pph9ohRw9YseWB2pliZGSWk9rBVh
JQWNbEC+aUzKvfy//gpX6m/j6ozeRtv955fButy9vVixc9pIuOLEVK/WUJE/QmmCRHsy2d7aHLNI
1iYzyo63b5rLuAv9kBz7C7zUYuKmlxv+/CFt0GsKbsYLiUUqRba9sHgGBr5Ljn1LUDiP51LGq/5C
h3vKY3L2f0kFgcNIO4ydIbTdvZf3JqkQdRfdyE2jDlxCsK5sCgJNJoBu/5R9bvpvsHxF2+IR8cy8
6cZ/Pnes0mq2m/0cmWlgaQ5O1Fnrl/YLxDYQ2RxsZJoxYcB2xZjDUIi7C2tOpCoCIPVBFIWdPE2i
a1fAOR4ALzEj/CvyvqHxOHCCkGF21bbDFuIUm6/Vuh6FIoXZKm+bTcTs56lqu9ZTppJHFuBOvoVs
NZFYWiV5xzP8eenNVACjBbE1jNtIJKclaoQ7AphvU0Gpy56V8jL1AI4TgtVmeCNDzjjDHLMDjiHO
HJ3J2Lav9L30EvCIQXC25VfiZFnHVneIg13BMTZBRjolWGXFxAiu6V2GFMzrxo19/sWPXxNVkKI2
KvvP09sP7EiXoECym5qmN+D2ib6bvAao3edj2gpgWjHgICWXh9+5OmZYP4sQIG+yUSwj3Hqylm+m
i6XQnFj9qq+jVLf3c4kz8L3FlVB54LklxfIVzZmdkI3M4bIDjYRXxR5pzpvLRZ/Uz7j5yoPKKv70
mRSKL4FtgWIbupEK5Y8b3fOYYc5cN8sbrtfwVx4HEfC3mY9o2BJ043R7bYLy21bhwu1X96bpbx31
zhkN/qjoYPNGEx8I+lyUbkWyxKd8k8j5cmU333jlNHLh56b+mf9Gzka3HhM6/WTwa/SbiDo5pC8P
0zGhVZAEChLi+MrzmNbH0szOlYyJvWPgpjgeKOa7Z0FHTikWfaYhkHsoCqdtbx4gNQLnMlPpbGuo
0SnGJu1cbamlQ1odGHeczYBPe6RmGCJg2/BwgPeAQtwd6QRVluAsxE4skqpVkE4c5OIwzsV2uC63
3f/FM7b0yjQuPGpqBMjjjv+fOtBgf8W+okDBQlnuQ3fd0pXQHKQkbxYhP0adAKik3Xl4WQsF2x1O
p3U9xF+HcA2Qy7F7cLnZTzRYvBzByK5BtFbZ+Yr36Aq7Q0ftC+a9dQOu5KClI3Nu5onCU9U+Cp8T
MQRqTIeW8jDn9qOrL4PHuvn0H6XkfskgK6gGF8zXQtc9I3oRB56Sv3+enDYZcGpEpnCBrwIF8PZD
CXArmHNgkebxTNq0WV+7q6gu3z9Mhv1q64whPd4kRD05bk0ryWucTFtjfKDvkrkeP4cF01vvtbnS
wI53A1hwGKPrcdd840Kw5tJrKX3JTXKi1lpyBNzDhZjm2lqFg13kIiBc7bhTiVA81fw6zzBpKafY
ppasq/d9EISvVqp7JEoqPUbbbBdK4bOuRK0F9jgOcLDidwbI7ExcTcYYHFObaMzsx3D9iBAojmA0
ygozYpKa/CKJ/t917Wf/bnWii9mtPsFI/jgGkwa16tOiu/mmLA54O6fmJnnaH8QbhRG1o6P9bnM9
kn/2/rDdWvJ4qlizYL37aY3XpGfkk7pCCAohx+eeaNm+29srB8gCcboGbfNFmaQ+toGejAdmYI4M
uODGz5xKMz8qbXtN99kHDpJFXcPWACQrwA/TeRCg4yQQEn9uqwGylSe6QiA5lx55PjCZWWjYKeWN
K9tSyNCAcS8UM1oM9+pQJcvJKWu87E6gKCj0RWnwQmHisuO6cpwZY8dY8VntOe4TV9fiecpGUAMM
T1LfV8sOdTg5re1d+XuQtSFHSJGiL5CZSxplGW+y+Lzv9YRI9FnsPq4UvKYS5i1PUXjT5hnXfPP4
vG6ff1vBwAg370EWxOauTyH0+d4TUfi3mgiSwVfRnP6MDK4kLmLedPYVMvi+mTxAlsEaU1HEYpwM
cdJltkgyVP3sdHk0nWAWAKmvv6hw9O0Qu7Pbfpm/jIov/VGP99SSNaVElgnj8yUpSb++CPisAIpO
4a15DM8taww2sNwvB+j7ndzjx3YomZ4XXiVWzfUpicDO1UHjeMj4bELLIXDAA05/F2Owwf+It4op
a8xggNyWfmJj3NpPevV1GPzLzA+eZs7SoEJZcBODB0hfoBFW/FCvwUQ0PQE9cNhK/aPOE8WA6Q+d
J4MdOFSZTOwgCkYU8EVIrW/aYAvsI6GP7UjYNmhoGRXb4G43M7DncXMN3e8s4ittsraslzVSbGwn
zjOQWvbrgcEveprngDwddSXjlNV/Jd+dSO4K6Q8u6eg8uDsbKQFtop1zAD2LCKZZRAfJ4gguBWf1
1ghIn2e171Obib88/bIpd7mY0jCp6Ne8DpaW9xjZPYDEcHwIngMhZoY8qr/WOGg2+Fdq+DijWdSt
f+tvLUif1dBuwcPBVy+RN52WyW3/nPcPmhtXkhthxRq6Gl/1Hn4vemtCwZP8HYMsLkca1ES3Cf6J
CyWOrAMYJjZ1tkzTQA8yFZgQFz4DqLQ21jZSTje9C9hYDsW9mI/sYW6ObRs7htV17CUQz0/CmcWu
kfqIFiezIKQQIiBOjpozVWR9RQvXoG2qqHVMZ/ma50wXLbi6am5anF/Dl6pTji8P10gbfjypUSSS
h88epGJHNOtmIIe3EKD/dtG/rMP65mdMTEMGsQH7i1DuRw+kYxzQnPj76RX18CP/EqFyWmA4ImQQ
qtjdUXMEAa1NoDrrPfuZJXR4TxAd86MvYVhqVbOPIP1Rr383G9SYDwq+gS0u57OekoyVH83Tn29n
LJ9mlq/6q5uwq+35vkU4E9+8OADIAENJpnYAjs1vdKUXLWCbLlS0InEeAvCVIyvOkBcSibkS7zCL
NSyBrjgLF41HZIv+iBL6IJpuYlzlo5CEad+8SUNs3mM95SyRrOYfd/aDMkRupwLgA28uYTTJG6WU
HSqMSw7zx92c/DVSxvJo+ZnyLFbw70K+GsRZqe5UJNakK8UeNh+FWEQ1mRUOs+wiTiAmYGjy/hxa
jHBl8viUkmy7yugoJ8oXyen/ny0/QyQS3ildCr+q2FRC7el5oH1esogFqtoRPoAq9tExWmWSy8CF
ZfndA5nMnCiRcKaQQxtjz5Aft1xKGElS43gkN7nnVRMJsFZcSm2jPJglxBlcYqdbUFcMo/UCV6Ay
2NXFBsaeGtX8sPMogydngd6MIeQptL8Am9Ser0sUCUbDOo1+fs+u+HVbJRT9VvAGSHvO1wbucSQe
vm9gBqEfYk9VP4/mJrD1IYlgmubF9NfoeC1MyFdPDqbfm+k8WeindvKE1Jg2IbAT0tr4npEnXVJb
4q3/OQ1RhfXXjLNe9xwfz1N62wqCuNbuFfMBG10e+ExD3HB2gnELF9ecHPqCs63ffWQh8RXXbinY
IP1ts6rMYApmq8+bqiZKUnhVjtTNiogfLUhqsdI95aav3ELEUQ4wqYQjM/wdnUDpD2r009QjIypv
cCHaonv0bo61nq0lZMCOLlF4Gf6i7EmESzll4+Tk723b2raLPq3I8yEjtF5lvhrhm5mUvCQUuhnw
zg9ApBYtGv/zp+YIZ51TDYXhqGX7MYYp+/jcLfoi6Hqvzz8bqZG3roi5JUGeALDjo5IJjje+Qc+r
hVezyzJMUQ0c+Dm8rtuOgnlrDxQQenGrxuA3XoYE2W75eosi5Vz7KHYD5rpECXCPfJC5QrQEz9WP
BefKxnM1t1fNJZqH76FxFR/eS2G1+CEEkRDagARKZCcPz8srnncQYGExJuVFaC9Wo32NEoM4oWZ2
De1UGrgAnykCXinunXpI7EkmueID0dyOOsBjYV565gidtsz9DF5XCpkUQZbf+aNMA1mVKBcabbYa
f4QnCuSnkf0pNsbU2R+dVXGXGp5K4ee9/JSF1XNDuyfanxNbYGgezx4WHhz0KcoXcVeupKwNgeEG
LEoYHa4bvB5gX9MVKNMtWWmurL9MxPhdHWGBi2NxUJOdDkGYBI7WkjCgbwsIGvwFUj4ghUxE17ny
esQ8JxEw6zxRnzCZrBhRhOEAXgcHZX5YWyv+CCUaqh3vHAQ+ByFihapAZaEKYULd1lasGowKjNrK
eGru9aIMCqDiasTJEDEnPaZe64vjAxVtS4eCRe5YIViJ5mT8yFl7ywLztqNomQGNG5bnQbA3HXVo
5bsZNAKiW4d6R2Gccknr2Uuj2RhCNztMXSaFhrR0D7BEmNGt8v0Xge7qgMOi8ouZZsQ/4tJN6o+w
ZUSFMfqipbc+iEV4tKWBterD/crs/y9bVTnM/H/tb8ArOYlO1953KSkywx5FeY0SRU8dRrohIUKj
LNQfbrCay/rK5VN4lWbchN44mtR5wCVvVwv6/ghKfxQpxuW/2g8yfTajjSOrfXuh6L0nsMNmE1dk
FK8a9tQIwG7C6oNAaqSbLMqcPUuNZ0tNB+noqLmbmhUtXW31boPI6Ga+u7vPFOg2AQez9YLhCPOv
/8hoDPuUvXbGFzaXX22a/G0RHL0jpgr+45SIr8/gi9vXwcIjdHEj8f5GAEQrbExXPJ1S90aZ37d1
JzoPZOXb5F/jMqbZzE7ZXoG954jzcfX90Ah4L131MzZAKhqIjBx6jYRhuDRJzq/PG0X1RpsRK/VG
sbTN4YyO43apOIeT+dmtw/TWOxxuRtQJuOJlR/knc2b4BIXp/ScHnawBVl2JOglC55wMZXzNjQ00
S+tlzAXPQBvswPIIiv3hDGZyGQjJ4+Jod9pIGamlK7HKP5Uq1gMjeMgzKKqM1QsNJfWIucM2d/xg
UgSsbl1stEwQjCNU70bPU58UzDCC7KWhMlheprK4PfDpS7MGiHPMTHbFU52RbxJG9CHJdyV2+f2w
AhszIdomYmv4QuTBDgVUxrdwJwKJ69bN+lcrORM3iRjpNMjCl1hcMCIaFjEhhe1qGBFokyGFrvDv
77JZtW19TpEr3d1SNVE2oO+gh6PDgBFTTJy8pYeCjM1r4XPU58KJ6TLiho6gKgL2K+SMS3ZmdBSW
MF3/RbmY717Sws+WWuMDYK3n8gb+AN6zt3BTzskplaBPkioDEW1KiVXd/kh5An4UkoB34OT0RgD7
N7HvriivkNWtYMD6Kv9YmClWV7B8tC5uHay8FGmhNyt2vkREALVmtukCWT/Fo8PKlWw3L5nT8nNN
d9q/wUBjVTQ1GhSn/jL2ttqfaYA7kMtv/CenqcCiels2Z/h0nN2+UXIoatB8Z/TpGP4YUgrkxMTR
3UWQQGRxB7E0dTr3+JdYX7f9FLTuhkdheqp3HzbZbBpLWps72U64iTICzkNPzslGOg5ULa8YqjMY
fvazCJp29JJLS6EdRqGGKDzjV0ylxuvAjBJGeVvlMrQgj8O9b5DUPeO5pkVn3DN3JvldMQsaBUZD
enwDelI8Gh5ebeH3RxIXqBgf26TmeBDijcbIE5C4oxpbznWg3kpyEdMuvd7mf4rxby/3xnyXy+lX
1p+4/8yXA+1KMrqt8cYzdgLOuojxxk8EZRvpBcRvhim+gkl16VXVxOjl48q5Q9bROZrMfXKA3hzF
yBCe+s+iT7hAVIWZ2moWWfhxGE96/sc+RkmbnW6xNkYRDj51ALubI0PTUy6iGG3dky+4+4wLIXTy
Z26j9Q0X2L0GsCAiJ7ntmthKCzJ56Krr4ggPK3NAY881Mc1XUsT8ySlAxCGhBh0qesphN+Cl/1tD
D2Lq97AW6APYtwg5hqk2MxfjJT/saZNAhiPdYQUckAqnAVxxp84+alMEVOTk5eVFIxo4eJKXArr8
lXMV8f21kDruy1KEOmuu+HNlw3kR8zCo53khVO+sKFiN43o25A4PVSnSwbXOqEya+J+oPeBgrZ8z
/VCJnTdSsA9+KVfJqVFTjaCUratAMHzwLHHus43VncNepOuRCEljuLSS8HLL2guPmcDs99sxG6DM
lg1ITZdsQ1SJOASDTknsFz6+xg2ATo0oZWZv0eioDchNa2jaaI8S4+0oImhawgKpv/gESGTleWDg
c0AkW5oYcY30LCUUhvPIQBSVtxIcNZyQmMnlPNM3PzDlH9Utpah2Yklin2btXmgUKrtFPJeZCDaq
d64/9Ngczr0r8M9XB8v8eL1UEd5/MMB6v1zDvurFLIwStuIelbVGjZeB6Mu25uZWEQN6qJl34bOQ
7IvuhDxVkRTEILD/G4HQVZrwu3fr5ItpMC0/X+LnWFzHfecWypRW5JKEV0Y0A1PBfAZPpiqKperk
/A4MeXHtNdndsjRofWvGS0u/LsTXWP2qq5cA7nzUSbrm2vOUB+Ud7CI/edGY3PvF6G03hAvxHkni
bMR5atDskIl4tR2re+DYvtq9JtTBmGYZfWMOsHeIiZDQcStfMed/VhQHsu4MXMEXQMTrWtAYEwMV
1aBcUZl7dxTrJlP2pYp/LdcuU5yr0tgO5+ltucsIBfu6HQWj0kFFfR5Lal3+2GDIxx6kRP3AUyY1
LAiBEYY40xfZxF6LHqSarBL3cZurZk0VJC5cE6UeHSjcRYdB/w1TWrW/NoW/+cqXUrPSVZPWXCgs
pnyENWRibYdTrVnViHvCFv58fQGOAAvKL9+Ax4tV80cj/5AwbBDZbTqP7yuYjdg/Qvj2QyiBNXCF
R7hT24OfXkRbSc0yH417dazSiECd4ld3IZ+KooKeGTXBImURJS9CrTymEJQbSzcej/MUJOv5bGP+
BblFplv90XwyEttWoPazptq9GmMBqlHvUitYdjTSwWdLeE4fh52sS3ikzYgZBWJLlWpLnRdd2Bl4
AGY9nri3v/YWnnFB1ZLwszH7gvyZZcm9P9YEJRLmk5zUC/xkBFgqFTy0fOvhu6sU67zc9HJoBxc0
L11o1hZbT3oJcXcDSOM3xqkNutPQzcAcj+Qv5vDEV67PHZR/OAeB7KKoYLzzprpA1Hn/IHa9TIlv
giEbCY6eRDinn4Kps3amwNMgfTXhdN0KliSDtqvj8qMBcjbejwKriAB2OgJdJ2e43BlVl6mu+nJ+
eSvJdCNub31hMGbpPvyUWlXaSQlZr4SJ06VFg9OXGOhikKClV6QBdvXXYu91KUgpnJDWsgfZBUFd
0Fer/2oakZTbPvDUqGDlgkXjidfl0s48SMN3e55Xeu9zjEf0w6uHL8q0hIXKc+nHmkiD+1JBNHzh
1thsPnQJ0gtQdpOV5Z00LSG6U18194vJWkrGytRnAvrRUVS9ohLL/YaYRz5477ppy229y3j3mcMo
79njOA8pRuh61QbnGTJRGSf62QdqiLXCEqoPL4dXO2pgb09dozu+wiSe6fcA1DXaCFjhJHPsgINk
R2HGu7OBqSL2tEq7Bcw7y7C8wWUFCaePfkBsxwv5c0fb8CzYwuXuUd7SW9v8Vl32dSyI0u6Ypor0
CVo4g4tLyJEeNSTb8nM0I5P9EwIyjoUOOdopczbYlfAAl0iSg35vhKZVLJuygJZbdDShFwcVJE6t
i/z0zQ/dbDKvHqTGaR4S/ehdj2t2tK1tGOXaqm+plTDSRDoVrfEs+kFYy5B+kvS/WWsYJnt2gLKD
Sx7k5NSYDWIV3p7E2eUkV8IiX+DO5YXfO2eNK67P2G7JVDPyYj36jzkKJvJJJcM4/om6Fc4g+Dav
9odzEK+pU2UvTkikzZg8ISbBaayxNcPFVFrF3LzSUYTypBH0V8CqbzbXbz+y+69mP7Bi1r4O7Oxp
Qwy5zg4AG+E/UfjqrbximiS4AkF04wp5KssLnRaI5zm/658nrlvksVHuR+p4w/RmYrwJ5XFu70Go
zhNm3IzSICmRspQ16JSvXIEGxVPVDE/RcZ9qsR28jkRrl3u9hq6ZeeMW7L6zMrh9g1nt2MALG8XZ
FQrpcvZs4lYPt3ym32TaaIgd/MLaO23HziZyREIBl5+KQhIyXHL/avetqojg7E8mi+7OhWDuHeWw
HhL6L3k/8vghWwK3F6M2472XLLOh+FkHtZKSWdX8aL9ae5yCl1gINxyedfZqCUZ/9PZloPs2KytK
oM6dmOZDn6pJfA9sp1K6YZyhU3cZU0iw5VcatnagTIw9x36c6gE1N4snja8rXNiQWjgk9Ve4ulPL
JQfwtKWvkZz0SRy/q+RC8EiBBqf7JRZk7X+d9Fs2ks0eaY5m3qhkm8W8odZF9chE9wGEWLPWJnRp
LMxd9Fz3aHwV7IdP7GNMvjrrV8a5zpza0ITwNnk3dULTpVbngZWPqHhTw4qSWUZNsPTPwi+CzRtR
CyHCxRihNXqM/r5ehiZ5AzxPPatlUGyWuXXDr7oz60wuubxlAHc/Fff5liDPCivomwx7jpM1jUyx
nloWF4gzqsSvEsdJqfodsdUv9iVXy5rAYF0HczqwusBUOy+iA0K5OnmCWK2P5dJcjvbH8hLeIdQX
QRfRo2baIvecZTfeXsSNdrXJZj+33i07t4pbUFV4CCMbpEzJrtnnG6MCO1LVKudUFUkh04jDHXik
pbovJ04qx/SSSh9Fj1oPW71NFaAh/ud7WfMUXc0838fcs9axzXHw8MTm8qruWClHaJYaBRwKIfUo
JCCwlR1B3SFZE++69SUGZktq6xGUfBiwuBSjLv6ZdKALKMmiEf8LoygVEOWoeYzksGFvxnsghC6z
PBtR/gF5rBdeK4dk0g3M17XC0pc8s8EINAGoK8P5Gzi2W20aHdl5UODyKU5IH5de9nnjGd7udzEX
68lkYw5PxTlrpMGkNa8VysES++mtztX66UuYxjBtd0OGV4ynYcEOAuiJ0U3DdI/JcCCc7D6A/PB2
NQiNvgc7YdMh5TJRt8Z3Qni+X/qS0+VKLfAExBsyhW1/7C+gVqbeMMxeIxx6OxMM2oj5QMN64wcU
P3vhqlBsGZQn4ELgOLdtEPENqpAN+aUEsPfQPuKQ4TE6bABp8Z8RyVD4Za3NGX3OIteJqVTbT5o+
mrCVWh4f/29i4f2pKNvP0MvrARE2snAlZM3X19vHCSqXPfcQyZ9IYGZmkvMb7buPVxjTVj4J3MlQ
N+v/CVUGA2QNyimryzU4mbhaTm0Dljv7jKKXds2nd2awhcKjvRNAfPYzrXLlg29BoPDqDIdjeelS
Eyy9vsAVsNc+Ex7+5yPrAOp08j1tXgZXisWgs8pxJ28bIz9CHtk8UHJ/tALUESm1FgRVldpeIUp9
I+1x7oyjqS8bLwu7EiF3t9NCpqOtVkVjGpcQZA6YqTBpscAq/YYRrL+q+fjlToYCCoLwYpAUU+VQ
BshSiynJ0WPtoa2rvA9yT7mjyShh+wV9SYZr862O3VjnU0UL/uvD+npeSPSJ2auNSEOWS5TtbNxD
Kr5mOjV9muTtjA9/aL0kn8cVfg7UzwqY6VK1t4UuO1DUFSiOM9OnTb5vs/l3g7wpCAM5wYrJwEq2
q53OpDB+q6G3TzdIipWuqFWV2L6AfyWnFhfgkd33BO/+sh8WlTgyMt2qsw2Dqrc1VdIzWBuIxwOy
/FKcopbHUQtAOKsHFedlgdQNpLgGbasDyxNSsCMOsvGhkzsOPQkB5IiyKa/B7aHbyQ2OJ4DHzRsI
DJCZ2ObPbERwOQlMz9CfTRBryDASpMDajejgJj2KsYinNyytcjm+QpSA6ropcvn3BaQdDWqhvtVr
VlMuFjDcEGmJ/0tTj809cnkS05v/u/zVrquIRr38eM73r/2omcwUtdARGCUc6/41CWcW/dtHGZ6c
uGvfPjkTaKtTD3OBsfnu4MIuhBlszNR3RFgjk1I4AXGYxIPadyxR0fKfWteCkBbqR63Qz4OyYZbZ
WpNl/uZa1nAi1M2nBWYbaoqMZZr5f5g7GkUtO6/+OsNZk2ZvplfMCwytsVp81SO0CYhQo9lFIzs0
tZtVVxWPEPPmqWX7HIxr4r6nF1M11cWTAcrGUFPCfJOOLkIkqq8I/mTr48AmGfqnrlZyeYg/19DU
EGXdhUo6oGPxoB8XajOPP8Z+48NXbEAojf5zxmMdfw2AbXuZwhWlKu0UByiMpM3mONBB8qXSdJ8h
OKH13SUsgUpt3zwEm1cSxScRyIHpKiPjH/2wILQqZIC1izcrDOXLhphpR+eZGpD40c4mzrkMLedi
XLdd/yFJOCFo5nSymryP9K9sVzRi9Qm1lSR3BVCnk1UxLWGgnYIorOhdZKl3XOPs3gseGuLD7TJx
y89M5FZHgerWkfr9RD93luZKkjo22mFZdFJv+xb17jKkUWYdgIEe5N5nzTvBYwIgpj/bmleDejLb
ikSdIK8DBDImIzQ+YETE4wOJ5Ih/OpaAuAHX6m6S3f3aPtPvYAHyThJ4t5DaMXouHH8VSsFrcwlZ
jZVRijjZFx5qxI3I1rxIG2OQBqviecbHUrwsAWuNiA0KbE+7aKb+LVX+HEacfFNMGiKGUX7QUS/u
V/6Ky4TVlTIzoszqEJ8Zuxp82Zzk6UOdQA0OEZ8LCB1vbOxieQKYNHRrI9wUnRNR3OOCew7LQlc7
ZMkaLEEb2+PAsn6YUX6Ut/Hx2kPk2ozgal0Xn79mCqGzNLb1odZer4hdK6lWtUUOVr1dPfmLTtmY
7FoL3xNMNyKAi5+OUur2I4PWgowNcAqFYbDO5B2PnAro8EICwnyokGLT3yal8He3eyfOxyXPgaRr
+ytgKU8UvsmMvIqqyAY3Gn2mRWdUe5E+jKb2QWpQutORsbuzKijud360JhCwT0xcm4LtQkKVaBVp
FXZSiJIMaO8RP2rLrD3tMMzTBikJV6ak2sgL3bKP17U51y+521vwnox0RnXXMAFCIU638yPT9cLn
JOQHMgLtXFzfnz+gndiUzOp0oWibZZcKO+tO8QVMW/hn3TkDkegpxbRx1pnP9oIplyauYII/RlHC
ItguAAbicEuDklzkiKMx5ak4OEejiDN6578Dy8CAZFGmb4TGH4YvQRTUHhnwgC8kOI2cyBmZwhn6
KsHOA4iul8902LXl0JDkf40Y4PLQqS5WOfPBuj2BIinUHuX57zmKgGZLCmWFMSS5Wa98yByu/9ZI
ZJgEMNCyT4Jd1KSQ5/oq6YkuLIvesb1O5htulkiN5lCdJDNh8fsZ1aC93RURZKekmbd2dHOeRXqb
hPi/gMdU043kzD3G9rfqGu0sE+BY5IIwzSBcZqioAxg50wPhDvo4r66GRN3CGEsPxicC/gkvn8J/
WCvedaBPNx2vc/yT2nxi0IpFyQieNVsw/j73PaUHFbZ41GCp9HwU32N1hZloYsBfKnlqKeL7jbzS
FtCjO2zJghFzOCS+oUKOix+56BmddO4MVX8QkTZj3V/YVAvw7muNwuTB38A38inZmp67UVoDqtir
QGVryCZDZ2UmyzBzFILd3BEoZd2zHD8VcfuNoc+iCL1PsddHGQswjQbK5cBb/cguRKq9HAJpMnoU
VRc1WLkWMcNdvB304ne80p9Y/v+77PG8VG5F6of1EVPJ5Y+Etjq1JktGZLumpnPaep6oF87UEtWq
KEIIPZqy/1iJKzgHlsO1MFQDmhmKwXCOffETCXWw7j8qAhPsxZO0juswFEsl1mFUT9Kt7+HIgBsj
UDYzFhMHFM3SWiNqcx0SPeNLaWyyvmSg81FoptT2HhEMhTPXkQjbJLdRgivsE/ihmVq0yQFZ6rgc
cENBqaDRC5QlneoIpl2svLwGFHkdwqboYtnaH0v416XQogfGE1gJ6JTGxvWj80sd5j3Sz+SwWy0F
CKrApv5Xv/r99+QIgEagPzFL+5MTG7twkb5IFb39HKAQtj07+0i/qHcIKAAlILOnv3gjBjOn8sSG
3yYdAjunJYWRPeyXjZUtrx35+rQLW3tQXuOr3PuHt3ARXv9MCGNKSF/HDmaxNZlubbK4f8b9gzZ/
13eN213JDFYonW+m3dC3uYIgIFXPvq6hmOrNA65Q1pKzkuXpJ1raZ94L2/dsReT/AbzXQ3WyajSu
V/Yte4cjJ8ZBtcb/mTVA4D+bAHQoktGSejwnjbjtPFb7wTIIS4kHiIP7+VBTlWMvSiz9FabgbQu1
jG3Uq0M3amMxfImMRNTicWyCCUCJF/RHWlJhjKHPx2KcNBMCZ1HYpjNACQxMIXj668hkk8e55UYW
JAhk0o6pML+2UA0CX8yZRv6UPetCPCraozewOayTUmuGCDDrWkJQz/20PHZ+TvTzfIwVU8DAnNQ4
YvzOs1VEHT70MV+AZvfUcs4wezcmv7YTDCIwrz8p04z3xNlLUZI9Jv0++jNEOytbwX+rBQIeTPx9
ZfQUgkrRbWgfqC6ohDJw//+knVMDcCNNgfTvKvDOH1pUgcyMNK9K4HYeMEji8PYqnapARuXkC5Xc
X+n8oBvTMm2zvqHQiB3fksxQworWEk/SKSwpWgduB65Bg7cORDvnQtVwsuFgkYRywXjp3AsBnhct
HXNFQOiciixON6Iar4hn2Dqm/5mOEz+js8/k16Z28VYKbAWMRNUIW+UChGS9Osa0GXyVxc3URMRN
HtH2R+HNN4R15UyWRrGt/GhyMIBtyMxOp9JHuf2K/DA/yvSZPPZ/39Do21UV7oxXTouf8JENYpCq
GikTtySweafY81MAuN85zXND7NMjGU4Z7ejVk8W63hXhlzNW77y+ZsFvr/fvselN0O2DR28kkUsP
s2tFzeVGA0rZLDylk/3yJREzguNleWIcyoBqBS6Bp8Irs36W2h459D8UZ6Qyg5u5F8SJfKFlgPD3
nHAy8Aoed4RZsIBSfTHxjWtDxd4D2JMQNp7vvGLd31ohEL4vdyj9zrSOeZHkfk19sG2h/5hTHCbV
4YG048Wt1FzQuIc1sdkU3mQaolIFG8VoU9cJKs7hye6ABiKjmH1r63C7P4Tk/FFrbaPy7HPL31C0
izaESh+ctakYo8AOlqyqnqm2urRiZO/UHEIQbeR5LtrWPNsrmuxU9noQHgF4rkS2FjdZnOZvpvJB
1MMzsZpZsSdJUoVj+UHFX1CEOs6VWj+tye9L3my8AQyT4BYagtiFp755wdvnT+EFH9yeQHNbGMjb
jta8YXerTXdTHnntK1lTLVS7gSRor4hn3ZNVBSYvPr0KHOE1DQgUx5yAgogpDS3qOtjK0JmoW5w0
vKhmHE/MB/IxsQ6Mh6PzAHsR3ToEgZXu9fjPKFezQGsoTobox5vSaXzlwLjvQ9Dwx0SOJajk/jx9
IHXdswYOp2GR61VnzUpESjC7zqfQo0sDqgw1cHLVurZftYrgDkOeUaCnOsCeMpneR+GaW0vUGKHU
ZbdVMaUBuci4CccPj8fsGpk3gFtpkxZp5NK1z5VLDNRqqZ9wyXlB4NbQi4vUv65x79QYxKmuUp9U
BVh9oGQoOYszgPK19ZC0vUc8uzgoqXHTISKd8m2E+mX1JolN8Rj5X2vQWpBbLVLCGtbo+0hJ/fSz
4RAxubpWpiNeBIMYr7qtN0E9ySuiiH+3mjpCXLLPhirkIseji1GYsRtLR1RKmDiktgQk6d0sxW/D
BZSuWuMyrKGTJ/dAbnxqjKQy7/0h7tof1MRmirZl7oRePaxru2GntH5QAULh/ZCwOnhSj4vJh57t
It7R/QklaSTX06CKFZZ/X4GpuAByIkog4CmHYjAr9E5UfgmXsIwCWHPCx+TZDZFd7uSRJMNxELu/
N4YxjS5fA+m41DCv9IuSqbKLh6JzyLkfCYsd8d9z5ZV3qFRgonWL5pPNYxxho+5+/BP2cpW0gNIc
tp+RkCpd3XF91RkkvChp/OFPHBINBGHSzrcPaKNU4sao/1tcls4nvTTy5v/Zi5i6DShrSDjnBefO
1K/WYDSe334TDH/xuT3Ya4g6Ty3hS3MC01aXUpTrHpAYMoENFiiHk9S1VwW/wmSbKRbl4pierqfb
1Cam4FuY2Y+QfVm8ee1ml/sGMnWPSmKewT/GvH6W6IkNfOCyzwnzF5xox0OFyzKFixI5yWhHEeBA
vdWlKkMSF/u/ScJKEbVS098/fnNCGuPV1St2gccmG/Bn2SSsINf9EBon3JVzGJq7pLBaMWFPSe2j
IKbhxXNEpiXz1ScoCrfjoxBFav/8ZIfoleDqJkVnBNwmT48uzuqG5/7tjsdtXvhLME1kBPrr86qH
ZPPUKDdFKjU8AGOYnx09bWF1BkJVJUjy/RFq5ll05qCRaD4pLhTm3p9X8m1y31xvl9qgmSI3mWOk
DCnQxNBT/GyO2ceytV7EKLknHQEydczxw5g/Wh4T7QmwWKBQdLEPRHRVoNwH833mpPD4+SprFnKo
tgHIqXH9sZDon4PihwjhQpy7rUAH/CRQz0lYQCLVWQmXw3xKdYo+pZPyrJnqfuiCPsl/FZ6q2/tN
yBTsZVF5XdWfJdKUqfLNSyakxCn5kUIh7lnCZ/TXSt8Qy0Xibe2nHxNX9m0uVJ7XlDK9Qu7mZWUV
0PgMS84cyaBrYhMtA7AEFWmDfQpXy8nI/pibFqnPKAhPogWdOSWff8LuxQVfXyfW4BeQ8tIEYfB8
/BEaS19W5xb6guMGt8d+AG+/MUetUZwG7BFcfdMAxkCW7odGEFt/mUNMY9Vv/seyfIiIruvspbP7
XZVFazp42oWmnuJO9ZGg9KG1b7pa95QZBuPcR9QvmNr9uG+MYJaQPJak+3RKXHntE65xc2u1hY4t
9oT6rJQ6QzCxFDAacJ4rGAj0l8UKllda3uc2XF79+0WN20EEQHbalXeFwodMCT8vzGz1EGN76Kw4
AHRDE5RRb+ivgtTPfNMqsW0UPYRVEMeuZS4KJOyev8RPE6UlhV3JnXVoF7/nFAnYESwapKpr9UtT
jnQ/FPit0B9Y6fbiOznTWXnu2P7veR1dgQjKtSnwmT/05zjcmZqmM+1E3b50otNen9jq4llSSuWx
jI/9GC4tXhk+/upFRylUEZKKTAjH4+UBB+dibJgBp7YxmxlisTlegHt9ymKV44PkBGjJ5yp/caQR
GtgD1NLVwAA/gWhNPq1zsy0oQRXb9YyJuqdG4SnXLfZrWzmwg6IW6HBAHkqF+mSiPRclz9zVD12N
zvgLfe4hhRgpo208hgUF+uTKMA6qw6Sn+elY0waTfqw7AEWH2Y5yZRrWHbtFmOUmZTNYGoWWsC3D
4W4z91sReU8IDdt6kFR5hAA6McwmkdYa8zBTfuHEqD8hAPOeC55figmsteen9AsYjii239vytmXr
StXDESHnoX+e5pbbtNWV02z+IzvvuAX5huPjRu2OKO6jl2sGLcn+6pn2FnjnuIUzIYzbNTC2c/rT
t3MrT51Bg8eJ0zXo54FuR3aBCoIgv12uPONiHhvYY0aqg6rvMEXnbjy8eLlGuhIZtJumArCkCVGJ
CGl00pwJKEzRNbK8TwdifGiaZvmKkdRKAgT9sQ9qJ2WjrOX5wuJvSLO4YKEpotMeBHCjwn7oE4J2
RCRT7gZ5BFzkbo4oSHBoAnzfcLJVcop/Ik20VktbUhSgNZBas3JvskIyOv1Uwoyai18/BrYd72PO
XvP99nE++/iu+PXxXRL6+yXk/xtSzmvgas3C8iCD6PeGTA8dspdkyXtBE5gjoMSOJMMc7AC+i+eG
6q3krO9i9/CLwiG85x0/Kn/miaBt9ZmgxnyjHi81xs8d9PwrnHI8Z+tbkgO5p17ATYVdPGmNOKYH
UywO0tveV+h3nr2W2Zbdq4qBgOUUl60cW5pnBMaM9EvZ2ebeMAHa6mp1E1y188hVH5tWbpFck38z
68p6HiYk/EJqg4AG8D/4on9os0HH1W92LiyrVN7s+ttLwt86KptKh7ZxCr7GJIUEspb8h8SmxAuG
fENfG4R+VUy8QSB1MVbXDFaIhUblo5D0xDLKQtQoztiMtzYLNUgpuB2NtJyKJKG/td6S9GWzyUKF
q1nbTzaBAg/n2gjE8GgrRrBOjhhqwtlv5avRUMpTPx4Ic0rY74T6GJKf5+duNAhHa1B6pFHYQGIs
wSXTKoZi9vVfB3AjJaLQ9BCJsFgyCRd7aJL6Pls7ilNx+wTzGF8X7Jji4BEIsywnF8YhkXGV9oxw
3FS3g/+UzEYyZkpAjb8Lr3NyPAPMjtcmk85ak7a8tn8r1F4pJA7QwaHzpTuO+zWsaMLP4t9H8jCx
55zvJLlFFzroYPDzzFxZice0aSo5Bcn0R8cZvdyAymCsgFFg1HLKVARbC+563gx0weT/Mz1Ceeuz
jJtisRWa5G6i+17GmAqi4rEPzja3v78I6zR20qIcXOf+cSuLDJ9BtPEmcsZhRNiMIa1miwi0EFjF
LmJPXMztuAeAXR8qmKLWtQlWjRZDjI96qYl/vD5gJK2f3Zvts+PVBHFaqVhoKqMI+lhYNYARc0IU
RvxpDBW98Nspmh3UlVkowQJv7DcZM6QSkm8Xa8kft2xZzaMcYO2EwBttPu4I+zAaiqA4JSx2b1Nt
6/DLpP/XJCrifa2IWlyMjp3YP2cmbwA3ccHQc1DnnyC+2KDKXd7XK0FLXNfLKXkiRrlfDLsStd53
NMoU8SMa3PukEOWhmTULqVf0UMjQq0gUJzIsqCLs+OJTVJ2YmShRkTlOZXvoPH0UKw4tcp14kjMC
co4W4uq75411wZVWo7qmyXBzmu5X7/D1rbK7hChxgj/STtlirrp8MgVek1byW+BJaBt5xriVS3eK
sfYRuTmv0dJsdXaLB/fO61UuZT+wTsMbSolLt8BuV8u8NIyiEM3aBgknO0J7eKPLlMKLqVpVkpJq
eRESqkwrSzrr7S03UV+bGGxsK9SrvrtVkWFmQYcBZoE0o2aZxZ3JlTbf38g1PJn/LPOmcrGWLkzF
fbWqhzCiFikkVeL3lMwFHnXNJPfKSx6H+91ExFP6mReCmJEKd+cEAYPyoiecEtcJ+4T3P8rC5t+p
hTNAuyN2q0o+BUMlfdST3K5KhA2YKSDZnfcA3CERuNpxnXmivlPR21TpTklOVQGa+HvMKH6AX8gG
Yhp4zkEUxJyBO5kf1mzhAAFpWBDetVHDj5kt8R/HiAe10JeYe3KIQPDOEyDKbnrxiiYSZN+7eKs5
bjPV0lXlc573v6MCtw8eWY0So7vwcyI7vs/q3Utxpngh6G3OREWyVJifk88w9kv1gnVEkJwqkyTC
7mEmVz5jalCx33riXvUv2oCfzyfkAQJnMRjmFccoScr25TR3/Z2bLHx37Ct0kjcFgiqZarPV8aRW
bb9qYU8TUozzyWRORfBPP8ttJD6y8zhy2b1Sn7LqqR05dfXNgQz9q/QtDJKtfV52BMU1ish1F4Tk
6f1YIqHyXBb1RvhASmYyAQy6BZNPoHawFJWNM6WHdIiFJC7jlvivZUBZNhwZ40vzP+jS58iatxxi
MmRmHh5FFGBJhZXXCZLSwYVDluNTAJt4uh1XMDMgnZlpnY69F8xCE87OKD00nt2gRgzGuiv7k6Pf
gQR/fxomZ0Swtzn52NzctwKuIKIsomTqg2HUiTrDs/HzVDzzAzKomZNMwYKM/LaTpSJh/3//q4yN
CltuPL0M1dzxKLWE7gq+8HMzzaISmrJZyOHkny2n8aXOEMGkQNBOiYchAXdHh4vQeRM6U0cZFqO+
/2qSNZPSKl9hacxuehZknZmREIn+aWijfMk0AlaW4GPOfGnX0BBhNHSgzF05hdoTi+CyU5h+kpgc
VmcY76HffH1yr94Y61Hcokm6XCmqkM4OzMUnB9UCJF2XtfdFw4JcrZAnZi3exZgGaCRKfdg1gpYM
JhQw8uQwlMPbWR3z4UhLF59SNUae07piU7BbhNmezUjHaI9DwU5m8RVB+O5z3/K9w2Z1wpK3ATZH
DVE4mmCGwo6xGwiU1f6KM/We8ZVyeNwwF0XicEMda4Dq5rvnA5gcOqUvWD05Vc/74eiiu381oWaJ
QY6LG9oPiHplGC5d/1tMvGqQpxd1HPtiA8gxeLhbcChlCTSIK3+tZnkMcVZp14pBn5hNAnqVe+EZ
1rfbSRZPQFwC2uyf93Lfnb7pLw/W7IDpEqF9FyJfj1aHbn7RGr3FatOdrZUmCqXE8bXFefRmA2JB
55GqRZxWQ1On/yrPX+N9oyobkJbFK+VlWsNRf3RennkjzoxlD+eoAV/u9yDlCrNLIIm6n6ioXQ0C
vfaYSpaQ9fczMc6cWvqKjBjcAgKvguQI64jrzDN9P+rYjrYR6LlRzct/Btrj9YQiMsNpwFzghXIA
v9MaCldKaSr30t+WwF3bshub1uraHtGG7gj/YRsjbdH4Io3h2I7bw1NMSLzz2OlbBuNUX9eUirtf
N9m2s4TR0ngCS6PxFbrOc0kz0kB9kqbI6vKrc2Ptoej3NylN6YA3781Nvepv/5OwyOKuFQddBWAj
P2zpYmkKv5GJRmAfJ502htk3JTLi0Qhx8ooFhqomaBJ5nA7JSxLhVwLsucD93WtrSgIocNQvbQYQ
HQcxZFXiQLtpjsABM0Qm+iYyN6JxVInaV9iH58x7UTdwJ8FBSa7mYfz24cJE24jm+7EgdaROqhfl
cNmAYTRSwzGRYO9iJid10Ce9sfeuf1zea1QKcx5a96IG9qOQp+TFahevSZnhk3An64bcGxlZiPxp
N1tL7EtTK9/v9KyCUlEIOn9fIJ/qX2Fzv7HFY5qPRnbrWNwOEZ38maga24C1ZzA17EoX5MVQ3kC2
ooo/BkbeRRsDgFUUYd1KXynh2Bj0Ob1u61DjZUQsMDP90V94FzQivPR3T/MNgjWXXH09Hp3tV/L/
CDz7i34yMnn7Nq7J4g9KOUVX9tMwONATlHNAXO881BkrDwv4T40vKS0N/YgzIxh01GHBb0596trt
wrYzNdqlT+nuvVsQ6suny+AVW9Rm/1cdyXBy7ZM3WXuedqTld0DrtEfLdRaZtu7i3lJpDMdHW2+4
W79sTNFWrvUr9vyq3sHUIEAmZZCUjyP/TdXPNcAUy/wQwINel44xAtOZP4i/LZHXe/iQCMxrJEbF
23l/yGz+JD/t41gWnUJji0m6KIFDYQLiob8JJgjySvCX5oOd75C5iU4vkm5HZg0AcQWq9iNbrRUt
3igZGFkjlZZKpf8hC/FiDDc1bzwvTqEym0OB/0DvA4P7YJxGdLYyabtQp8vmJJgi5Fbk80+aTwWv
CZ9pm9j9JE1Snf5mBAtdO1w8o4C2/81C2AOv8HCiFK+U4wLoG6tqCnL4yfohCef3WkUerfLkWLHi
1Bbsrhk2kBqYULOIsPfgNosS5iLyiIsihiciBcMEHOht/bJ7Fq7NGG+GCyWIlxWEvDeqOnrIump/
q8j3ocBnKZlxjHsttRaUvWpd6q5J2z9ZVsinyjM2TRiQTU6ywyRTRDW/DU8CHNXlDAhCb8cxg/o4
fXvNb2mNjluC7oac5AsC5CulYsVoWYn2EMTZ6T6OKkU2Sv1rpbhxa2b95/1kVyFras2CS8+gxLws
yn8U1UeuSBxjMai3oN8TrmUWxyaovJQ6fqeoojwdTz+/DhylPsDnGuqVzSFBtzAGl3Wm5D5lAuOU
tkoyzco5ghF40+NlDcw2mrUP0/s0klgVIX088G+ekcYTF2jxgzQO6XodWPhkzBXxaPfEbII+VpkZ
ehgTZDk8PL/Mhdt2nYpUufH8CjdQtGuvWHWk1PjFCgpvKpwuDWohpbdDi11DIdMDpRB1Z8vdyE1I
DJgqpIYQFR9EttCuNkeHlAJapJRrFjRlYrTpdGZoCa1XkyFDbPoy89j7O1CM118w2D9VX8LnBSIU
38ekqeKquaQAf9wXWaYuDTdtlI+VypOJvvDZEMGLfzX319Onrt6TyBSsJzKShGjgVspjGJlkrUHM
D7HDELZ9LbR34k3Fu2JdwvftkbaLKjss4nZfRl8T+8mLc6xlCrpMqHc9WlsW3uuKQbQ5Qcyvjv8L
OqNCkdvLs5dp3m0awZ4VjghLZ/VUoRcWjEzNtbR5Cu+Bd7yyhJHHpOgTwh1HHyTIEc7VD1YAHQ9C
8z0UFKdGMn208TRE3MkyTBx59EO/PvLD0bvjaOIehKM2LsfZii6PXiTGQBMZnP/iG9sqlW2bgCxX
uZDNJ87X371xH7wSBL0NxozrS2LGq7yM3rc417s8XIcJMZ514ma+KRMqXFmOMFfH+faFvna5ONIm
mxAIKA4s46x/WmcklPNTfW10WQpMspsG0KUH6T4/dNp/BklPldWNrnqZBYo8eBy5k1kFfBgH1Ap1
BVOAzez7bG14B4fKHdYM+7nefFCQ0sRwrF2w0siWykqmRiXxOdLyflwXbgqdbgV9wgf7jIHXrYH0
FA2LfOT0623PBBBc8Hhk7zHn/kbUC4//JaHxIp11r2I9SFHiWgcpqZW8lrOUXxe/C9qsv9TgfD97
qri2fIoRxtQU4kOs3t9PbT/maA3IMTrawkcBQtcbj0IoRnvbwMtCUrc/Vj1z9vsc2zAkFrO18QGr
QA/tPV6U3+8JtbXdVHAZCnY7fLKF7a5SQc2RY1SlsJBSXh6SLnkmbe4S+ML/ATzfmo66J8mpsgCw
Vng0hsjZ3vaANKt0phW8Q0WTT8GH3HF68AyrsDIOW74eOIWa+FLtSmdMeKpac1nn7y7HU5MnXRcW
D3hxxD39BdW51lCTMgOTIdaPcGEXgH4/9U9hKrCAfd6PN2oe8+uQ7L48KEfqXlfvG7aANHOyidkA
YAPKTSl94g+EK5+rwzr7ahXq6hQefTeQr5nLtBvn5/evTDQeEOp0HKEqM/z//Vx8nT8QGs2xrU4L
XwhF2N0ttmzR/fViBKdEUSIf82FhWTMdcAkRAu6y3ClBIJsGv6WIfcNflxHnkWa7bvo7zgX66BAM
5Vx6PApS5Jkjsv3hnHQRchetyPK8Sto5NjoRc7izwZyWkutXYk/aybX09K14uSItXr077tm3/s3o
Ps/7QkE1zxkC0cw46oQ2pDsE3uztBspjnVqHZ3It5HnrflEUjVdP2ww9xboyk6t8xbGlMluKQ3Jq
xOrPtd0aAt4V93cvVQtHFM+wrQXG0yCXmrwmqzafiAUB/TSGMbqgOXpOmrPOgMeU22d7Pj9pMHWU
xyW0+6KItkzM1CBf2nF+OwsfrvrH7HasNvUMyxUcpt2tlw3vWrq4ErYx0IkC/2KXXtD+M13Ry4DC
WUgnEZTtoCjxQhGK5qNU3J42XWythuA17WtMHsI/RaLlQYKSSGbllxy5zUYfHSehOiO1BLOAGPod
K3NmGHyHk8x9twu6msrY2X7TWEUOXN0QQ4QpuGN79WaamLtac5t+JC0lSwGB9dZe+LLrl0BH5h6F
FJIfbzwsSnUVse2OIcjYGuR9EYM5Fsy5MWiC3/rlIuYuPmhnbKBzuLh1U3ZrCJIZSeYYKOSA2cXb
eQXuZ0srz4SG4zUhtA4CjSl7SB8oA+66Ja2SND+DP7vSG1Wz/Z2ZTjheg/lsBX87W4u1tfFHCt1X
DE1EUCFd8IBYcbHMAYUOJc9SyzPmXJfwiAZ1TB47kwuyRkKJ9SYIuZActllR5D5PYa71O4UpU11+
iHGg/urxOZLKZ1hykIIhXwMrb0D3svKS8JJcu/tPgp9jBhQP3yiB0S9VxnlySxT8NZVxIIWfeklD
ZXWgijFJ4laPv13dABDwNaaL19BQoFY2Qm4x3fQDRMwIlctA9wPzx+7dXU/UzhVXQWIBkmUXWBM3
xILTkWtqcqyMcCZ1shFMB2TEqnnkS0tB5cM1py75mg9FnHwRpdjFH0ffEGzeh6uztfwLHiAZM6LA
RAiwQlElkoJjG93ylPopgTThAQxIW8PfzY3zMv18PRqy1xZhIz19vwhzpLnqJtzLOyvZjOwbKmw/
CqK8MFFEJkX++OXq9FJIVkGc8rS3ONcfauPOCBYWqao9SO/9yiTxrrGDgba0UfRh4DpKAaQXQzgK
T4WgqM2oJtGc2l9CFGTjhD8ZYOW2o6Tf+dm84xXTmXi0U3efnSqysPl3vNdudfa4S4b3NEiy4Y0T
okds2/8YQ436cuBrR0LTwgspN87xmzxNBhx+3Dz94gtu9Ni+KjqoySlTcOTCve1vl0unJcYcD5P/
fAIcuY9g5Q8Z+Z2OLh577AKAPN539DTN6CGWvIXiyOvI34Dw6DwtyfJOYYXh3DBQNwaB8SQvA3tr
sKu0qA71z05kAhUsZJc9P44RUjuH6VHIPeIh53Dqog1nZ2TWbUWDHpOdnsmgspl1AJzn2NeiEzM0
NhoeckNrK6dTS3B6uhORah6xskCLayHSAur6H5Dv402a++wEt75n5QII433ehEG4WZBON4/m+h0G
yM22+OeB9Y7G7UdU2nu95lzFT+PLZETj9i4LhUqDy9rMWOhEWGfL/3fK018qF2lUNMEuK03AcbL7
YE2lpQYk7LKeGWz/ZybCUAK3grF1h/PcCqoutF6hb6jJ4J+LTUNjbYhb4UIWR1fkvlj9PSUFKBqq
28SlHDy5fzXAue8doM0VX4usgznCvbjhtGCpd81iepPaS2w4d+hVOqe+bTBqTQSXUO+vqMsLyDDN
HiCHWWrV0o8AKLZeTs6tIS6A692Lsm7Pj7xLbmnMPZUHSItGZcpCduWREefbhhCyerQCZn69W5ca
fWpvmQXaKBb+FDbuGyqxBXQy7jep2Tn+Xi0R3LW75klYDvtg7zZfn8CQefu29UxJpunpTnb3qEIz
X8iS+WRCWEqRHVR6GaYqyIsNxI9QFHPUUlSupv9jG73kXK6uk/PzQAYN4CweE7tQxZGKrqGM6RcG
KBh4hkA1PrcsfWDFbRi8Yg4/l098xLn3Tjm47UIJCRWxZj4hyrm9yyKQe/29BNmvZxPE6mZUHVO2
QsjnLjIeHjO3/oA4k0EpqLOTesnH8XoIkLFrutQD6MKFx8fIYR0LbiAAlt/zl2pnsDLEiZfQ1gp9
eDC4kLdB7JMI7TrhP9gRrfDzVFgrDZ+3iLeKdslpM7ZjgdiMD1sfrZZtZ9DFoBI4x7+mkaEGtPmf
q1p/2qiDmL6ubt2VptH8itZUnEdl9FLPOjSwfNPqwuJ4NDPNGRFIhqSsFOqHW63Ay6PMJ9vipxLI
PnPnIOK7Pheq390Njz5Bfcg9Tm5jw3yl8t5S++4LzD7T1r2yphCmE9sxBlELQH+AL4HzzvN98jo3
9PnRvPhyPavcA7F5B4cRQaD4tPn6IOzb4DWY8MSKt/+MEGX1xcTL0A/NXjU4s1kOFRf/vWPQQHja
xdkUE9kPVgIaLowfUEnJYnSJihvsQCIDrtChWMljfa53pYnVNDryH8owsxZXSmpT3g4rRW7GCt2N
vT9AeVJtHMTHw/HZA9NFMa3HLjUAYt0xiLi5GjwT4kYw162YzhXBdKoteGd7IaUa58znwh/p+G2N
Q8oRXjPCozQm6WGMXogIrsLzeKyxYvCQc8a8QT9RKwYTT1aOtXsYFl3rKci476lVgQR77Wov5lxc
aAJFHWN/FTDqyXK9m6yRPvQz/DR2kOiYqH7/qovUB+6QFkzxlYX972CzSFvN7n45YzXKVVYCyPt5
BJlYstz4suanFtHJS9FA7PCmJy16u2eBifCLsCTbhXKb/CfIAZvKAQa9IsP7x2Eo2MkVMGCXI/Lj
VVtJOGRg1mNNmpN2AjoO1XdunTxF1wxVOun8U0JyhFQtRPMGc44Gll/MNNGFc1TO3QxUOSGxiUiL
efqdsxY/L1xJvIQ7eciX1xuS7AHLYMm5Jywb8fLdYeXq2DmBw+I1ldpiH5Pgf6chCyg6fI+aMGQI
wuXQeSHFoiq+zyvPCjq/zB+bedxpi+7nyYQTvle7xi9Z4BBAWqLblAnNc4OebjAPLMb6vTwqLnGT
Y2cPx4Gv41zAFDsHJ7auIzHWGU4ZJ4ATt9yIriZ98DB0SW42dTIrmx35UexCGArmwIim1eN/5Q6j
jBRDicln2beeBSC0ocigNMRKO8VacNwnyQd/yqweEDGW//WkevdecrZAZ5pmdFbZuhMprYKlxXTV
MKKkkX5/ergU1kO2hzDMqqIXUna6ANswLW7drZoqLSxNPwoRbe+xsdsb3ado8sokiBzfu1uQHDT5
icK5j57T6OsXhjNkhAeXPY5wPEcXWq0xdaNyEEcd6ihXG9GgWh6l4gq0tPjNvBEQLSbd75KMldL9
Ti14fO2ujEm6AOo2nrIgMSW15MLodiUmN5z/LMjFo3xZMTh5Cm2lMkiQrwkAnP4TjkvG1bhrtRWx
kdn56pUGbkKSa/TT7oI2BsxVwju0sq6Jhxrh8JZXdmD5AKrrwdSvavb1imSE50/fvwxnygFCWDmM
tq5t4hMWIyOgnQgJZZzSe0AAThpsU71biAvOkiErkvfeVwAAkGH+PoZz2GREhZo2t8AttV7pT0kR
RvsVDDTpR+3bKbL5R7AUlNclhCY5e64acwvpwYWUihFzjOjH1HgGlne+RCva2uz/2/Ey7e18r7NE
QGyLLPT0rzEO3ATKMvjUOsjSOwX6a4i1aNVrW8ZuQ7YQjDVbabF+fkonbURR7Unw7IAcyjNIpgJo
SD9aR4HPJ0n172Sr2DA2c7GyXismbvlcDlf+kUcyEJe3bAj35XpyTvM9NroOKJsxjSlrkCeVM+CJ
pnkaGQPYFzdPXFzb8Lb4RKU7YsWHRq6FPHiX6V0hLeYXHnejymnL4eTo0XQNa+MAwWAmnPnI9czD
cs5FN7moW0yphMWJCKJ8CZTURAARqGa3fasKX9ocGGvElU6DGTjw+pMVEmMHTmRVlK+T6xn09IMk
jK6gQ8YgZDZfoRy5lwRLd2yI24FAWKFc7f9h6HkO6xJkgcu+ktwULAUs3lwjfvDY9LHr6DSwzW2w
GqSxBmnkbHbhLAUtkQZrkKcrx8VUhlpJ3SgMBEKh4WoaoviF6hp7YOClOGs8VWPby+wxaYMwoO4l
wiPus8GeUaERLRoapN7afY7N3xN3fAmev5mjAP8sMr0vgH4u+TkMGWGx7R3HNAJKjkihlOj7Dl8+
kXAi++Y9fBIX6wIS/ieGOo6ptpG7befueiLki6djIlClnRxEIIUVOdo2Opwrbq45P9ZJ6oTYJqdV
C8pvwd97AkII6b3bJ1ulGnBrxuLpxmx7DxabNu8N3iLNBsuXYUjoP7mn2VQMPadExv+nBop4RdLe
kYpg3K+xivkks6MxzwdEz39Id+/b6ycsbeDrVsghJ5DdxR0yqvDfGLNC3+eJq44zV656bupkL10Z
BPnhJ7NnazPpM46XXwLNWld9v/nEWE4XP/GaalhPR21oFgJOeW+QltO7zlNBt+CUid6w7Px+D9dE
wg6dU/JQ0CpL9di3s0XdyAnmCWNqOwxsnAS9TeQxQuUNjUDZt743uuWiddvMiDdxYwrL72vRaNr5
RsH0m3gBi942anzJqKdlFtz27xZ9xM38eBCO+ol+4CR0/w8w8IWVG8ETNH8wrzF1QgmFoZxWqBTA
IVLlMi0lfokd7VnW4l0ptX6KGdKxl+MNeqDnxrVXgCCF1a8fv3An+joxHjHFwLUN+2F0Clm0bwgN
WEJwqzbaKirgPjAMwyYr2xVhpJJkDnQA8boNMUxK2Y9JKlk610selCJelRjjk9SyyRG8hMCfZDhh
V8s/MbaEdP4AfG3O52QD7+4wSdUw1pkQywOJQ/cfbaRuVKOcYRVV4aOzEdKCrxaMeIr8W9e5OmFT
0txL3WnS68OqjT7LT36iNuaiJ4FhBk8jPLr9u1fs1DpuPXRUZEXn7tfsFeW8HkmaO5xQAYsPgZzQ
sP4kyN7dsdWzk4iTTXlfYI0rfHQvW+mREoKdT0x9dsqgznRz5XUpc8qDnB7tsuGA8KOO8pCtoInm
82aP1uFDN9Vj1DKylfne5x6JKGFguDrVgV26NggQKLEYgBE78CCkJ85egx4gYmL1N6yrbmLJiNEr
uwh2ip5Txlx5IT1QST6HrCqSYbL71BkMRm4xx4I0CecDMe8g35vrkjC2hrUVvM992cKFufg7QpTZ
0hkcSE1yBHExmqhuFAaelE4dFVHGA5m8020sJGp2v7g2daJoD7uFqs8BRzzA8OgAd6XbfjZWESjd
oNpRZMuLzZuXDhFVJsDciPFlX9H82dnhUXlKj04dRqPRQgDpxNPollOiMhWuduJt8BACqap0Bbe+
57OoNaRdXnizxAzTyoat/QOihwBkRXqeazFWYSPmcDVCVMgjKrtdyLWnjVrptdL2OzvJZHB3SNm3
pQuaKJuOVLj0vTv1Cts5cBlkJ2RgUom0tQZyVKe9DBG2+ABavk6elI16HtPfJ7TrKj9g5WOUbcRG
5tUrFDkzaLpkPQCKxL7+VCLJUxd8k7OrxcBiYOpcMi1PzYmzOHqS4b7rjBx736sRWVIylDxl/FOV
DzzNcouC40baK89ps6aPm4M+SwYMCrIqUBySgiw7IbDK4NsI101V2+EmQfKcs/SlK10M4ciylB7c
sy5EjEjqRVIPQGli4nuiwXPVmYJQxAJHqNs0izclqsz0X+AvdetqCchinEDvGkhDF1PuQDRpTSqh
7yCZVcykSSeKWeWE4fD1J7+SpZngrIjtsWBlgOMBSNSX6l5GexEoFzj4IFyu2RGn/lkPEJY+493L
rv93nnqsCSQ6cYIcWv6J+qMZstToglcSJrmYmlDkKNgXbADzRyExv7uLZiKGK84hDetZhIZlvwqe
wlfrgVazLmNbOtHjUd8PgX0N6GLV4nZtBZnXe8lxhKrGbFbK91KRQt5aBGISMNIaVIyjo749jSTM
klKB6kJkOtGHfdtq/QPl5QfByBlpziDtraWgboVCQ0oaS+mzgrDdTvEZqhpiABi1ONG2UMDNDhGg
l6uKlayOne8+MUeZX48vcLPDvMgrRQp7yWlTrQYkc8eC+p9ejY2XctFn92zYvXbArcKf78CV8HVv
T0ISCcKkqJUYHzQ8lUKf3tfuZnWfDVTLAWEDuDGMzce40asBNHRqMXsN9fApqGTAX5ihUyMuSTrm
YlhBv0EZb/VWJb3gc/JlmVYA0pHSxztyg2FkNsStPREpx00tmXjVXaPDng1tZB0ypMMUiuiHyGrx
CHUbsddAtQ3pAnhglyjbVo935VZepoSWnONK4nL4J2ZdjnFICpAs5pjCgntbz/9DDzFPbGT7fazj
k4eoDWXECIpW1dMEQsp1eiXVfEynXhia1/iyyCfGR3XI+/rCd7d3xNYu0JK2uHld9k0ATnfXAcsz
M7e0sXhAlumm1/607oh26dc4Hu/jrwhvgBx00n0bt3uP+LnS+WDRdixEBrSvYW7VdeND2EmEQk8Z
YFqdzFjjjVJS1EkGOc/VZpfbz+j1wMhMRs0Sq05eTeXk7SxLYyplMrXX+saQgQlpMmqjcdZPuR80
cbumXaiNKlq4UgMjA1ZooF0AuhVb+PypnhVwHV/Oy46KUoYzpm/MdSSsk/MF0AamEkoHhLuH4+W8
wo3oI65wNaJbmC86o0THML+D4OG4p5bJFXZtjc6NWPlMva+350PI5EapoawCzRnp4SuwTr0fZku/
KySJY87jXvSKh4nRU99hPjV50LYIfNFq3rtj//o5wAucU8BMbXZ+ZliRf95Ni65wxWlh/OB7/INy
SJxzxJoeo/io5yAJf7bqeJFtoIOI1PbJapbIOlu64Daw+i1ZFvBT4QxlRtPGWCxbvV/astFdXzXg
rh0mkGiy2KGLZ8FlLWWod49/7IBfJb7nEhhYwwfxZ2JxIX5i3ezSAeRUvNkk8r1SrQAO6UJkwHmJ
4RSs5Dfj0jGQ1s0t1OnX7ZKheJGBLrvJAW68h2GmgaopCgXR1+3ECH5h8wkqkSJ+NQ87QcXHNOTH
8ExhNoXISPG2oZI6e9/1Ss/22svCUlKqSOI+8NxjDIYd6iO4PT42TQQK7lrr4IJ3yBwOc8hgPv5f
XPNfRjdgcFq9cNApZl+kLCZbHpotkxM3ZA1y65GMlupI6gMXw4K5scx3lngp8rZwYioirWXBZilD
mZfld9qyFv2giC5YNp15/uU3C3OUzfVbdxegATL1wyGV+j99SLkLxCt/ptnAY6fFnqxiEyWIiP4V
4ZMZmpYCqBc0v4BageqySolHFsVvYaqT+zCp1X0iJZEPAI4Y1kTBAJOpNsMoEgUC4ZW0YM+VKojV
oTcCjIFUlapzfYPky3/7QBH90Fs++dreSYPekFJ1X48EEMOZJV8GYJrVpnlfTBA205hm+NcsxPwz
xO2e/F8nXj3QMkiYFWTEW/41XCLOThz+Z6cBfTFzw8v69yshzIojehbTnUSDNREjhkcl1dVtcbzB
wpYCGL2Ax+t+EPCzXwN/HxSCVD0KzH0+f2ph5fPh47UQ1A+T7bZAJG7Y5ieZrY+cFf6KTEcDP7A+
G95cE0UtXv5lrCKLit6wcbXdOc/JTvrqak/m/01bMqCi5bsVss7cUH3B4QYOgC6fkh9K3oA3a/Lv
okn5MHPh201MGR3ToyhHSzrWDibAZpABmAQPHNYxgQ5wkErw69MzaOEuqqxBL2mMa7Bg6mMkCzyn
tttBZEkSOmII9sU2KALzXBtNKh9dzA8GlU/DQQ7EpUiDG+kYIllaTQDKaTypbOYf74KNuGhmSpTp
qjbuKLRaoUjlflyFZxj3EIsAxFF1v6yDKpqda210FPMiUJ+SUj7RO9nYlourg+bemqtSusmPzVtN
FtXvVD8ASXsVDlN6i4XKiaBkc+9YVteVp+xsqKzPeyaiUHCm9iNsArq59OB6Gbrpbw9/URgte76I
AxJXky0jEX4nXCmddHsL8DkM6UvQkjrNajeyXcCGpl4aq4L8GMsqihBjeYb8/u55Ife0bKzYGXb1
vu+hzaG+4+YqSa4z4Ioe2mTPCuTV4AjsK3n5f2AcYqQe9QAOvi8lnyR3I9GGjggfDabt2DbhNYjF
fLYYRZ5FcqclVdcTYUgCn4ESmE/5bkCybf++yf8r0N0C2/uX41e8CHP+Eyx/B1cg/SOHNwJCb1zt
OwXpEGBm2uKUd9EHjmWB6eGK4cCJHfcr9+GV7Pbw1S4/zsOKwQX8pScQ5xEKtDeNTCiy+Ad9xM8/
uGVR5cLKNx31EU5mWQ17DuVntCYSeyiKRNusnEhUprqqTc+Yvmb+4h/QAyutOlLoNXoD/206gX3P
EtTLO7ckLXgVI3PUF+ee7lh8BhK+8lpXResBnwAzuQJ5/A4gkR8rFS+FJfPHb1ZiWLKqWU4T8Gvv
EH7O9ErgRZddGJMiNXH82aSX5UgVyiSdWTvrtZxmp13kH5MIvTdVocCduQPqjOonUWweukOO4gVS
s+xN0i66XtX4bOse9y3VeBI+aJXwTI5lA8Lncfek79iRH1Dj7MYjBWKoR3j5e+1G6PISBlY7fO9Q
p1EYXAb8n/FWjDwb/83666EdHFjxcnyIgfwtuFMs8GKdpUFGhcmwWe/qvkB+k4bBjOE9Cq0DvOBR
HDVzTDPfjlcKqLAOqEqazFMLFzT3PbEee7IzOtUXVl+E6CAQHUsd6iT1mo5iHRX4Ly/+RGtLNBbj
5vQVe63xnlCpjPQ9HNEGa4VbORop9QYiQ1a9ms1Zu5AedM6MHFqxEppKkbCdQ6y97pjDAT5nPgzq
CgF6dQwAeM3Mi7HwMmoMBLPmDh7o++vIwd4hPeZV8SXZH0dNM+mJdXssb4E2vAJ31KvUVewzKoMe
dfEhPQ74vvwLJu9zwbbi9noeTOD0UilZNhQvgKdC+fbhu2DWmv6ffzvk4SZ1xiJXlTq7nfVIKgq0
QpQvCU13ut8a/loUP5nVhXZKktsPJgHxlXxBSl3fYfVpYO2TgKq6q/VG8yF12iPNwGqw9rp7RJwC
LooNC4EWLiIUlA5ErP9d7Al61hr2vJQZE0uFDmZp4RB76GB+uCoiyzoHc9QugVErIKrU9Vj9Qn1s
9YzzA1gbxoryC8u5luFKcUDJPwuFarJm3mvRFBfp3leclm+hN0ExFQDA5vh1TCCyjbLitwuehnnQ
qXVHROgarvX36xOv3IhNrNh7tLdb/TROOyQ6spHzGJ7ByU4jlh0NNh7AKdiYiFyZljSoZZlYuPT6
tN7jUd6z/g6Al67F/bn44XvYVJTdzvgF48E0sGL8AKESr84OZ8e0S+Z+dAn+tmkbwxsMatQC7XFr
NTyLpQC8/AcVNw+/UxIVZaM8P7LArx9NQOPejj0YRUGqAzEJgSlTnwABLTIarhbO1FAXc14K/y1m
lsGLQ3A1glD4tPc6VCRLxP19oxVTZaBv4Yx2t8C8YkZHaehppAfta1htbl6J1M8fglZ0UrJV37a2
zLT8WeDOB9KYx1MsVGwCzvF2Ibu91HOODvnTq3EyuowKuD+3cresJ+8RU0knlgOdU1xelI397fwA
lf0C0e7Y8bYCOFKvuErxCjknNe318GMYwkEXEHLoVqNcytXajZlZJxkdSzBGEVqV7pRSBH/tDDzS
KJfZdaCFNzwagUkBAjz1Jhw+sm5qA4nEilkJIaKoaLMiXLMuGkY5esm1h5w968Li6tbFUcZvje7j
7IK02LekpXECmoHqaDCEdM3DEj1RG0yM23h3XkezzGnUoaaKBYb4j3NJUg5msvDEFOjsTVdXdtxc
m7tt/fN5KE1l4GFs2Jnan6u8CydVIEnYhSqI0mICCMbzclEPrvA0bMqHszmSHxiAnKEwZWzc1/X6
cVmPNyCqn9hKdugdh+4zZwGqCNdVEi2CZeocEzmBoNdAyMZcf1F9/KBSVpkzBVHQ5ixtdBF4CaPQ
Tu5UrFRarke0L2+swriuEL5Hj13siVOErqUkuGs8TpyXiOFvZcEnxaSbym754kQw+pNbpJOko0fK
9esXXrypgZIuw3UaCKtBOL5cl4AmyUVc/qwYJB46c/XG2QH+ueSBuMUgP/YguuLIa+jd7qd2Sl+X
xmVta7Jn1GTlziITueQTNySJN7I/oiDuYTWcl17LvMnrgy15L/IumkqARuNvYhTQUZc4MXVyKQYL
kjRH4+CmNq1GZbh6d+E5BYq15JI+wPeVR4Wdakbrds0oso/ePHm9aKskczDaU37xHwGOOYiXXPBa
p6Nu5/wfOuNqOWJeVCOsgK++GbdLkb30ca0oSjsPPovCFig8fI/uNHDaMZsLXu6nVTkkIKCa/EFT
W3jQeaRYthMJA0yPuCzmjmOiLHQ5Rn48iFjte6GZ/eb0LRFRwLaWIAk/pVt6zWg4xu3fgMQFMajJ
Y5PACT//bomtHPi354MB4oCo1WYOH/rbbL4krbz2DTraaWxfGcZY8zJiP6TXQefy9qQDRGklL3Vk
VN/wn7p8vVXfFNszEBDV1IDExd9ba1sV8gfIpDH4VK82lqldvjq16pTCRdgUhxECJHT0w5MPj3Fq
dT2V+Fz6ZNGr77pixjz1l98/77zGuGZlk6pihi5GTbVqC/zVq1WVscoO0d0Kc6MwMOAryrETA7P3
0YOiGHOKy1484FqnWUf/wTL1sPokbwzZXPq9fmjVqPDiw9Vi69M5fNnSTwPGkeclFlVZxwkSH+Ct
e6Q3pOVH+3faeI3kdYXVqKrB2ZpMORpeX3XXs70efux00AVNyb+duzqAsPUpBD/2fhk5ANR9vmQW
112pGJfK4Q6WNdlE7jNLff/4GPPNeeTZeFooQ0CDEilMvDlkE0UxdIuKQFozpve6ldZFNPIspIdP
KjfNI+Kx6EczMV7MV1Z3bFoXyXYuPg60nc/hwofAACXwdhlwUaOx9G6Kw8rH2CCjwfkQXg9iVWyu
ZJCPXwBCKGaVeVWiWK1o1tJhhxtFmlwqZw3VuQw0uYuwmq8UK2yl+T/XHtjgHhj3zFuf5Rtgb0bm
P+q6KYk1qgXdDQHNIwLSryGiicZSrjpPQ7KPzuBWXT2SLnamuvgvwD2KdfAUjBzDXHNxhqznHjhx
4nZapkwkw2+uYGi1o9SKtYM7pQL9PktvZWZ7VLsuiJn/tQipmgPNRYdD6ztsXXVBqygk3omExqV0
gkX2khhzCV8N3FWG6LEo+BtceEqR8rXoR+VenBeeuGBLEyp2weJgQ+DJ2/1jKGHB9BrEdtaOBI5p
NcbViuFrGNT5YRnyrz4OHN5c9qI5mAY0E2XIVYv+7IkvO3cKKVN8J9djQb4ra0HcRBrVPB39IO8x
2rKwKKpU0FmZWnhbYB+KlausIWIEX830Sac36yP8bhlbrpq+Gyp8H/NIyvv8H/3ZAAyUPN0W5Mdn
C6rkwmK4vpry0DaprAaKdkdG+H6Ji8U0cXYXu7nqcscOcvIp7bYYYqhbBjw6MPqsyaTaujl8vofo
j+vY2YGxeKMyYD8Z5MOjmoyvcjiqEsI1sZU7PDDMEnINbdh/tG4Gvx4Dq+vQjesMqJfGuAtHZ54p
smQijZ0w2n75p8FXRgLQNdIPPL6SxY44h9niNrxrIEtD8w98r+9aeoDHvCpd/wCPjiKTbGUwrKSR
GwksGJay6KcPR1IeqQ0f0qzhAXjgY0Ih9OLvUZLPJ9LSqwwunjneT9b0RFaoWYT14ONe4rwrfL9x
qIRnKNBoK1ELgh5lHm1XjBwCMC+4KFkrpx71/kRlxkQKmuJ7/S1iix8vtxMSLHAb4apdQvckx5DJ
ReNJbu15jnaOaCIcdgXxKURcp/8HleBoDv+C530EV2i4g4RiuaLGdOQxvKR/1kg23uCmcKFlzFHd
pfHpcRLrUhBgPGBeBgWEOTlF9jwK/gg9i14epUnX32FV7q+T7h7mKfgNSkJPEJFCinFWllfhSPtC
/onViMKHpxUi5ck9qpiLH4ITVgflr/zg6OH520S4qjNHwvthWzbTjEU+JTpSiWhn7zm7OG/cZTBi
+CHKg9Iu+3nVHyiAhV0OQBsP9DUxIVeG8yquQQB4EzYJAExya3Fx3YCbkz0bPOkCLKUm1D5RlfY0
ljE7+rR7wctYATIzrAj3Vpuch83zKVECPMbd6SMeFA2X+F6CwlNigCo4kv3Qfiptn+9lUdZgF+RF
kmu62yiu2EMIy44sQ9ZArxUKcUktE5vpt359OpcMOrAkJtq9xcLjbU6TTpbaSlVCgaKU3rmArfLA
suNXsKrtb9fbRuxBSEa8hFLYehz5JymPQgUi68hAx5HWXOpROdyciRBM7LCiAvOEUmuBnmqjYztL
CQPa+XRoFwYkxzitKKvhuJTErZdhU77Pcls+jOq4zxUOJZuGQOFYheDdiIWXVdiWhKbh0dIFWokm
uk3xTX0U7yDkHuQRl8646kzxXv/At9r5YRX2yF+nYRDyq6fjp3WU9yNPd5DhIgRhfmLhMF6JRGpq
RTnsEXl3tQsbHZU8Trq0X/PuDzAl7QCpbMW/uGDdDCPNI+qXqJVQMpcCswlBAvGiSHTrAN9OrQOT
CrL7ATCABsDpV6ViiZ0rPRVX3ErPmhnNCsZ6HY8P+cZG3DQHPlyrpimjCkA6eZfG++bTpxPZRltS
foj9gckQ5Z7D7XK2yGbDqUL/MN96KQru4Q8N5O5xXeE2K58+xKu+wSUrSvHdqaD5GrmAxu7CKkAt
WJmgYnb49rnbJBOUMHdLhW+xdY81MzwFeYvHRyNzTKkTop0WU5U0g9JX1SbyD/x8NkzQarQokrbu
bBW4B5kiDz2PvXRSStr8tXM5vfvfdR32NLRWfN7+nOlNxbzQtMHKuKqrABVrcAnkbKAHqVOxNn6g
GQODozqNwdoGObVPbZ7FUQsuCaYNz2iil1zYS5QscirqxXVWC1HN7WwhNEM+S1TgpP9J4XX4YL+0
g0zy2ZRN547OvKpQIrEmVnGcDSW1JyaZq2Hm3YDNgRJyNtvAROWW+85Za5V782lkjTYxEx9ZBMzG
AmFLA/F98eROl6omX9WaA6LlKJIMx//DmnN+KsxCvx+R4tP8B/5SHRJKB2gadh7Y5PXFgn2Zb1g7
obZVRyy5Bn3ynIJ6GviBNYgjrmePOEXEk40fQikgldwnPzippf9R439I4vxDeWmJgSzG7/quWX1I
HQ1sqFNj0WlSviY6KaFgD6JMtvqNsyKrtX17CznoOJVhaXJ4X9OL/xleXW9hBygBADruoucNSo7j
B9XBlNM1ANJgE2PRNHHZKxn0WBUSRI8h+0c2bvUBs4Nfp+Nky9VNBjWiYM7epjJq283ju7DKuMtu
dzVRCFlhowwdiA2FCFsGdn+YDfY35HpMPhvEc6Qz5pM+rEnNq9KbVAcelL2/MmmoGB4JDbibNDjy
duMzPLPUIG2Esvz8CCq5l+kHIFn/yMW2y7QMaBnpblwKu8jzRKNBh6YsR+QhAnrT1LwEuTCZoDp6
ouKWeQ2qdrDZLaBT6/gqM0aFd6jroW6eFbVrT5qp5m1thldz076OQHwXEt17rTNl2T6FT+nY/E2v
Y4xFlOqHUHi9Soov9CIxzwnDvWP8ZjOmGHKy+eDVz9UHlyAF2uJKI/mhgvMjg4wZXBQgcT/sRgKq
DZjNL+hogoi43iOnRVZX10+9S0bVDwQXh06MfZb89BIhmhD8ywEgiWmOFCPFUOVGkV5cqtTdnm99
deQWpnr4by0aS3Ztck5Kc6w0GxY7p0w5erSBl5sRfhX6IpxIb+uj/K5qCZnfEjn3a+GHIWxHbivN
jNPbYMYAg91j+lBMnMSGoyfQ1krVsrUnxhAW0/MBP5wcWZuJbFuSkEAsjA2x29+DMvnIcMu8HTE+
FVpb7HSUrVzW1a7sej2G+LNQoSfH7Yl3IspAPDN6sAnfF8Vr+rCMWX7Gyw+AKJkSgyzKRBIwUpqo
al7RQtuIU3v3XezbBAtILg0bZ8zmAqwALjaEk5CWHvOdXjciY9XhS34RbHbZtYAxSo5tuSEa/YRz
OfFOkvXXoAjnHt3Z+CA/oo1G+kH0NK9IIIRmb8UlIDOrAJRvTq3h8DWCWht2yAUqOpPkRpcuVLY4
vmmK+vG8md4rBfBeK9v2ogaxqSXDZax1UG40OcktuCcAQ88MyCCPLJXZuWeiOlQd+XDGvz5JlAIn
JvEgARWy535I3xQbVhLoFaRnaKNpVrX+cBWMJDAsJguNmdcFv6KAlch3tmFjdirZNcNb3WHfzwa3
7fREDICzdSWgwGmcqsHRwarJb8OiFU19PgcFBmCflxssd2ZZlEt9Taqfx0RT+WEX7zg4KVcy5DkT
efmABokhOUlEX8qJ2hZAuKAVpwNmSDgZc8v6wQ98KUjXt0rTx+W/S2jT/4kdVRSiJqOIghirosj1
l+Y/9wEdDGM1lwXm/kH1Hz9QPno9c2ji/2wz2bEUrmf5AVKudxA5ldUPpADjfbKlf+XFWDtHlSye
musWJ5ZAh9KS+kTe7R54MAnUaHIesj8DSI9S4DiVo+nAG3ueVVpDasJQQS+7vpgwIsoQrwMyybbB
T6VeJEfeDvI01rRAl0rgX6FykgLJvGjQMcka4HJngsu2cdx/pXGytSxGrcWrIQy3G6MBYBBd+iJP
GVxVsPUMRvMFjI/FSzHvLU87GrijLThbdU380dvXjOYP8qWNer5YNMYoeijUcSdHJOjsqq+KKz35
/sv27b+RU7u47bIa6QNjEv/yJ9eBixmgJdl9XNUvKSt7d0z+JFEfK1sGJK7we7LXqTXY+vE7jZVR
ikoiX/oLWFLUHwPeN4Zw2jMwKRFJwoVie2QsrA0jDEt8JXYn93xU+rf1h/WMojAefoVoJ+x+mYxl
5gSv80ttG7MegNVGfrHYxLkx/+gx4BIdspH4C6Sbx8QaYbKQfMgThS62rUTI3wc9UEOZ13Gc3AG7
8Cin7WXpejx9RWj5FK5C5Jr0QcxtrNjNrJb/EevSjp59W9N2RXLgiTX0qRwu12pVvYoIg9xBnTgG
9NxwzSV/LsffFCIciPPtkUxKFZb9LQxjsKsmDyI3NJxLibFBS8WtryS7ombnviCani+LEo1gqgyE
NC1DQtZOGRF9VuZdNpYQceScXqG10x0uDkoBB0+ujfsiFEZ08nYoEHgWkoniZxpi0B8lvKOeAMfH
wDaOSHq0vBCkAgvHHGI25UQ+ef59gsw1iAbFwCw0ia85+3TrXBnlZdxhIjZwQO8pJl5ebMlXr96w
4uJWNRqVtKCe00qAD4D9UzwS0smxbVyE2EhUcCrhf2ikF24CGg4Q66kSQRyUWeKNuWXkYWgZOlqZ
MncXNGT7aaIioGw6dOAoQOGxGfABGNEjTw8KzyYAqSPI8XVuuvRjTqPkMilkVonj7pphwwH5I+lt
cPqARJZhcyBvhXdM0Ud06Od4ys+Qi2wrEd3aD8yzIVRIjjinvjoIPVbAsUTwf5PsuqJv3EcUED+f
5/rq4ydoGn/uImueXfEG6dkx8D/r2Hxh9PsoaX/iOV5JFRVMZfNfMzKmNQ9Bi3AvyxAI49ENfi1k
D0srWM3Qu0hTAQHoSwcFj76fCMAcojf6xaWV2tr19QI5crGwReQRkHyzoFJdEMJCnsO538nlcxr0
BNkR8BbqzXTIWM1G33EkjDH117BXnE8/EzC4AAtAw/U83h1tSmvuBdKlHcm/BoGLCUqv7cf/K2ty
xWyinRsdwl2fOT5bV7F5bDH6obEqx1iOYyNt7lYPlM4TpfStSCSHlhB7WyPYCc20cbgNPkFQEH2F
lzNFNQ4RKfPNKhEkoqYSgL+eAzkOlkGilhzWXZED+JJyRsSpjtEuKIrhQCXn63+Jk5TIT8OvRfV0
7qj93lOO30nG21ZrSzyzMZtfCSY5VfjksRF6AzBTf0oqe5uAYoVwsEKJz6SrsHRTiChSGfWWx65I
qgU9xTsvIUwYtXFZX0guoRfcpMZBFeeOuZPGwQ+0/DzE0lNazFA4KbhuyLRSV85yWvT8q7YweHOI
rkwlxS0a4Z4Xl9xKpT6KaVeUHG1ji4rCJaf8TF0oBGjFs6TV/RtNsQUzjXUR4jzbekmEmTj5IPuN
XVguzQ4eelttNiaV2UrlE4/G4CObBuYubbLNTae+BH8iagrPVXJVmVSzSssVdX8cBn3auQ+i1yXc
tYJ2DLgO2N5wcP/yV7GUqvjIpANj4A+yB1KdbvCDyPsx6RFqiLMmKblQsmIdMO+6KjHaJRmvd87t
EzPJ0UddRmYOToWOAcqCG5Y0Ky8BlVPlMokmY/joObuwyDHb+swU76yXQtTUF6c1zfirUH2gmTuc
aazgewXt8uX0bnRdh+US3S+EW8UnMuT3tOHw9jDDAT+3fQUuM15AgvJEcCRs7yWIEdl7Mq4qB96N
LFu2mS1SL9JVT8pgMEXEHvIaC+tz1tnubPWt0JuFFForzZZiF/qN8odRW9b/MB6xsL1ERsMuo8s1
8l7+bi4qYrPzlufCQjfy+R6kBTQ7W7v9TtoyuiDWE2zMFZwvlaKGgQe8hOlN+80t2CWXj2G1za2Q
yw7AB8Q+nQnh9CzsoFOCYr4epXHxEBgBYZT6GIu0eRAI92sfAIbxaOQErHmqxZkX7aOF7ZNtcP3d
w3Gyte+cHzSZ9ZlijH1gHsej0AZYXBz0lJO4dt92vL5MKrDObaZv7oyREGa77YXZYp3s/3QhcaAD
eqXgdlOSWHSmHMbYxu2BXuacJDt9T7mgeCkt4+FUOSIiNBwRCGv3Gbpk/QlzWeDiop1vEgIN3QcU
v+H1F4xrpYmCgBpbuTzn1BdWA1Gtz+PSs04kO6ea9PFYnbbHhfqAafVUZJ2I5tI8Pm8mrAj8bLcX
F871FDqtKak/jX6tIyvldFJnV6UbfdBHG5lgbbapqW8akZJO/UeJt/F87/xfdLHK+db9dyBwu7O+
if10HQR7x+i9FnxBye35tb/fEelfPajeGUQg+MmoO002YCiRVqFvaK2NAoqALIauly7ynntg1NHE
856DbcmoRO2DBiwO1NTQItDihHPqwrEdPROdGDeRvURhFc2aap4GdTS1LH6W2fzG7OO2TVDPxrjv
MfsVrReipAAR17gYbSCRX4+a/APAn/yt7KLiCqrg4kOsZXS6IACPdllZisgdpRGW/ehiqUj7WWLs
E3qR78Lu+LFERjPI2Bk7ajTeXN+FdaHqzGOvcYh2AiUrkSur70BBByosjffv4ij6kVhGOVDD/mgS
FiQ+40JRdTUyY4PU/qns4E+/KMW7rF0OT6PJvPL7CD/ccxH0ptseZzWxS3pwgxaNYuYUsvMpM/Ja
fWg32Nv8snSUkiklQ67KTcMMsndrYSNc0jg4oxHapLLDDzdJ5nLcrUhUw/Hw89lStJNDR+FBOsP9
EMN9z+ENkaRsmSjzcQflRet/owEQ8aTJm4QGfgn1uk2/sOwBNJ2/OTMtWGq11CoG272gnTCvklDJ
qa65k4QFI324vtLT5zKFCUAmA4wHEUfgQ/8ZB0xwTgZWcyr1kQTH+/Wz8tpCe8GwAZU9PdNRaFm8
i27KOtJqS3YLVF4Qg3RF4hECmBsxuxYUgxrjTm8bdX8x3sbMGoizL/BuImWNTyP1cZiwy6KrQFlT
8CVmuuhD+ArtJNErTfy1z2F+JGK4qCMlFxZd8pCSbDLAmyOxCu2Xg/4gWN2VSZ02rykrQu8LCg96
OTQVfG/+VMKDM0W0j4rGatS96DFXxZVGOp7yHKOCRztFaCzyvhoCp/zpU0JRuqOE9lcnHYvAjA09
lE7eNQCmhJUGOBn0hcRXolL0acf3Gs8a89AdwNEPMAHclUHgVGsLPVeotwzsNFe+YkRl4jKiNVF0
MJMckRuxln37lk6qVBUIKaKDVIJjD4pIny+7M/h2QKVbaURAWRTs3ci6iUl8DN4HUVUz6NdX+BSK
MJgwZqeHv4OhCPwu3Ds+AbB/sHkGlFBASVvyAy1PH4Hzw7Wi/8kWDhT9NQ1x0rldGLqNJwpuzZMj
4D1/LWCiG6idu84bgQEBQmjgem/SRmLfS8LLQmTJ663f5du2v2PG8aTs4Sptz+xY4c3Ks96v3CSs
bj1UdabkRYOZ1jci8GHjxvpmuRd9Xr+TaMik3SsfIkv9Dk2TUEcMn9iHhuuLNpvOX4t4s52GvHuU
QgaxVDQdQaRotNZDyjZsFZU+aXAl7xpWS65mjnsKx3siV8kdERpRqAXAyu1KqAGN70O7wOfMXw9Z
/pXugP1am+uvbchlFfUWqfZWoxaF7ju6278NYHxpbfs9+it/2zaWPsn0BAH0kJx14ETlIKXUIlwg
SADRL8K3bErF/DX+Ey8p6Fjd09cvL+R5xpIMaY/91G7CQ7fi5MAsKy2uE6Ba0/imUwjkQMljRbe+
Vzm8rLg0zOs1UC+zKn+OZ0S3sZyKo0YV1MDuMC8T54BY0DplB6kNwpf6XKGl5cnJ5mx4XzIxbw3c
qVLu7NW8dge9ldDaySoW4bvnmyAzIUqnd742qpHAROyjWyJGfqtSb0vA4KO9y5OdqRGe6P6AN7Pn
EXeLDL8a3L0pWoXPd2feHyGieEDkNEEHK8tzTETOTfngMrXp+2uBraQvqI/jUVmrBiOcuDwwVz7C
dI4fOhgtzLWVCG44n7C2XCTDrheYOAE/KRlODRsjI0I2ZbDSVM1Xai53n8oB6zGejfutqhSMGIbk
55yTQb0IBF2ttsyPKHp3/iX7qUzbrHIMWRix5+MdQt1NTLbsPLM1mJXAgbZDl7IS9OgofDAvrp/l
jJZG6kph2joNcWPcL2Haph4xpyxkz9ATModXWbseIdIxlQhOL1rLeUKMPPLPC0GrfCwkBAVZj4LS
JTKA2m4w8JtVO1NJidHDkwuuo4H4Xo+UTwbh+7IMRUDhfbGGphe7bzZjOu8FUChFzN3c4opiUZBH
0SMIOFGLSmsgBjws9C5GArcnhyUIMcYdvS8WooJh8s6rJqmenAXEWaZRUZSDMYtzuWkYAkZKLOJg
Rk0AQez21qAe6KlvALjD7cVKKlbEi691dwY26+OsV9zGpIFrUYkkwfXMxv1EY9OQOWmWAQRQGFSk
UbeMBZKyfCTx4c9nicxyzheA6M9iliy/Y2oaiwNbv+fHWk2bUx5lHpjC8BwkIfamWFSjbVDx9Bk7
JmTxynXneP2Wo3MjSzzyEfLPb4vdBVLUXl20hHl7e2W5oMbMDJy+AitUc8MGBYwffoyN2fx02QJJ
icgXDVlMiNWn6Te6AHXvkCqBmVjJwXaePTn8FA8Rhe3n7mmqUx6ee9FaJGpoGRpnFs4fnuHccZE8
UG52dkARX0/q4ghi5KK55XQOpDfNiyKT5NTrtdaW7qcQmX3u1a1+42hpMHNsGTWc/3khXsSyPdiN
ec95Q0SZdObhY3jm9DLOycmASzJpmR9uYvv+uitUABaQotP9PwL6WYQw4FtjNqCRWsg0GMfoFei0
+q+tmgcNyb6vt2A6ARNQkJ7N2mmV8vPe8PPcL7wSNEFgj54XRR9cZzLNrduRzIV5oUAlP9HTrJIY
ayQe7G1D+4xiNhVIU6jXr6DiGNC5gvB8EzQxtjtV3FGqXsnbtDpII7yi/BrbL6q1ThNLkMzTlhA6
YTgfq5gxoxmIZBbFTW9w31U01nXrQBYKMRcmMZqR6C0oHjQazoufcAC1eB30AhuRf0Yj7c39e0VF
oN3EOK7/XJbgbeDGxfc2nkm3RGAj+8Cx2KtMmNdG1hxTwvCoIFY/KxRVSg/NKcxXSn9LMH5W8KBT
zlDQ0OeD3AEFNccut4mYHPvK6mU5ZbF8WyYnFmOOFKHAxN+12giU4p5Bemg+nCfgch0l4UDJRmkL
mRW8PeV6NbE6SMSpjf+LcDqdJ5RGOlZv/SM1ZKdGDzFFPdZEvXypg/AlnjgGaornvqSOFA8hRvxM
k/WGzTc4OxI1J09u2tgPFIrSrBsLaOytCE23e0PGfJeZFqQU77/tTjV1B3QLf/qNWvt7X0bJnWYd
9TxgSAOkLKqmzb1UHyJWDhCmP7tZVrtWaLPni5ebGj6xythFPJNXLLyisFuk+eElLOA34L9x/zXY
zjyu8LkzC0UPz+V3iK76HruAVdZ4tlYzF2odNbhy3trQh+urvv3q3Pe2rS39Gzw6dJqG27A8Iu6M
WS2mIYA1ZL7dXxbKGIAmlaD/3/DH6lgTaVldmG3y3ytkFLwE/pSZtFXxMclLV0KqKpnpvkMdEGP+
/hpkdrrebcfalUBNUkrgbpEp97pxM5c4ajrj26+lRt3FuTtYZSwvzY0pJDjITzo442quWkkZ+okY
uI8pJEEELWeW+zemrjb4uT1oFFfZgds1F9biW0AUxxUwopv7FRJJchQnEz/T8aLTXvjROtZK6kla
eYvYTXxGIgv74OBR6zhy1ulJdrJozBfSleJEDIFrHZlhCmWo9WchkAv5zhq9tWgCuOaU/dTrbcmZ
HhoD0detCHStGxBVH09nXI7JS+cPDq+rSkWk2k+ZIArJVM/p/B5D7Uai7Om9ruSdVPZVFroyfJz0
xAt3mD3MXq7kOP0GQcW3YXP9CFpJh8Bltjci68RX5Qps+aZCNhcKHvE+9Rp9Z3mOdvMrJ5Nsol9q
+V3SxCPvGx3mW6ZyrVORRu2ZQdz2Lssi4ur3DWfijKySj9PXcnavTjUfJ2iom1WEzqQDWWhfr1cQ
vF80T74obe59Of9j6MMkVHYt53ZwvXWvT9+5q2aQH8wsteYk7BLHAZOb2mZz+x4g4WkaZakXPBKa
UOClstUSFBMVnoqW0B06+0UhDc4l978FDS1r0fM4BtgnxGXHACsicPbE45ZjaumdXm2CnMyrfXMa
GwbXSbiynTi9fdE6Bl80K16eY/NAjYnLL6QoLR5f7E3ng8QteU0dEDQ/7B3GVEsDe/0FQujh1v1N
RwGDto1Np/8Tz8VRh8M8bcKWIeD8mU5b8Pvr8gJ4MtjLQu3tQIsD5CrXO58AsIWXmrG/iYKB3Svc
ILbbH3fXl8ulIxN3CWTKYeFjxsCy0DIkLYC75mDSXpgLeqI701RmuHuxKvixxr7dsYh5+u4XPLjF
6BjjX9r75lJS4JNI+XyGKRg1tsl0TdtZIyXPXfXLSs2biNzxwCC+UZC2vNPv4RG8aHbeFlWgrpg0
vKxheX5/tIBAzeJfq7ssQC3aDJkx8ife/VtjIb7aNy00ERxKZfwuGTQRlBh8tP7zjh7siv7bU9Xu
+grESQvVZE0Ptle1ixwF0/4q65HcudAMn+370DMtA6K2dv28x9TmfTDkj/jB8BbA2AYKiR9LfxKv
EziSt/FxfmObiCd+/fzIOlJpEkM/uC8Mq+3avne4txXBtBl2sjuVb2RVvhDXoXPpRAVPnRH94s4+
+rUbGbv798DCTaHLt+u4VhGYV/jO8ncYS5saUPbmEhrBpbaa8v4+waEmQ8dC7dmmG/dXgg1RV9my
C5ezTJBbP8CwL/U2QXcLAxxpoERHxFP1fsA0dqBnggI4FHGs8gimaglP1p4a39C4/cV0TspGJ9f6
xBZF0dDp4ySwp+7vzpNFfH3P7BT4TTN5+K+JgepT8JUJIWF0H8uxEnMYLOtBDfimA3nAE6tEo38a
XcoZfgPecNB9S2Q4ozpmYrI0GLIl4aJRj3PkTKmgwlCqBglFR1lCO8dRkSjkFZBnzKzRO4g7WD2Z
I4P7zuuP035i0qc9xh3p1TAcORdSmFSPOKBTXL/g/hrzy6SWj96Xb2R/8eH5lXsk5LX3VTr0LRdx
1Pm9QbCld3o48SsP/41363yyOHHe6CcArO0UleqfoPu9oZxNNdcvTZr9RULJnRClx9lVQNu+45z7
Wd/ThW6nFf3ZCP+/xVQZZrycNm0845i1dkIpIR7xPmCk/jCNO6eS4/1qybGQC84oFRtG3NoufpR6
B5t8CtE4NopDtLtJKlBwCGGNN+24Nbs552Kk67nXskpmPYQbuJUYbtm4bNTdTjyqg/D48U/t59BA
BussH2ok9HYEbYPh9jfxH1bVq0QXRZzbtWdtPE7JVtdhQ1iCJ/hpyR7Y/e7mFwAzkFUnWDYsur2S
K1gdUCHbHuw/LCaafEMfSEwIMmqurQgY/Bs8gZlqjWcgd/cjGp+XNz05iDNZJm9NsDK/FFhZVgLS
8bjADUXLSQJDSMP4BO/wUt1gFm+d6YqBeVB5D4nXUmW4j8QUh7D7+fQYlpl6UzJ5dL4SDEcOsiQy
lrV6trV9owMV68EtOWzncLpIZfFdLm41PUmKITsXvKvznzyqgcn1BN/19whiWFj/e8a1dk16LOPj
DAw3eM1/GQ3JbLQ2QoO659+B06ifRedjUpVr5sbcDL8PDrGCpEFW7y+jUK/xhG+CHcqgyWJwW95l
H2kDluZk4xotFrCeHSMVhSjG8hczcyKk8TV8rTQmunUDOnrxS3ICUcT0/LVXh9n7UPYTV2TVawDp
wsJ932CHLbU8haMTl5jQ9LA3TyQMUDMkmMErzMQ7rTs8XPI08z6EPjVonNBYzw9bLeurSndX6ifB
vWSa/sjRtwRhqI+ozmOGwmzdqBUt8qqJPybR0ThKO1BLtlouM07Fr4XkL2McGXuXurnflDJVLkOY
dPUGgPvDU+NmcWE3gDJ6+sfCFWFhGVnqubByUat7TMPG4ysx1+FACqJlalG5WKt+mh1g1Vwnlm45
xh1EgQ4MwXqtk2Tpcxpv+pbiAZsAYxs8abMzYoUhpTYHCpsNuq9yyT4RlgFtYhMj/Ojnw7Wd9L8v
IhYtMLYFBmGPnlGxTB+xCm5xwrlsOMbqYvRQ0vv5tTqItCZPGWpfDCo0VQqrao+9Kla58PDx253s
5eyoR23bFn9A/0/h8LDw5GJ1yULyOgw1gwuK4BRCXcv3f2WeWzVHM59Iv0x+Mqcq/ELzuNlJtpHP
GDWyvRKBZLeqxKvRragRZbCMwptKU3dFokY0of7RAuU10Q8PwgPaJcjBNJ5EQJx+knHOdnrMD37C
dwppmTQar91wbTVLRXoAsvkBV6LY51LXf8xe35hAZd2ot/EFsVSbqdwNHDO7e053WoqBKICpuoa7
zyHKqR7vaOtmreWDn9eLWkmZWG2Xbj2EHPAIxD7SgaMcavyrnLf5V4+QUoPAf+E7+C102ewSgLmV
rDhdZyZfH5eLLyr939p27IvDPD43CtoIiwZ0oILYLeCfVJd+WTi83xhoCZEH9uQTAADQjaCo0SbU
6Gs1au1eQJYx+cd/DdWy/lYe1mL0AmELroyOfvMBZPoAsuYIDQjTbjuiE5bRvPdqPOzd6AmK7O2+
McVCpR3+d0KPvVyZBF+lrNPb8WumRq42JIP3/uq8U8pdbUkoVZHqFC7vREKsjaPU8lyNkp/d1RJG
fU0IB6nNRzeZOrYO+UjUsMB9cymB1YSEOXxulXw1quQIR9RZ+1dOjwlUjt5Zv+Zauoc3U99jN8IT
WkLjsR8cq5rjYAIKMMUAdwuSH5Tg08le0GYBnqNf4uQbLWTpkmxyOR7Gkoc6oek5tOasYWLNP5VU
r5lEC0IcKTS09gcMNAfoTgQ550tJrHqC4HiD8HC4/MqMLevi0faH8aiP70U3Xn/f5N8WRCXRcn7n
r7p0fq0y6gEoNm1XnJvKo91I0aIRQoy3hFnUVHsMmKOlGaOccBmyWMqyM1D+Vtimbe0ZnyMQ2sx2
zofyjwCi2ArcGvKmBUbCW36N9OAz7RRaHAKRliY5J2rtgeCHBlgl/HBXlpahDRg4RH6el8YbnHkB
o90pGjWSpwCF6Fi+cW8Tsi3U5yNKWxatgJks7LzlGycqvatt61K8AwubXAH5VZe28mXd6MJZyfLt
/0vnepIRdEGSeCxIogJG2hRoqsTEDzxqOBrRJZ9HKIN8zkB3pF0rmhK5DYRZXS7zG+YwSora64ZN
Qrf70LPfFBRfWmFOwN2VSLz8Dwda5K16zD/dkQ35dFKlnk0NrHjr4fRD34zlsOpWNRkmtRohQUaN
Wokff55alFfkMg79RiPEV00DND88csA6CSJWa9jtjhPoF+pCQW4vMRafoz1H7vca9Bfy/dke7RuN
4rjoBS1NBF6yYpsXfpJXzvjzpmOVygaCXyuuZz/D3kbVNp1iDHL3IR9SvqSRCz0ENYFjxknXLEoi
6ot73wgH3nxNSaJww4M2nHAKUJH20ay3iNw/imENLyjT0F4cYUqYwTWq5pzHwQLoGdftEUqsCu3E
uK/nBIIRA46ofkM9egtkajRUhj28TWN+EMdTh8H9R7L7+DQB5v9pXlv0NiILrA3Jd4eYlQTBqrR0
M+vkVhMX7hAM2YF6rtaqXLWPr73sJnpgaaJEeV+Xybfdm+OoITELigZ3hmHwwcN8zav53V9KYX9w
H4ybLiXc7P1v9FxAR7w/gzcXr96OcazZE6XF7CdtTWGmhZYUuq1XK6imW+ZsudxQ0/nzNGF5A/sc
Xf4EkdwR/nUWttA2UFqpz8VeqQHBUDbwRTfXtN1kEQ9ibD1CLkj/lRUswLHEpswxFRukWRqyp3bc
yxGLFo8LorYPsPmLLwBjXhkxnrPDuwZZQ/Ek4kKfltpPJTO4e3IWE7dMBpV898TcB6Z4YavfKztL
h8Xn5i9mJ4NgY9VCNiyGf5GsTFI5AKl3PnS3cOtLiremVpeZk4/bdhfSc01r7BUqYQ4i0VVxi+Ao
VyY0i8grCRGa5GJIoNxWWggUmBNqH6Q9uqNHmGFGHROQTMROj6Ar7ePiWILMC7QFjLO4B1LCFtMA
GlpojBTSvv2+LwFeaDJacHK2uDnYfKF7Im6rJ+8CgdlN5LKuf/BONbzIxMGyuNUSuEbk4tlOex6m
bE2dkz0DZ+lN0AsW7D8+qPrYvG0bCd8gMoRemicT1v00BpOvYW3k2XsjaVUFivQvLfL3SS1fShJu
EUc+BVwhYmRl6zid4i95AXH16yeDZL5uZ0SBshjJ0mbdovNdEwJ08u1hB6kSDRkHDhmVLJRmMFmD
KSrAgm8KLPMWYIa9qnF6BLcDF3U/Zt3DQYCgjNpBxtQqbIvRn7TaHkCMIIH/IP0dKzWEevy94tSZ
qYyASBqwW+pGv5mEffko/LrUzn0vNnoqf8jDMJhchvmGxGaZzsZclFtYgQKKWY6j1WcF21bkoubk
lhQKNsCfUm5DPp+9eBYZuk1djKgvJV/0Y60dFfbutVkHA3VYXTTjUgaBxXThhUNDo37evZYGgVA8
hcyprnFwjPpy3nDL5VRCx+3a7aq8anfUjO6tV4X0PsHD8XGcsOS9pFptuWCaM619bEzT8lOkoKCb
GXLemmP/rnEUTe83gPWr9P+G4Yo4+CNWT7ScxuXVRZySk/ANmLFjf+JLoEBHDp/Bfcf5zEa+1Cgr
sjudWyeophonsJzCAqSZMWRSj/1anSJ2pssXYlF7d/fUeyiWfmAT9K7cMKlBAySZxt7kfohxPZL1
M43cnp1oPXaAeZF9gZVnoBbyBNiVXTI8UREB9wuvjGRdUyCslW2Kn3A8T6ApCX9F63+ycIR+Y7c0
Rfl0XPCFIG+fO5bN9TcgH4z8xyOHqGhWHpBp6qKFkPNEJUwnMy0GV/NeIKu7Iii8RxYlEQT/dIqu
QCpvQUeEp2/EYhXhbwFpKYXU7mzdMtUOXXtocrrY8TmevWwF2Z3Qbmpg/1EtQI0Vsy4gxQysTNWS
rJiwFisO06FobCOhS1AoTua3hxtXLnLhR1MK/RpD6Jiiu+imlQMMbaov/Mf4DEdk1qBovR6NGK9N
DvzBBtFaOLFtjIE+Ah7l/zww1fETScoZUltMpwOqGb+skIvZjCiLMAQLInLzXGnswchTe5e4taFi
pwM/Qi2axJOq/C7P4iDHSAzGqTx49LvIY3qnDG3Qa+x7zRCKGXy6ASGnZ/5878M+JB2QU925HOXj
fZ6pVWShLf+BmH2KYZHp++mRxnwiwsmwNE1HXS1jNp837X0Eg7AxEmu/2Tx39myGqRxWr4MqWhwA
6kXka54ofD3Q9sZCL0+JFBFOUNfmhUt+Yuo1MIEqyV1qhr5Oplw2WJ3nRcg8ijB8++PkpxM1h1tu
JOptpbfKBlrD7zSnxQT82wJ8bs3CdzQhSKniiFFDTKWsBdxutv2aB+286tpowvI+uX2Q1kIcKCxH
bll3fecwFX80x5SFgqsRY40KaCTvLB4OOUR2N6e7MTsaY6QVbgzY8b90w1/TuHmYkfEol4eOXHFH
jdxEH+CljFxYNT9/rR9kiP7lpMotIPQ1pD0F6ABOhjppRemo+quqPlyTtpnfmFE3XFgbE28noyy5
WG+RBckJlpdbvw5o3uXgHOQ0XOWVSab99lLbTu/uKSrnGJ0jt41RDzKpuEY/IgIO3yMVbVwp8gYm
4tlBK3wg8IS7M3cpk2eB5nu9LUSb7YYMiMnWbkaC6GPwzysq6K3OFSyLGhI9D1VWHRZGVEEyXTB2
EfnQbyKYufpKUPHMkyJfARXza1O5qJs5I6lVG+lDAgVMUspOS+IKnvvdaKFGzzM+I0zW8Br33rkJ
YVibxdtxOO+YG+iozHXVYecaMVVGuTEmUB6XnErwKI/tooJ+jw8LfO9CgubygQOV8OKpKcwGBk8C
zeXfbyyQe3Hzjbx/z2SeI5c4FK/4siZ6qsSAmgaMrnPDMnAvOWx40E+9BgxCwn5/0EsyArdIRVPj
yHedfIqE025tsduwH9BORrsU8s3ZjnhuRbXW8Dp0TRsDwVZ6pp9KBmGtNUOp48cpNG8YUCujY/bQ
tq8X3+o67rZQ9Q6bHc2WE1oKRUGEHFX6CLj3cbd/JMYufBsm5E6rnffdm+TNU3WGWnLB499xHsKm
ZpeALzxuGRYFBnw8TPQBunUKbuUsJXlze1IDYlJg5OKky1+GTs219b/nVJr40kz8bVXwv7nUN0dq
W+fhY4/cVOku4fAOp1h+GO7atR/xTwOe7+LuBYIcTpzY8wQc/L29Rpu3KF++d+tGbufXyAX1unWk
JwUOYqiLvQcwbOoYZOi1KCsnC2Mpvbl0kkpc3Xo8IuA7rMQy4FtCN81Di7YRCzW5mYFogzBBtdXp
eq69jE31Dbf0uPqKsXvOaEFJZgTtuGQogaEF9bsT+2TVBE78LfEgndr3a5jVL+QVjNTeYSJC/BwH
mRSbMQUFSYQZlXiDHDYa6QewCBMd3D+ZxdLpV8ycs0b9Q249eU46J0EYoCpkiA6SRSVd8wFR4mrH
NLYK2mf5bdeWqV+sYJptrhg3rNmv3V/1Rsxwt4fY7KKDJ8BtKnt084blgC19uTIkiJ31N/XZhgaw
L66/evBoNXk8PqgWpaLoqkbr/P/ZanH9coNetbgtZQvn2Izq5pJYkViCQ7c35LlXigVzKYnWFiOf
Od0k5A2moaDbtSMAHihWRA33bLpaLqFMod0ZniIpViKJh4dzUIRQRc26jU++Wn5uQnN8PfkHX+Ix
XanjrzlslEDoA8t3H+OwfRtnH3Sf5Xlcx5P0TbIjac+qExg3EnmN+/mANC931XJGGgOA60AGP+ZQ
A7BBuWgJe3b4bdJANbQY8oqGnqSc4tZtuQ8cAlJl0HusTYmLmcAvYwGvUlGN99Bpm28Eyd73Ez4V
YVd19U2j2PUFulvAHaz9aawbCY2HHSA7XfFP1GkxSzLL7WAz4QHU2Ce8l6Ir1xn6iura54CND37a
nMhmMfXzBBeksFANTOnfu40ELFfzl0/Kwlir/EuDCvabU9PIdwbsYT1EcFLbc6nBKtDoSBlO2/sr
E8aAWfa8Wym6XfAeiLG6j6Y7uhiKDjD1Y5CMTqieXDAzxiM4xuivrEG++Z07KRvPdIraOdUJLYvc
A3qsBcY7JFnEJVoXZ8Wnw9RdYz0CuJoKyIESD1FmRLEAk0p49yJpB1odLchc4bLiWKMr8IbmeDvd
zadrweNmAasSV6I4uOEq03DXDQDNbanMz08y2UcFPJMfbXl7LHuJ6s5/Dx9xs1KCVodsieAihbAn
lbQ6iJm3ZykeuR/VlPhPO09hb2mO5MgZ/s5qunjxZhl4FbUhCdvJIB6BFTp5cYJ8lRERTjmDH65d
5qVaqMwSMXoBYdWu4SfygTlxBITQzYBB1BIKL9aBUgHrZPZWUWM6Ykxb0ZTgeLGIJXAHUHfh5Pgy
cICx6RbfGRzGFOa+ztJVL9EPS61k1lPFTwSZ4vSB9+gvwbh+6H+4gMvT43bi3KDEffaQ7EqfPEk2
SaM9EdycIVsH1wDhMyWxDaQd5b9Qfo487j7WlpKKrCGV8N9QF04NTJPkB4+IIabYrhBtrFnQTW0e
vGVx0XYg3LB1NnR3puY5kYSaA8JfMPknt+CMmr1aQbLuoDwAXV9eHNqHOuVg5lBtXJMyqsNaeTuc
d2WsilbyLjgzdv4nyTe6T5cbTrsmKYrunMcoNf+WVfXtNvX5WocpxV/JR7KOftYR/Rz6N3Hh+9N/
wuZUo4TEr3cawEUF13DYS4aHjyOHEeald+Pk7XKh5gdIG+aznqN9I5OTKPkcE8LghbfRIfffFCoi
R3rsV4pxNebxX2APahuc+EfZ6Pb9wMt5IEvfUYXMZgOG+3mSuvVo+9MGk6NFNdqIPjBv5OXQzjXH
acczQpTXArSMjAE+tSKzz8hwu4pohK8obtvBJd0XVYvaDgzB8v2trfgzCpgEa/v9VksDA0A8+55F
EqcAiBtVHWd+cMH8cwDSNrnarBJGAyfB3452krXu/zmPBj+exeHDeuQeRnxOEIBF6HZMkhBs1XfB
kPWBZk/qB3lVleR8ddohr+6tAytwrjrMCL7GenUKAWWoIWMkiBHAdUsw+IUh5JJlVM9pKA9WiUZM
VHSEC82ufbiRUtiERz842Phc/tuv5GEhZtr2QbtMyJnq7RzP1W03A/s6IHXVIo8EhT5LkAhqTqRR
YpgPVNVqt5ANoiqFVuiv+jEayyiqTgJjR9hqE+Om+aUJInHOC7dUDWGIeDttRMmg9nFTgKI+BBrq
OTuEUfHVCi4qNopG8+/O8c/yT8Dxz9Tj9dDZt1B74zw9QtuLrO3r37ZmUJVb8fY6BDYOSKy+x2wN
DjO/cLNyP3Enq5cRlj5XWT98oWf0/QughZNnv2jxxHsHtIZJLiDG7sV0uau9q+JJxiYh5RIsrVIz
LZkGyfY0J+d3YVe7tpPXUPx8ArymR38d2Ox33Lka996HbGqjB8t9TaaRMq2JrES5Pb3E0ZhczdbG
fQ1b6TxMhVoFzWX0MVZ4f+8b7ffpa4mJs5JCFARHt+UUQIdZuoYUpRXfdKQPi3cgXsB5iv3Y/YFq
8ZZDCg1kknONwIllOUK7Y4p0S+QqK5q5zEbmFGwil64SujvkFGT/NgPUC3Lsif4GiBc3fJhCpOkA
lQ9Z22loepgit8NUCAtwXHMB49Cy/bJdJ9MkBVWThyDxO12xxsOCVUHtmD1ffbqQyvCL8lHFd6Lk
npgdDP+KLfG6sFkVSZN4Hm0yMJN+61FMDDe846wUsXBYauFXOXnfgUNDXsXug6vup2c3JtFeVG6L
7jzMJdZoKAH78532ars01QpmxtebRkxg8XukyIeUGQmFOuAyELQNx+TWeShnMvUHGcUlQyqgt9/F
dvOKRwp0PjrxFAjOL5irUvYMK2AfSB6whgyqEFIxsuNACGOwgwDYhBxQkfhjKqJhwYH3ZoKPetV8
qpUbY54M2DKJv6pgGLSWGFc74o7u6DE4FZFvRQkJQaf0oFxj2SNLVXJ/4bJj2GlUZPG/JaCmbp73
5qSwjaxXozh/PCup/Bid9vgXN3kytH8JHMeaXAoPa3AgANozLxQpjcTPc1VuWnRp4AHGdizpkx5f
xxred4oteO28j4E9vmVKnlO/xnzNq6uUJTlOfbfZldqR8fSCf3oGrNlKBpQEcsJ87yq2Losa4AFP
jlfISNnui8EtbOXOuMfneMMP1ltZokkBS1rHEUG7IrWNZHDfEsLb5q09yh//hefz4U/0vSXOhWZz
qhB9ir59x9dYstK/Mw4x0y5GjGwQ9mIIsVV3DuVZAfdj7xsAprTmIpHw+fVA0eCWpGK5OvDEnEAL
V0t5ngdOy5g4EXGtsLdbOW+Gab0OQYwROPtCMHXHdfkoJMYH4cXajo6yg0TCFDfVUwegYrCFqdSb
/i4l+qnwGqRsa/sgDI96JlAnBbrI7qPGDtOSMsuHeKZ76gA2B/plb5JaJWCikVn/jZeQbTtnhetz
BNpPhuwVB0WGfAuT92hXgukFNDb6VYzE6cc+FLDwrB8ufsoQNuDFUH36fOdfzHgHA8yV0DqMbKCe
Vu9M0hIPnQOzyqX0g18tPnllrTOaBIi/64GM490FKXlzlxhdLNEs7okqVNtSQPxKm/GfUzUqIIMH
1JmiNfiCwCeo9+QuHjlPF3uDCZb7RsSzfE2GK0EBkqOZafwIrIklcAOfhHEx0WQQV+JXk41n66gw
KekkLHoJBtBp5FC/HeAInLh9wQI1E6cGMYv7/VHV7OT+jaEi5ar8WvufQ3F5Znx13BZlYxwCK9or
cA4dkQiA1qtSIIwSMFmfuBOkFSzCPbta341lGpncPtF3SW5HSrofNippoJmpuvghbGmg8hlOIrjB
uVGhlCsXPUurHZ6mMvR6h4y45WCyA91iSu6/3c8gl8OfqEio0i5HYm6cVGGrL4TesgbfiBQs0Y7X
pZFIv8wdxs8NkLzlQz6dw5KWOH5c7yndBUkSw+u+CfTf6G6DN255m64YKwjoQeIawQ1RGJGiapk5
2qUzz1IdDYBkI1XYaX/DPFBGPZyQ2rA3sEBwLWjjWClfXcp7VFELLnD41lZY8VwiIB+9bz2SufSt
IScnewxaoU5FixW5p2NVzFtE6scSebq+VzEKcQJkUX5sgIoFxiBeU0CGsYg3DyoeYf4pUxh0kxj/
UCm4VQmVSS/C422GJPMUJsf/Woklsi14ipqs1qzFELRL01QxhI2BSDfr0GzQ9z+rQ3d2kUyhm0SL
mLZWewJ2AXphtHhsAaaMC9kKQfhdR2u7iYS4z+yV7DoAR43LDRD78wtUF6s+tSzuG7Ch8LOwD+bP
N3qZGgR4jqGqA3Hbdp6XAXv4BvZgENhNHZFcSjf7//TuSdir21byJ8TBs9E3B+7+VkcurMnC48oU
ljrpnJ0/VN+RqfoGG3TS2f7jvTHQuF0c7QuuUsLXwoobM3DEmjU0xuryVne3OGKU/2McEA4UfZ4r
QrUaPHn9kUVPYSpPAsNpwWfS9qaliQ9yIzISlBimq4LT3rLqNpMZkPjx9xT+9ODGyDQx/5AsTM6t
nYNaPDWym6a3dh8bh3RinKpiQBkDgHb5MkL1trdL+PNWroi5YKG5mjC5LZ37OD7+v7/MC8xnPkNK
em4WIecYgTZ15IkrFa1fkpzlOz6+IhnoNnMFw3nBSNPKknjj5etWWa3r6j7g+bdv8LKBlW1qd6sd
gQnpv41TSaX6zITQP/bqQsXtq6n6QWUy8WRKEwyWsG6Sq+FohKPV5ozbWc8uwlSDKP0niUeGlmXL
zos6sLj3ox6ZElb9I++qfHi9OE4gcBATl6Rwn2Zc/Z7KvlY/X4ASdodAoVNx6+QWp8xR2noIaNAs
ZGWT9whi0EDeueY7IEDGIMuqpJynDM2fYoCK8isDYN+ACCE7Sk+md7chcw77DPoRKQMvGJeNoKgh
e9f3lhhoaybAlKoAqWzEQes3ZLt0KhtV/nYgHVOCjDwXQCVgmOrwBhu3Q0RWU+KfGfnny7BIb4FX
dhHPm8z6Jb3uTJDGNjDk/x1MTBTKLhpnpLK8EP8XdNf/suWLd6xEe6tjA7SP6Zl1B4QaQQTVN56b
I4j79I3DMkcfw9w8sgNCdQfWMi86/EwUAMLglzNtXA3dlQWrOOKTbiyvFODGqi5FZKA/PT+a25DR
hJvWIYRCGikHqPc477ULNAAbENx5nhy1TBvLdrn4PgiV9sW3zJo9qTnENDGxgmh2pIEwIjrnki4x
WtMMVGdEDFajZbD56+BbsKrlp4k0raMVrrEn4CzAZR74PWaMAilqyuDXuGeRU2kLMM8Eo0C9uJrM
k/0wJB+gSNMzLb+NqfghGdakRqhw1WFCeSThKhMRquW83iTRg2QgS+EhFbD+yUi1zzLffApJKyh3
OyF6RfE1IbBM8c30rjv4whBVK+Hc5xt5hT+uGPbCI/t7dHGvSNi7iy3XKz8QeO8Ry2dav0xYltcA
yq6AfQCqu7jgsRV0BvuOMWaxnzbOELOtixKfz5FLeDdJHyonD3r8tlpjhpzVXSj0M3rfMJDKfKld
/P1UL5jf2TG1q7pBOXKFz5KvQ+kJ9MZa3oX9lMaz4YDoEKfsBi6Xl7XHJr5kF1OJXUAZvr82JbD2
AOziGuvwyTmI5PZaxhguvnYXaNq+Ppna72jSIOdqXCQmBa6LGVbfo1RenPJlK15K5jfMgO+Uz9a6
xPFQ4HdSN7XTkgySONVFL/0692h2okziTl5bL1NRaeuFeMvtcBY3I+qlUY1nN/vGLYFrUKe5081T
KK4J8JaXYd8FICvFFH5itMGj3GZ1sRwFTb3U0YquvdgpnJF2GoVnAUWY1YlqoeHOGFE2Tabe+mO7
8Pm+q4wqnNBBvIJOUpahvGyaCDAbr3z9bAWL9i+lOZ4uLcXoH9MnfRZlo6Pgv6o2s7LIDtBl869t
eZ0avb0EeAeZap/aK8rRATl+/CGkDwchTxY5cEbinCEV9pkILILDlMdy38moLXYfuB4uP6Ca4XS2
qwyY/EGQwEtaDTkj4HZMpycAxCFXOKYB7fyR0r5Ar7DFAjVyC/r7oti8HVumE1fnw1+DB+A4tRI3
BOouH0igDXSXB3WlzTuR9sPV4qZUzYhsQ8Uf1gxJL9xer/KQ7ksXpHw4AImJkkdL1y8Yq/gFzw29
w+zZZySD6pRag6rGR2ZeMaCDQczCDgQuSs/Lb7dB8AxrYY4AsOXux50n6RKX1mPQn74+DB+hFETD
eDHyC+QWgmy/GfGN1qWuxITaq7Wk1aHahR0OWBSG9K71koba21CcUY7qFTLdUMf6IhBIeuXXud7h
Cr5lwWq2HFgZqRBTYDZaUncgFQ0bfAJvUWWswR5CVrooIdL765D67UVD2LBwrUQoAV43O9fS2ydO
U+3cS5sjWqY7bYTqXK4lyC4eEilwtkJ4db8of6bYxpeclMyK7ulep8+kM5i3Ut7AGx32oIcEtGQ3
HZhPE5Dn3OEZ87Z1E7VpvnUtJQbufGmAz47JtGkQkf/N3kyOr+o6QYH6mBu5z7HIXKOtCK26+7JF
l3YP5uC4cj5QyZghG8N04iFPKOegeGWK7u1HSZekqgz7ljFIQjFWp3sk3Uaw6LzEG7shwSywbcgv
SYw6ZW702VsxSJAO+OtLcJcqg8iqnHP7MU65pRTs4yUb+W97lmpORHTHRSzBef2PA+Df4lsEx61Q
/9KTzESEqfdZeh5rD10hM9Jd/ytHTg3EUJRub6fhtacasK96DWm+GE+ysxS6jAQe/0G7DbVBVBeY
mQ93mFRpaNV/z96eKLZiHfcTSFbCO2gxN9wN0GMDqUoqs0Y0FYlHF8q6HXLIZpISRCnJoJEjbtiq
IqmoTh61BMKQbHNvyJ64R7UhIolouAw2zMR3HtfaPEE2TdHjuL5KZsO73u1d7lfPJGbiil5m0yqX
2GfcQhLpE7sTJ0Azjzkh+lSlcEzdm+raZevYmGNB7DQfRKz6+I77RwSvPG8Ev97oObjkkk0AGN8/
vR7Sv/8WJdZJs3nWt4m6hm5H9pmk/RPYwyUiXZ0wfxRvZpUEksiYdI8l7mOSWiyyax7/a76ewp2z
+173EwsXts7Zka8jiUKrwyqWTg1pyLLMHeND1XvA45CnBPxiwshgDYEAoPYJri3oaDtJ0ib1oGl3
EIBzGA0fOp+CClSaRVUo+ZDjF75lAAAQx/t6xRi7408kOnD5Vn/Kb+mnufLDffkV2fugQBcNQJ7n
e76vL3a7Nh3yvYjjHRG+yvC53xxxKRBxRSoQokNv2AgwBKcVtX/B1dVZEvecO5nqzag+Kt3JJvel
MEjYW7ODVnW/PKUCovuFCYkfxJE8jJwQCy21na+p6ln+/1c5zi4y6UHF52aQMaSv1BmR8wO3PCBZ
Q8JGazqu+g3czexoQIKnoWQQJoL2rpYrcK9T3Zyq3bzXzdhV3tzzE8J8HM46Nio97D+E/8uwNOTz
HouQ/apO7t4TNJy/TcLtveU+MrJSaen8hcqzzEsThfbFkmH6HYjYvRXqkI3j73U8+7WwKX3qi2NB
r3GtAS5Ektq0y5lyC/8uzU4xfDz9a6eSSILQVgrsehtYQvcahSdWYgr0beByzzN13fYbVHS3Mc7u
dIGuKhLEh2KmzQ+o0QktnJh47yhPWb9pAapb9SUDVWbJEOATvQbOKKdZhzXPNDe7Ft717epdbpaj
anOnIJS+r+1Sza/Mgp1F4GrO1VQKFkKPPrEB4GrxDh7KqqkkUXwa6/IxF7Ud16Bn/Sfj7DSGn0Zq
MPRtlezBzm/VXwVCkYM1ndchVtED+h2wpu88QWh6NlDWP74wDRKDw6gq68QEdMmbi4VqVvfHf/sl
OmHlbrT4w9eOiwRJADsM0LZAGbyBDYQXf9LxikTpEUJWW8winpJv0gHp87NBKq6i+j06UyD+8tMC
bvTav0ql1ytJQPKJ6jl2h+YTcVl48phERLQ8MQf+AR6FgDKVvXhHikz0fA/iddLYIckX0dJxKJlF
b79LnJkFdfArFHx0Xart2k+lQRnV2wr09OhLmdlBldvoG85CEPXmQ4APt+fAA8qRm5B0aDHDt/gB
vrJRdj6jVDFdQrANrY+0iPePufIocr37i6metbzgpyv35xJpAHYLEhzjiE56H6ydQwLtahijdng6
Vdxa4A6HRecYrfsuB7ALZHbKXqdYLvqqrVtHcigP5ibHzV5M8L9JY0DUMwnzkEEu1YyoWMUnJZlE
eVO/jvPSLDcdko5DIIX5tnJi2Bbkw0ctAu7JensORpTcDgpGmdd4tLLmvpj38m2yF3DRyG2QAwWy
CPBNe02BaBNcNHlZW/AJZxKYgyjJVnFlS8WVv67NPNvC8AUsg4gTsuqkF6yUY6cCnph5psIWLz58
AsUuZ22v174SghjFM9qhKAzAFd9etZE3t0ai1kd9wt13yZISUniQBlYDwypLYFVT0SZNt7wFMH8S
21X4FNWgxVOhIQ7yf2/hbvT1rssgAc77uSyY0K+O4OEENZFhytdmqYCmzsxh5Qfd6Wu0TmZtCoj3
2FLSmLrOwO4Qv9R7w3wSjNOEQqeG28IrRc0fcPsNIDpvu4rOTCl8T8Eak9GjIFxPibRrr2ahQqSN
0u2jt1Tu5c0W9/gJ9RY/h/HNkxB/kQiQz785kycoPoPqvOvgKOBNknlXwInCBYKKvU4TaP4b6zaS
DTgY5UacB8ZGqYlezxmGwjoRMxuVhl0NvoDj9nF17JGPx26U5CsRxOKlwe7pBMsHkm5lcZlCmbG1
HAVe7eL7abYzrnkh91CryALlr5Pskvzl0ftUEFrUqU8NCy7GNPYRXHNtsTU5QS6DyYlKc4buBGAR
SXPNHjk81EI17QeIGmEkOM+F5vwwOqfPBREmIQCby8k30JcozYPOjv5nNf0+II6M9Qc312cXkVpV
QlWfV0gvbXF9kRqUYnAUNwmoBSKsMQbDbr40la2r9ikUBa6DbRnXeoQEKfKxcckrrKCt/D+9Y8f0
SuSHFXRz35EL9Udzv2I5XSdDdDmpKMFi5P7wERUWazVvdiLk321MnvzfbrBeLUO9TvUA/VhRwWAt
sBTskGgKKgrbwhYmpmFXxzbl5QSGTa3AJ4dH+0b3LC/UbeCkE4QdznOh9Z1jE3mO1fyMpMNew1Ft
Otv845sRwZX67mZnE9EYJZ1n5/rQADphxgqVAJOEfT2ZB7Jt7985xf6+pzcVLe+U2TepcaySi/fi
ha6x/si35gDPSPYH0wb4qAJZ/S1Z2SFjRMhqsol6D8WccRg30BMfqpFmoxELHOD8St9HII+90I/z
24HmzoGXmYfWtfHTQnmQFwQCzUDXzbX0qcIbos+wiLY6iViroFK7zYgGK/MEq8TVJCnSodwCNxRu
zttnhT47PL7bgk1BLBKqvoXCeTeYYWlkF7x6P+LBN0YAoSoCXJOWF8cot1l3Q5Djhtrgg8Trk/WN
4KBllBuZ8xqE60usa06ZS8IlGpmTt7QnZ2w9Y7qPvqAy1sjzKs9SApayL26RWfwNkUGem8TKKqib
2zFLvfhedV7RbGKg5HjByioNjzw7sYpFBmeznT8BvjJKCgXaL6U0BdswAiB2zoz+pPo67E/cewZS
ucHpc/XbkApXBu/jGiwXv/pjBCDM8wGeEJSXKCS5y4f3BbIY3y9ojU9Tdg3KiMnD9jfstIYRq6T8
0CPgN9fk/Qq5Hi+rIibHQ9NmJ67nuzVwAAsweusPcZC7qeqMW2+4cXn1udFZKWXycILHQK8i+/Zz
pKB726KoWvu6G4myTDszyRjBXCy1X+2KMV+jtOMGzOeVVKT0QU3TnmqLeQ4kX4hpMnKNpNUfmuft
BHO8Bt88MNsFlo41redMRDm6bCnN8wPVckbMC/q7E4wsMIyiPG4ziJzlaJSB2f5/MLmChl4sq3jq
to5q5AaD0spNdmMz93C1GINEXYcedBdS91eZFGOeTJGMSMOPxC+4o4h77hsO0xk00I06lAQlFz2o
W845z1Ie1tHz5/d8fHj8AXje8+cSJ9ckYrj5XQpq38sff9+1TSNYfWNSd7oGRCvCNMu4WA1WaveX
yfmEon/dnpmLHLHJ4sShnHk5siLvlthn1zW8eXxlhZmiuPo9UkJww99QECaym0VleDKvGxyJZy4Z
RvnOmQFJ6b2nN/7rFoZC1skpn/4GwaDP3eaAL7wRZuGl4qd8PPL9E8Fp+kcpPDHeIFkuv3ZkCLYv
cFop0wlCVm3aCftBcKUnCFPed+IodneywZP4rKGpYb2gfBYFwWwPDeOwwOS9pukjt06o28mcQBPH
sJce0DrDLksWFauVIxM6BAE9MctnM9djtm7SXKpClrnLIBZlCeBoqErs6CdyIPnY8g1HkZxUeuhb
DXKpBaVPJ1MhKQ0lIT6GMGaUeOymt9+9zEAoRBwicjDi6J3Iw2B8tSMUtJ+sx8UuMd/HQFEPjlYs
TRHGhAhbBzjU9bmecyo90OJEEDE8JXk0aMw2ab8Ao02XwJS5KnQMC+QAK1+cLZCsYU+uAp8/kWJX
UoQBdNHjWK3uxwghV/v6Kt7dOcGXJHOSOXxIpnVfbwdprAaSHkeLVOWL0Az/Bb80T01d+k3sARjT
BC3pzLs9oKtpY4wOvOR/OLfB5V2xuHcAk2bMQ3l2ZNHIDl3sM6TJ/FCWG0ljKIHYNGoc+aaz+UMT
9WgRvuxkxe+TnK9LiBv9hG2uMdeSjN4CHGM1TuU77U9pVf5bkikjPG4nCeG8q5TPBTEWf2XNxuLn
mMKchSwXmgZzuZcL/5eNrKdhHThbSv9OV/4eH0PxqAY6efNhjJ1oJBkiyDCo//rnZG8sWuH0WSBJ
49/Rd/chLIHxlS53+USV8UI3Mc99zWZMilmbaypHocLXEKY1hiYlBHrH5hELYiq3EJSwlMA3wnSM
qPDobCqMpOmmDhI1xQfx3a54T0mzjf4pIDPu2H/idGzzn/wh/OvxFa2r4XfrchfT/EhkWRD0TWtU
7lsPLVsxgexuw9zgEkam3kblsMxFSzlEqj5W7qBoMtUsScfrR2+ARmneN42kjhDN9gguPNYs0rMH
j3FwfU2nLZaFCNRvpU3mnZ+tGhjITAjcdMLyvpvJBEfH3SqPG8PMEbtH3EKOBwhDFHoDDZmhm93O
EsYNt7DTAQnz9XfskK85v7NF30SfcPnfyIkyM8YJbL4uuPv6RSNddQYzHR637eQTMYU3PM/gtyfw
FoC4W3gws9HS4iFK2R1XwIVKZRuXTOUMF1t8KB9h4vOo6dkEh+QW2kWcirSV7kqxNs2aW4Olpx40
CUpdCxBV71HoE5XHUZDNA+0q980fygTQcujWTRIW0QYGSKMETxLxnHqJZQ8AWMJb/PF7CRBxaO4b
TBY4NSPLrCLCWNNMqve/MTjTYnsKwnCMH+pd74Hbi3DcKlOENWvvVZ5ovavorVIWMI4a2qId1TxP
c+RkdyF81/tr2HcjTQuu/8m8QxRuJ3IQkAlh4vuc8TcSt8+iOIaKfD/R1QCKWlTsm2AqooU/WGjY
RNs+eu1Wka0BZGLuR1C5Z74PVdAgAGtkE8T+r5Y5e0O1Z4ZZclJ9iJ+EekVwhI58vZ1Wy0D8N8/1
MK2JEbDOq+mVDcOrwaVOngs9LxoRcdW0uRmiqtrIxTmG6kIB8TEpVeWCVvpQVEVMT6JKOKm3z4fc
U7WHlM92HTFHkKkan6bMUEaWqOzkyOVjnXI7UEVbHmBUT+JmVtGbq6ige6vjh24aK2Lh4dNLaqqn
PJOIFhwWuT7GW04CWIQNQGcpmyhdhdbISV2ftQHmDPvjdp2vzTMub+wShVJ59F42w5mpO2lg1Nj8
QRMmYldneQVOor/ESHs+9Y6pv0ipWhHqpBsIReAzpRZ40z28YcUYz0qRchxZrljYuUjIIi2YJrIE
EAx+lzlAen/rBbG5g6s+/r9fso+Suji3LFstAMd5MtoMuFnIcq+CvkLkm4ONCNYXkxO7Xq9JV7LD
RcmxgyHStvzPhvgNQfJMqUOXJYgIOir7ch5lqO8SuqHlHdLuXVeesYZFt39HaeEwBU2GqgkNXJO4
OCrwYZ+Q+DMYhUcs8/XcGAjoGYC0PEzJOrz63jGxRsa9ZqBPIR9dKGAfs10uurm44BJCljwNJVCD
F+AisGh+qnVJJE/Y1zl43MML/IGIM8SYFVtTA0TTd/TcvbYsj0Q5epikLrR05MKnSHgUI/hUiRzt
l/dFvxDNzD9vUeGyJbBA5mISenFxOWCRGWLagI19JMKjKcNfkI9oA9g/YUAXWLJpo6DiD0s5KanM
LkCZ+NZsqgWXBBI3UiAdpUZVp+V8VC8T6qizsf5yy5hcCuOydIgmAB/ZiM6StDHEnh0epBGRJ2XG
noTpTOH97icdtp5Ow9Jm0lFfYlKA0erTUERTaVMBBYzrDsv9ijuKzE8ybETwz6pxIJ01syiFaoKb
acrijS4fbaCOGIlGxRzhG+igahVFEHnDc5rA5V6ElBd13BaXsIUYI3mzK3inKOn0de0BzHsEN0UP
rAt/FRaRvFGxi1gLRDF11WRL9xQxYXlOm+Li2uNgmVE+HsqBH95CnfWDcYRuhZWODmoaNLEniZZe
INcaXrnKaQQS4A+g6Mh0Y7GAbmhabBliu76lzZvOFffiVebGWcwAendffUhM+nx6E+Ri2wC3iBQS
vg5UN0ASdm9TBVd44Hugq/pO9E3X20q20huA687qUaT5FEeJHah3F7XPZ5JEP7Kcpu9WAEGTdi9F
mrmb3K5VTEFY58XsuPeUa7lma8cpkqkFkBpkHQH6Xl6vieF1c/7oBQBtJhqz/PhEYUKwWLGkj9IQ
ey6pUf6Ei2QKp1bVaiEXPP3fbkqn6pqP8vCRMqfps4yUWngsYGNhOb4CsGFdWOmHlfpiUAvBoJId
eceffWvZWDnz93DoCTQtZISKnkTUq5Y/gmtXcU0h3LslSYpAHdqRRs5H76vPLMg+Uk5ikM1rJUeZ
3GDJ4Ccn3j9PxHnlwlkSqMRO+0hwGnFxm7zMVIpYBAWvQlKB2IOT9pHeFvnB0CQ2Id4Un9izzebP
2BCeJPbn27+ZUT/surbcVSUdBVWaiY+ALX62ya3ILU+AvJm3uU5lu4YvH/p95bTtvTt81lQN9os6
U10jdQf4d9PrCF5I/PIZ2cQ8Vx4xkKfEE3VejhRAVdBC1/h+JT3b0idv1xfSnyzShVxcjGx7qKTR
RiXq7CYSEk8YGnsWhbgq9Gov7Bc4PYyZJG4F/sIKORtYhex66bEfGXJMPUt0pQAOS2AG/4REvfRY
5VOt31lhgxPCxOwlEumJ5yB/BEoqz1R+lWQz2Qh9m7QXwYCc+8nm6M6ONy50AaeTzxZDCTvCtPPW
MM8nVSg3y5sij+4AZpE/y7iTwKm4KlbHSC8SEI5snqOGMR5GcfxxaC3r6yOMxGV3zhKtejVF+E3G
ZcBUMXGLen8BUIFdvkLuQoqIAGqEZL2jqzBw0EEUosLy8b84lC1bYpo614UXSB4gjBjdGy4L36hZ
iQqC8D53McGeO+amPnD2PXQ7WE7jf1OgAiV0UwgBGmuMtdoh6nLT9VrjpEr3bXMh2gPuVmo4qhUs
Ha1grKukeLMJ3AWgf+W3LZggW+NPzgsUJj4aY8X55z3TmJeNp9iNxObICX/hDLx/49wG5RDbKf0S
Qb2BKJocwP9SjjmEFwkmjRTQ5ZFy5U78vwbiaV8qCgrxdNRpMPLjvz1uNGZamNt1DR2McVwMjE8J
7B5qeMX25av8uM5UQr57K/vGaLleYA4RlwYvtPF2Qw0HxGIigQ6YCmsWhtt4d11Kua5wLbHP9+iF
6vrYFP5ko+CYKCKNUrV6rZ6PiXIZPvMH6ERKfpYWm3pdnT1uU+13+kGSRmExcFSkuvwEH71Ffw07
17Zsu7j8v4FSJ1GsNEmmoJsQFa4cUbS59P3Gj0pGMSgAQoo64Iv7GRHibNwOIjHjC56fK/MUUHYp
S/JpjzIWd2q5lG08jt5TcGtqb1pOswIwSZUa5CzLWNsa7skXW+NwRlt9DGQYKxUk7TlCJJEWAD2Z
iZF4mdrWzyzBdNAV4NdhJnQWls1c4rr5FMgGblt3mPnYHmWlx8pxRprs09RK1H5G1eYhNy1bn2l6
vY7JMf7bWUVgng0yNswHokHKePCJUiKhDqO1OFHlP3tCfGGAOzvvFMdwW6YPJ1uQVCGugeYM42jj
mJv9Vvpt6gAg98uHHAuD6fHMW9UMdZwV3RRc0VmAD9qPtOs9pf6CBPbhvv7i+WRIWYRIlInCT3W9
gzaoHYGqLl4VEuSFiG/32aSQ3cojbngUHNI2E5oeCPMNYfOjfnWVt8FWbg+KA9JPp5kUY6YczVbl
QF++B+TggASTXzkBt2gMkbSAU7cu+Ms/wu2W8RbLhSBu9PVN20yH48AyW7hdLdsiiFxxaRV09YN9
dqG1a7Y6ZaMycsCZCT6QSjh2vt0yL98UFh6Vy1lIGHToYCv7biVSmrSC+zm+BN4HyLaOvBtV5+GV
SpvKSNHL55/KQ8e0wHubtEA76gIxKNNbu+1RgsXgjOB9Ez6W5tHvahqRsd1NJOwKbc8PKi0HeP3C
8EeWsQNRt6fqS9hjMcUvOYwBx0ZlsGvWonAmVz8DiRN8pe1y7eHTP060vo/09Bqh9tqSLzkf7KcM
301RAfiyep5pIJBS1FtFTJ6sJLlP4UvxUFUfhfjLt/WoZMmrjKjzSP+QhI4v5wMam4k9i5yf3XUr
pnkYJW1LoWb6H28zAY8H2Du2yP6CEg4+i7L+a5/zNS7CfdqCMA/+2F8MdyHHln6hzP/+mOX5nuZ/
JK45GF8M6026HfjNLRTJkPtVFFsS1MMlm9SSKmKX0rJ6M8ACs+GvlftenynR+GlclgiDevGKQYkx
/8EBQZ87sWmdAORBjk93ocxyj25aHZIToKNW4eFQucytXRCkJU7mit3KRyOqNU4NGhwYYFA4nPQB
mg7bnroxAS+xe4hhMBp7TuZyDhCket75e7HDDrY/wNftMMTfu6H+GeysQrirWok5T0xBONJ6Juq7
o/CDEmJGVHUvLL3TJpXdrASOYvbK8sj5XviYu4CVlKQ4GGCVGJKBj7KwCsUXUo3+Z6VhFEsC73q1
7EjZvV9rYArMvIjTn4FfZV4EMMroNZw+mJaVQ2aWMBh05a8yLqOSeElxNxmVD4NHyP8P+/B7eEoP
05MC1Ojv/UiEnNAXCz/cMlVNBpYkAkoe6yIwoTHgwMapHjTNSDdMvkRPC14trvcMjHQfJcSN2eZE
dN+YVeJUe1c7gnoeyQIuv3WtBsYYnSYXJQlc4ehK9TY6WajpegyqybNt34ffZX7aONb/7u6a9lEB
xDqoT9YTnznK24K0CzDbAsrU8wzPYIfjr2WbFSg7l3BZP9z38f47RIif5Ks9/gg2EoDx79LCq4Rq
YHf1pybVk6O5pRt76Ngo4M57uRmhfieXSfEqwq2gh2hTEQF+yzGfVBjCnmPqQz19ETCRNmcEvXds
ZpUePEgcuS1c3Aa39GFPS7uF4iA1ZzpO7ld+gAFzDEV9kBavbotuYpKqRVDxEOSm7TAzggF/sRaz
3nO+FDJmVJlTfC4qptBqOdJLMiMWN/bE94pmQDuuPRosj209FgiNBXWs8L0cxQOpfsOIC0K30vGS
cuO+rqq5dmIwM3N3gqdKCvvMqjupP5S1fbgeVfuiZvuL5K/XjH3fxfnNGMgKWSNmQb0ArGh6Harm
YR9F/gKR03/ql2QNn750AlJPeb4zi/Nls80O3VHb7ks54XiMQcNKDV3V0eO7Ig36qmdK02F/W2Nt
C/8uer7U1uS7iYgxJjnvAfEqpZCqFfApcuGtsZzWbzWXZJFkpFcwQwa5/GxrIoQykpwiEEqZomLN
QIiRvJ5wwLRl1p4b1tWOExfIAxvMTPFBT4jW5K/o9si4OOeK/qW9hu6e9U35uVU5KGBztJG/5wZc
Z34adTAMxQJlCdw31akjIm29YXbfMp8Kivyx/zTEP3kQXievFneVd3CDaWUhSJgGYk4fcT1ZylDm
fKs4ucKxeGKVRDZbVOOT+y8Gz2hW8HTjnZQJJo1lfHmPJDwafKXUT/UlbELipMFEmM4MzJb9n6k+
R4Ic85a4/waxHCZIPbaMZX+GHlCl20ysqB7o15NlzO+eS41MHiRa3HBUta7J0Ib4A+rAlzhXW70J
w0RQCI2uZNdCrBgubzM9zkhMlF69aUVjqBMfAxYNSiTw0UZcD+qKYlW+HfyzB4Pxs4d2bkKL8QLS
7HAhUyP/MBlZKEuKkU0mAKLaD3LFDq+xV6iGYPIfwF7SBebfYaC91uND+VBcsjtqTZ5glJc18ram
UQpUVnySba2EwXP0og0BNg6IMDzcLwckdei218vS7qrMV5wKP6sCV81XQA6vJ0gD6zUdKpCAF+wI
WECBWzAOw9Siy78qG8hLBF+nj+WDbczLfb5PeOmTeV7UQAVdiVEK9YQ8aSbfNC2n0ZcFQ4YRExGn
udOm8nBpBLeWxit8Qy1lFtMLC8HblgE6hzF4JtGnnzxSQrymZiJhP3s7alR7qmgCwVJ13BMZ1aIS
UhzGQhgi65fBzNNHm3wCYZLJyrHFaPUs9zAeM9gDAGXzfnX+WpwWZT9NcyUQ+NqkCldOM75sf8Es
dbiavV+wQxif+gnrc0bpI9OI9JESnX858EM707gd1IsNHHS6PahZcKE+RSgEPqNLrsK9t8OUG+wE
LV/Ce0NhmiZ5FvYVtTGMYiOZiayG3Ux/9wOkoR3YxtZJ+03OjwF8cl2XPnpLyAIa+LLuCZAdB6FI
JEnvDHAk57yxMK93TXBioYD00G83Ad/1SLh290UwZN+2KbjOo+TDGCpr69+PpaT4wwMs0sTPVUB/
DUtftpcL1FJmxkTWKKIS/OeO3nttIBS6CXgESpIg+nmDjHaKxANBf6g5WEg35ybFjjv1jqosVC8y
hlREuCAa/PvgVKdphsA4jDr62gLgK2LV4qt2PfUnOtzfOMB8rdgh8UjU1MoMfYOJjgXDECtnRpDV
WAOS69eY3w+zTz61i8tewJnoyDFkuEkru355mC8gp2WbbbkiM1phYWelgTHa4SWwjbMA4w7OM7Yw
AkNy8Y+rtJsoruUZHt037kT+7iBEn4KlAhZ1g0y+l1ur3GzxBUM/idGsM+wpGNX4Iy62tji7Q+fq
UJ6ozBkE1mvnOY5+m/x3mHOtXate6Wdq5d6rQrFyPv6e8OgPVKTLIedO1iQcO9efhFIBdBBcG7T/
D6BPp8lca7f7WK9r0m3qDn2ZDqgk5CC/JVCvuOdd6xzMXcltwuGZDwW+pop/1kBrhIe7+sVhmlFR
GfvC78ZO08/khAaDd8gpUPjrFROohX7g7ofPIl7vNE7TFZ5dOTKFuEWzVxDKP6ONwjI+3mYcu/Ct
03jNnoNvj+zTh9YKssd1IBizoH01u/HjFsrmpmaGqShqqPCmwbDH5DAnx/A9kRVDVj2lHg5+2WFb
BQ1CcA5ZNara2uSBPoEscZROFXy3P8/hSEKJJLnvYQxAS07bqInliMwbzDjx+4IYk3n/2CUd9Ojt
hVD0wh9OFjLoOODDTgyR6WOunnc43zS+UHYFZ6II7WcJoEt+Z8mtTxOR2/U2SzKMXUBHSpP9EaHr
oiY+CKo2iYnZV4c1vWbtghUJR58MMf6cMD1wj88d8MWWAfII/it9mUxhLjfOYTvZNpuzVPRRaAjG
JENAi0OyOIs6+OgeBJMIRuNvttni1ESf7EySYNIfvRXz2AMg8L4KxJ4wl/oVPcmnQm92hxBb66ra
/dv7BrMnmLv5UfB5nrmVUnGov0XbUMUkyuvSRI2ANcZrihzTmT4SiEMm05Gbzi+ON3SS0GNC3ewx
cLBXn5hB6yRL2LSYdjPoxcMul2s7ZXvabobzfT/aVle28sEJ+4fzvlW2Pt1hq3GKK1z9z1qZ/2vC
bH4CijBN5Ly7lJ/1hNLn4ZZ8PaXjmyVJBD3wWsP26C+gb6R9oomBE3NwR8I3dcjSITK9DVAM+pQz
u5V2BAtifQSktdXYUhNzq6MORDRJX5nOzyGqbCJroGR3sUUO/D+eulcNnF0jceVw4MHXDvhzq2Ig
WTTbmBEp6i9wIwt5UVl7C2Zu/va60PvDGbvMT/lVlVmbAGk8OoKM5UQ/iz5EAcfC83H/kX1CpagY
DKuogyp1F0TNsgPm3e9ZmPa80TsDuuVu/gwufDwS9aY7hNmIpiAKfVW7SIcOQFufra9veGghikX+
MK5m8ZnrecxS0YtHotfBP3bXmgmB2WIhJIfWqKhVsQwK7Lz4c3yJTBErFNhvSjd4BxZZsqexyC6u
C42rwGuJ3K//y/oZbMTgXAd/ICzDxtuPB6UyiC/sFbFUHg7WzBMbn10nw4xHxLzp1N8SocbfUPJF
hE+RXBrg7hIKycwUWnMCY+zi3VM1CoqUy84tl7TOWXFcvyxTOS5TSg0nGcoTqCSCLG3DzXmZmwoj
K0mrrs8YCcqoNdirfYLk9VvxDJBoYWQe5bAUtFUZMY37NmWz4JIGdjuI0DEa2BvhPPXrbRsdKEcr
T1hLYfJNntxDqTExkLcYS/9yB5JVk+QvJctKdWTTg2LhJczPOG6Qz5RKzYezyxLNqXq9gbdAjeiD
fj7pub/vndVzVrvaMW7Kt4NSQHS/X1PTtjaJblgHBJfBFPrrCn9u8mN7hVaPeU3oA0l/RkxnnEp6
fQb6A/dwWiGmCt9KYHrFqLNA4/7NJHESNMBmmiobpJfvbF+ke/5dNYFNhY2E/b3thCAUhVDsa3jl
hIhp+nIsvYB9eRX0aY6j5p6D7PQ/2RyI+9yJFK8+LJeHyn74QB5fFJsVg2ceV/r0wNAMykNMwH10
OSuYSbieE5v1EsrWzzh+Bp2DxtDujFAbSno3w2oH8MY9bFuTI4bSv1cFCVlzt1tPYhTPpSgL3SGf
FJGWzdxnhmtIu6IBTO84SCeFseNuOOxf0mzdvOa5kODt7xYfE4FsBsrxuO2vcIBDLz3AuxVtUHxL
+3ua85zqLa+5P74H7oK0jM6srQkYeb3heM8XsixG1GYVcHpFjeSu7Kyx5QYvm3rHkDIONLSJIyuE
23Okt+nIYQO86/fj2nbpBlVX8dYuVSvLrefSJ9Utwy97CxKN5HE2UorEEShIl1LKLfXTtIvIG/J/
y4gZYRv8/0MiPIk6F5yHyB0U+DzlfHUmOuGf0xaHYodfsszUmxuHmo/wKH4S9HeE7+ZDaVF1anNI
SPRi6MX89SarXXpFOF7DIdirvxXjuBWBZdYX4e5sHaEot6ieEURodlHkBNRcv/BZ09ABQQPksg57
5CH5XWevJ9JRiv774nXlmpktVU1p6Em60hfA2Dp+0mQc+G3WuG1VUV+qVPLLGRCwW6T5aWhi1H+K
2YI+/xljvVuckehVJk8SIvc+18au9NfOuaxmbhPAPOYyV3yLfL/POXk70GJqbFtSPqB33Oyg7VNL
nCmqs/Dl2KiMjyTYDQJx9/m5k17j3gaXzydTKC38MISBRwJWXViNDXuzTDWYicxJczTUcBKsDNsz
VqqoPqswMMB+21jYBM6pJk4fUAz7uREi/jmBQRz9D6vnhvqhufDsefv+128LqeYzNa2pj770/COL
YkENDVbkqr2Ru16aV3Vbe/jwzqebXUPuYrDxPY8leRGVvdVdcnQVQG0HEWF7B7HYJXsA/5bcvtiw
ewwHxbLjNrqqZmGqEoiIX/wV9Q6yRhfe9urFgDe/1N/Ha1EaTPr0BYM0KkIlAg07ao4V+Ow8g4SV
UgeMYLJHQgO70KecxgRlcUZfFHdx+YkLwrTz6sNpNMeNJ2Oj7R3RaQRwNfsPylihWQ98N8i9ebR6
DV9xU1nxS4y6P6xa3jBNCx1ZqDeItOPeQjQzVxeKNK8o6h/Jjhq0S7Sho6qn0pL6TvHU5JOVTnMS
AbVPD3/u3ljpExvmjeYYslY5XD8/Ost4yYkvVMyaYGbOuS4gDH/FgdNlb4kLspklbXLcT0q4yy+C
aQkIKYQOZS7bh4RNRoyp6DlApCa4cJfgWl0kZBDtaRoS3VqUVtJmZDj1EraHgrxvzCvO6YpjzRGJ
Lt5957wMgyLe7x2DcrFmpgN3B+qEWxbkxKJN0wIyIOLFzaieaHAzUfBvFvrGT3N+OOT6rv2HVsT+
JqeqdILusE3ZDVdZLTwZOvKNPv6SyJiYm89SMwuIeJHhtZ13wAzjMFQ3iqBV0TkwNjEg3nGpa9Nx
P3Qi5J9zT7zQKVhyD1v/BF2xW48AoDCjEfgatnFkh41c8kWPGPrDRVJOMYWt8UmhiQgyTpRCBmAX
RdEHb+8GehlNEk2IeGrQ6tiyXrgLwDwpoemrqTHk1Mk7jT7DjDQEemQ+/u+rn9VEa6v1OEn1J49h
qGERFRsghQ5GLJo/mxdnTFL2VmX2Jjm9ebVc/Rdqf2Dpup7hEZ/wSDEDDrKFE/uvOLVC+TBmRYnu
3P6Yoma5/LL/QF6Hq9rgj8iaoAb+CYBEfGMJZbqF1+Ri7g3wkdTwq0PAvcM75YFYlDW5+4ApTteU
TXZgPhnx/UPJq/cQzERMPwyHZYUtfzk0jwPdo546qpaW92rapg0G3AGSmOhUyrN+dHfS2IWvlBXO
P5WsBZ6s7fogU2Qqu9dpGGsRUs/KYTgaQEEinzt8GRAJGVFwpMU/4MSGc7rJayymEsT2M6ZMc6Kb
ocTF09znL0/6GBKn4eWDIClS0HGi/5baJ376qRaBbTrULmwpbNgYCaVUR2jnZpRlAhhAx7Z9h6C4
78z+IZEGFSatQmr+1uLi05KuGpRFXCuIGumX8IUTHQMAa+5iFWO+lVewfDpMHHRqpscPwC8w37bH
EkpypUeSFYJYk5yWZl4dseQ3+LFi+PG9DrqH/PJY8nOLTMD64xBMatqW3xkh2GBVtx/M+i2S+a2L
RQdKRdi6Jb+WjN2BTr8H/DE7r8+fEawVvGf9KkNAQBJ9RMjATAjf0kYWXM7ZMi4rGfTXtw0zw1HM
lNYimwlHADk7ebhpT8zvziI6VNYH5bYUIUAvGlmjAU0r/Ncx7f/F2FXH3N2DpVMoS0efi5uD5k5l
0AJLQKMj5WWoEkmGher05O8eJNDzY7MnLoq/vsohBBckKuxgf1yWq8z9pocOWkspxc7yqfDRQ0uA
VQx6Mn2Tu+pnOBSYbBdoQAc0ESnZm3hQi4/BxYxtM/tK8y9bdf0xXnkv23RSol96qFNo7KE1U9TU
tuVYu79lqyTFHs+ogB1DZIScYax3ctEBQzmkN1fQU51GaWdRJLLXg05UXckxOQvE3AfB/sxR1elZ
so1DEAfXrvTeelEgnb08os+HVuGoEBqNpwcl0PtL5CPisqBs92wVzoxAVYycmu8zaYzoL29/AY6M
H9SSMVERnn+N0YcL1IsoZNSNBq4lt08mNNdVqcPFR+0VMxA8wNM5L1rI8aMcXrKZY4LFR20G3qVZ
8GDzf2LwnFLp/QnyeIQs0/w1hZ+hPiIawaCo1/uT4AH/NCJ8NJPXHyLSBOhziUJiv0q09v4FaeF6
x0npJEkYQKjekW2nwQrXjrki9TVF/fMZ8ayFGX4qVIFzvrp+zlanwZVYPh6YhKJdnqF1Zp8yCzOe
qA44B+EHYg5pwi1IR0fpm+W9kPxWoGalsy7x3xtyXhVu5jy6omFjzqxMZS/s1HLZ8ZXuW9oFYIyw
FZOP2kBTLwtFYqu3ji2vsT0jZe8I5DxN1Rx7RY6Ukp2t4j3jlToCH6Iu7+sBBc1KAh6ICs5w9taX
CENfVc6WO3EXZRImxLALEuFH9v7dEXiuSC26/+k6Gwn3Ekc/hZOv9GZ8/aApMlNPJv53udadUROj
KO07iQhWp8Q8pxo7kL0Rmf5TE2g8puhW6C/f3+grjG6MjyCRCDNC3iJDapqlAkPCZarnUTf/CMqp
IhCpcFDJpH2pzF5r2A34ydQSkliGFwLZfLlfoNRl/lUsL9nRUj9+E8yheldloEU9hLCjLaSucky2
YYlw7LshPVC6ebFHbsdTMrFddKTJ7hBR6s8mDETiGTYH5gzjEuLQrn7qsAiTUjhOmL3ghMkAXsdf
szLqrfN6kLSyuvkAS1NqNS3Q/pRR/L0TFTKG28JFkiV6pfIt7hapgTPmxOFO+BJFQM6KddCIFuJP
GRyjNKVTpVgEw8S5UpXaAdhvKa8P5yjdN+VKsi6qq3YnM/9oG8bC4u94tu66DLQ6qZv0Niw1V97f
0q1hh3CmZjDX2t9UimJveG1u92d7/OnGaSjoPSPk8KaRDSFwWKap3CdPhxxRzsNyVK5Ef3Rh48LN
lyGBAEmX4q02dccP1nEish1OOMYJG1yMmHoKqUktWIdUxjqoDPyJvg6CseKjiGB6NUBtnOmfJi8O
OQQhQBvWcGJlLeItDmcWz93zU7GEDgpqrEWb2BYSNGkpvBr/1979G/Cqd8nw4xN9510XaZBHsPvd
mglFyRl31/s4lc+VMVbLnZvhLQ3zXTDkngOcX1FDgwb6t24cjNw+A9x80qqF0m98SLFM3MD4d1on
KcjJyXs3jLwaKbqQLk7/kvrnLzIMvN9h/AcRI2sI81H7RTt56rye+REb6xiTeT64qyS5erKcyKvp
4987VQIb0Hnn8elEErv1BXvk9Y8CzJ5+2sf5Yt0KIIcZ7DcHlnEtBXPVm5g3MeuTDAU9m1W8bjpH
QttmpKlJnrmgFI4mtPBUpYrgg6+dOUwnsvrHJPo+Pnw2aP+b4bptznoOK3OIna9WAUxfevDKL9Pd
0kDfeZgotW4PxlzJQ/qw+SVhGTZuhAUuHiOVRGF38CVF/HothqqQbTA7YwGM2CjTKSOBGp9Vc+Em
dFimXQo2K46xSbapY0W/+qkK0Cf6sORqCzMTrtg3F+0H6NxOxAq6DDdCRrFZX771N7hW8TEin19X
RktfOi8t5wLVz2BSW6xEnIcaF+jkHYHIHOLT5aSuDEy1z/3RJCAbZeE+489WXecV0nqo0BLNbhim
IPg1VHhC5+itui/usSB7ELErUaUPk4Cf8RBMP5qbUJxZR0QTdATAiFssLKBP+aqwh34+3zAjOIHq
tthMZucKnBIxCnMY/Fr/Dysro5Nq93YC1OibvB5LoHI97RwjgT00eCsDEqx34mGlL53IHHf4Y0eQ
8aNeUtpCpvlZ8k+qqCkzplDUnnV1RohlThh/MVfb57R3h0IvaN3DRpin6Rc3uK+XbsuieUJB4O1x
VRZTmBsTlGrtvjGOwEnLH7e63aDCW3S8QldFT5oSPawXg+HlI7f+zs1zmJEcSESt0XIzhjoMeinB
AZBimG0THhL2fu6h8wbGLAjzJvf/gqfutmJFcD/uyclwsPYWtu53rBZO9U7W3sbWuCHDqpxdZdVy
wtef1q1yqvPZy5oe7Wl1lzWzTVO7oLqvM68BwAmyDk0imp6FmO5OWpqvtoN3AcGBF+FRfTsDC02I
948GubHQFQ0fZGPQiN1ONN3C+XM/CfMqi/fcQaHaNLvfagCVL0rqHn1/IwO7WkTULUN9e/npamri
hgfogIJJd+eKC4I6ZkrfdKXGHcLVzCK9jYhHV/SxgiBRQmhlab8G/SLNC6f9RYhfbZ4syJJ3EMBQ
FtYAsLITsYQo7IbQjj+NlLSosbmzrM0BshjxdCy/AHUucy0TnpHvDEABgw/nFNNnA7BYZBr8ScuA
wnOkOPbUwHAIiVRTLkNaZ2fg0EcslQ4rYnIhKXeMdOwsFDomKz+ARXJUlgS9pTUokMf3LrmbGzts
ZpYMyZ/fyQi+tjoDjbXt4B/gVgI6EcM7N7cSa9JP1FbIRIF85tWV4SgpGLPAAF6X+TuLxiVxnSY8
4MOEwyQDbw5CO2Zs09FRNsyYPr1yZHpsAgJQStwhqN8LH9vIFBOoFlPyPXsK6sSx6miY0YESJqg3
MfS3Bw8u3yrxy+ZZ243OdsBF4a4Ni7ANqgydnbq0zc8OijHnV4xunuVCaWkA9VcEdYC4plbb134l
rVELtQztEP6pp0ta630X2/akLm2cb6EzUdOtB39q6wPCGJCiP9JDTzAzLO2jr3xoZV0rH5SPEwoB
tLN/aWnIEHf+UTzoZxwCICd5I8Ysnf3HIIEr5/SDITyw37RPcsBxcNaILNV/ropAaag1Byyl/g6c
u6U3C2pQAHiup5E6oFhll8MRc3Y3X4WF1lNPftzD9XHIdntnrLB9DyTU9Un83nh4q54pQsGN659z
eVEiEf1l8pfLinKx+IijcJtAeEKxwHo+XK+oOel2zqILXT6kkU9X0S6GB2wIJQZxubwIpQxYKCnP
oV27l2jOvBahaG+JjOQPq/whAfqKqwlpY1r4lMHlb/8o2dNGTm7LMh2xuZSgR0aWplbbwlXORcaL
2kWbcEFWTQce5eekhxUHx6j//ubv8E+ZSy7MWCO5eD8OVKzozWF96VoDfbqmuHinoGSqwtRIwENn
OVYPqydleMuGE0Jz/E/++7KyKlwjhgEMU/eiF5gHgD91m9jc7QOaOCUSNJUqaJyhSOWwbp4YUzAf
UhjNBtfi9aHEkTmqaaPCcAxQMCp4LZKvjOepBSrCDVSVhuZkv3A5u6ikzZwULC8fPONP0tQ1tc81
PUdKx93duAjxfYj1flnjwCBTw6NQzgx3DjzLi/adCv5HsPq/KaoCMbK7Am3kKqIrvYR29o8haqRJ
Sbdwinxp7EMYP7XeWwjD5wdikS/WTq8VAQ9gHQtsRF/ARGeGuvzfzGgw1OrfDb+UWy0vm/1O+wAt
kvspoZVzgKCcZb7csGO1AOfvzXNT5ROpcJ2n+Nqo/Yk5clRCCY0j2W5gyypq3J9SpKmJMiqSNrbv
RIiILWvBWk/8EQ1K2OxZDCABSWMX1sog/8i1oRkl48mV2lRCKIMMx6Pifo63wIodL9kOXLB1T3Y0
xTVK4V3209xsByV4aWAVhOUJEgmmsOKvksTBmDbzhghOpQ1btSRQbMrgnQ/L0FQcKM+dVFVEaL10
VJcIf2pPlNHEtAgL++59yxBDxrYBJGz27I4D5Yn3MYKCSWOC0pcpOyZpyFqHKbZYXRJ8JPv61HUX
148mxkT0o7hAyVNpDG0cTx6/ZMKAv/JnBcMY/LVy3SWHyYVy07uyl3BMvvPaHGEOFohDrgZj00tb
Y+xtyTNoWVj4htuD3Wn2lHwqVUUYoTtuDJVQuH2dqwfJcQATUbHRcy8S1EPEp/XrLRoQtprVoZmY
wF4JUjJk+uAt/GbId0oIN/SBf0HLC+NBg5WTZeA2KC3tj75uDmCMwjpQXS6GYn2xrQpXP+ymFT12
RrSO1pSnO0h7bXARc3OnPj0LCHz0wyx0vPqS7pNRc6w0zj+gE0fPShf3d3gtLKeCLNiNJSuE3B9q
WTI0bnkM9RXul4Q4slVTjj6Cb2h5G7O9/5vZFBo2dk8TJyJbpR9efANRaGe4MhpyKmZv8SOCqBiC
2NBelvVEST/CJKFGKNHPYWNGWTEzMkOA/VitEyZmxDOmbPJ5CezFejxBIheSiorMCVuyV07rOxSn
Rot+o4t3cpoBE78e/A94Nbu80XSvCISeMh1YhFcwehdR3OBHX/jttTVQGtBxdNJR15emf3TnVQIk
+1xO0EdpyMVrPJPcSCjKUVx7HNKnC3C1BM4l+timsKqFu0oB89u1i+SkqhPgYbrbiVPQ3HvP1P+V
T/nHXtmKkDsO8ytN2weGTD8UEvFviPs8/CIywm9EbEQiv7Y54lluflbpJVg2n2sxbO8cFBR1xeyg
rTzwQ4E4oy2pPkPbUOdNIEzAuQo3SjhHMcsQELVHsjGJNuikrgzVF5Qda10bPBbijKKCvOlDtnY7
TbCxK3x9wYQ0a4lwD+9yxHP3cd7GLJ2Da7zKK3rk/TB3XGSqMHNinJMoGT5ntLrxQg1GYAS3HlrB
o2Y1ZKUSIL+JFJQ0JS5Bn8Q2A0SgRFCQ8+tBSu9oKYX374TobJuyl06+dg9k1kQbsZCYt0iM4Mou
M15csAql8bwV80VL43Yegt/8mIroaRO4Udhjf9WMZLdXZ7HOXacxeCvZzgaqV7pv6Yr+26bbicDg
sH7DTrER6ykVBsw7JmMCaMlgmNjFKNY8CIC5emhLIdZaIeMcLFnMx/o9ap0KEwMkqVISdt6htQP0
TG+t2e+ChWtguP2UhnZPp56vbkqCAgcqzKHP71feTbk2SaYDcyxu10lhQ4lymlxVfVqQ8uoQ13xn
5LX29nyh5Tg3Vn1GPRDttGvvAc19rakRK1VMSvHNSAgcIlhH+Ll1mDw+QhbJLlIZfgbIiPUlx4N3
lRVie+da/IvffkIiiKR8D6Fqef8wk8XO8lS1RNl9F+/lqNySREQEAaGiCpbtv06tkdfQXT9y4+UZ
Ln4ybLWZMOwffjZclbBeMh4NC152Ed7Sm+JB1wyOKvJIpiuOlxG8iRFvuxulwBevHBJamxAqG962
lVUgUAUe53h07cibnVbv6cNAY6eb8IzxvXUTOtj89FeREUUnCjicFL9d4wOKPXS3iF5eG2jL3hwg
LkGy2mHB+cHkQObBEvrJzJleBjOSRuiC21/il+XNFPXhwFJHJ0lfV5RGWoL6wfF3AP8rzgUUcicK
TNOdvTNpocuSPaqWDS02hJ30amorGm4ct/vUOVhJntqvBgpATHKhJ8+2+LM4kdXLP4jN/lkm3kxO
A5466ZJWva0iIdN9TYvSDeMAx6GPq2qhq6HkajAFUGuAy5VmVLvyxhh5lSLSwei1lTKuKQRBOlnZ
8vuAOsjfGZM8d5bzbMeYOgYbS2ZHjxnjRIP5FqYaI0WTYvL1hINIOO04OUUXKVUwK+zsSUxoDe9G
fa4uEY9JoDqnj4Ph74ciCbhSQh/b2pRZ80FLJ1ZWRhBhtxomNmjjgLvAWi1pRx8zEyMZgN9Ct1tG
ckuXXgBORMxDB8duUHLOhVnqueT0UiNNiX1LMpQWcO29BpxNlQrECU6IzhxKoOEEmbTj40CyQA0L
fiVC5gA7jSRC+QiloU2ULDFA1rSd9ddxOlqBbwkcSnuHGnnDR191PkpkTwuC1aPw9GOP/sDqqKPe
3XcVezV/XAKqckcljO/wL5xPnM+56x2YfhADj9hlbU6CV29ddxgHAj/QHIGRowEaQvloEEO5LyaO
rI0uKGno6LbPy7Pdam9mktDnL3nWmIPWx4Cu6VXs+FOtLrPYrsPnPrstzrRGccNGrKftWFnJFmdP
Uz9SnXL+LDbD7OZCT6mcm9snPko1gMMYD/Os5wBTglpRBXqS67iVZOUxD73XQOXf+auKevtp+EOR
MrP8cj51QdDL427S9MizngjBkH3JM33oPNkV/XS6y0SRta4nAcQwCLwc26j7/pRkUsdHY/8n5hw6
zzsAtxOkEnuKsVjiyAwIUb6/TT9u4OKwyCpOJug6voQ5CSw6ZQ+EnlfHpjbfYYNTHohajAuBVMuB
zVdma1KVtWwqnrXr466MTHTro07a2vLhFE75Q2oFPYshaUHUr6Pow6/yisz/bavhvOdB3JMr+w1n
wCymwewnx7UxGO2POn/UjeaeYMg2w8+fMvydjbUbEnOTZBMQml1h2Clr9jLVYMq9SR65bOu6OOF9
LrDi39JUI699xXyOeFqgTPZpo3RDIIesQTB7EJy4NbXpDYURKcOBHSZdWOIjJEu3AesaWlOwwDL/
hn+WdU4r9uux7scKoK02AqX0VkKkfCzRcWO8MtAqV+Dx5w5+k1O/9vKT7VEfFK6pUgxVWWKPyqCF
eHJfZiwUSC3PTn3aGNWf7IzTGksl/XFuRxsODC9O+BiPExwljhKWJzIEmSylCOKsSbNipxRuPVaC
RJXXe7iFeA2cppjKEiUXjEawws51rzhPAOAf0w1oh9r5+9aIOVLR28g+OJnCiU4iKyQEyYQsGH7P
MMIWLjTr/IGJEdLvHq7Xdq2SuK3ccBmLBoRK17Uh/m/DluL7CcmrfK5BARbCIK6Wfw5ZVqMjfm+F
4Sh3jAhie5pm1pj1K4gVH1k1Dd+d0XzzqNZDR/j0cXaYWT957CzANU9/OOmLPN7lQneHFItMer8s
sDBK7Zb/CAX86xzdYdL7075NcsAVqsGOVgCrL7IVs9ceuns357bNWykf74qPNZrNFJNGDlEXVxuN
4RB1X38j/mkUrl2QB3j4DtTVIy2btvsEMp+5h4rqE0IrtdYCzhUS15StfeRN6ImTF/Poe61q84C9
jXrJHCpOK3DIwiJ4L+C/upycVS1CDThpQ8xZMh5Ih3kWeO+5jh4WQMF0we+krXdMR7P0yqnjw1Qt
zxRne3w/CegSeZ0p1JbeSP7NQ7BkVjnF/MRb1jy3p2WmMIRLAvMzYhp1i2SLIBTk5NnevCvWvwqP
BGepJxXm9CWU9FnuSL7zoEacE/FJjrkZ1NDPYwwlShqVEflxauj6ObDHYfYK9yb3UKFsg+YPAXO1
znB7Ofif4xnsDZTDaWVUR87I/ad1lVQ6/H0PqfUuKyC1aOyK/G83DyFRBQCDJnsKhLqUucrhyjiS
qQjyHuBcBt8nZ1BBWWOppNMIDfCIQzirEQS29QpLgksg9qly93DR83javpqSK12jwv1ut3ux0QBb
tkl4uYwD4s94qpr6oi2KOlmbUwJN8IoxaBD6/6L7rf2XpWoi8ESSq+/sVIpxgztbyjUfilfssT7e
ld6u78u9tpk5nyN9dT0Xdv+4rgM+aLin0qHtQjAzfJ4Yk+hbB7BAfGB1xucI02lFfoKv/z7WULVo
fG0/4GQMBAVSyCIRw+uOEHghUrTI4HIrOA+IabNdAwQK4Qis7c4Bb+du9iV7QeEXVu9f3kOYhqMk
riR3gWMBebHPn94se2Q8aM83dpcBxrEfKhPWclyjethis0C18sz479vgtjLS4O3DULjvpIIjXkKH
9FH4L8GsOccKL8XGubCGyFeTf7TydozXeBd9gF3A96Ei9oh8tJdGu5vpTcl5hkb6k96SyKjCON21
HJM+Zqm6pqYM+hSH0A9Z7y51jo7YXL8rYmAFVKpg73jabAPgxdE40QWLmt4UAZWiQ1v5MiyFrlpn
bmubjIS3p0XHbZYzXNhDL9YH1x0Hgt7xsPZnWnOoimoDyt/BadQyjXRhrB9aytg+iHAkHD6blwWy
XFAnbei7L0sNP1teRQWMBZGFdOuSUL+5xiak7dIk2pGpz2CpPof6NkGcdthGr7ciwRQwvAOsB+L9
VtGeesy/FJ/J7BQEkb3RZbQXDBpkwVu80Ewggw9LpuLhMVKhjwx8t39uidCJLZokQY56Ks8aETo6
x4pV0GZPjcIz8PUH2xzlQ1w4tFcK4wmzMrIsOlYVJT+r+AQppEL6v+sbgMwQDErfqkXxkaip3zfE
FX0ilVgBKjhH0hiDTdaldhz85xmEb0z3877O0joMfCGO8jgJvn88RZs8OtU5MRLxEV38KlV2S5IJ
hIvVhKW/8zb3fR5KNOoKcZSfb0OnQulmD9vtSZya07F/q0oIFziTI1LeR0/iDifY/CTNrs3IKfsG
f4gqcJUjunCrNnovKwIkNT5DepbnprnHFxzN0Ta+LMsSRJ6NPuEoUll/uZER8zXETCtiwOkLUqdI
2Iss0xE9tCYL/cO75uvEuX4eFmRBzjRpBNf5n63bDNP0ENmVMAiSKi7VA7zoKqWj/UCMUEaj3Hny
d2U9mT9H3mjJWk7ZHv5Yt1VnYTpzlCKk6SsdV27bEbvPtWbbuzwkelGbrGZaCTh5Ar/4mL78U0R1
aLe9umq3N9kBu5vAqFZlWQkHO8idSg8Sr6JbmUdX4HD8rBee10Cbrb7vxMr7oa3PmLYmW9x9rOrC
3UULPeSSnFksrj7QoixbNu5vRHlEgDsywF4IyQIOwnRpYDc/V+t36Dy/WBApSoDJGR6oSKjDPRH1
Un+dx+A9GL1fmc3i18yKrWpWKE9l4pTFDMcUTSsaS9q60HKfJUk5FRLcDljZF88uFvsnnVhaJcv/
6uMxESg22paXDzakk8nbL4fUXJjS6RzsYf5Xza8ORvvuEVqv6BBF52azk8kssZ0ttucYZCTkRjNY
6sJU5xEGfcyBgbxTQqEIRDYGP1c+xrgEq2oyXTlb5NMX0fvyDpXfQBKKgWL/j/vWXJR0o8JUk/tq
nHcWXArQxf6QtvlNT9YW+MHDKEQHTYEWuLDxVbcISamibsBuO6I00Q0MA7zvPiFsT430FJ0KqF/Q
WuznSKXiynV2Q19iRuaM4CzAyOiiplFK0dHFXDJfHu4Ccthnp/5eVCBbvRyMAKduoOvDWRyioqMw
Yd5qP7QbS5uNIWJD3Y1cDSgJd61XT20PG3FZd1zhQ9yyuJKdWkikbce+cyEWh01UutXHPkWfck6r
TPWCtz1iIzsefHdftPAIuvuayYO90M8IkR9oZtdkQ9ym8SCBwt1u1o1Hy54/H0rLHOJsqeEko7oY
qz/1Vu+GRzic7/Rkf+dOH3lZ/KtD7VvQX/Jn3MYz14zpPSd4EstmLL3Yuu5NHG6/YDoiVRIQifk4
3mQ5h20jq81RFsdrq9tIEaVz2IoRFFjcEbabRiY1oPAsEIVhYh83m1NsQgDhkcxLFY7DOZTtJ3lB
SmlINrmP/1Pj9buMsSKwHsUhROLrByUG/8cn7ori1QH+ICV1yw08yE2p1UhsOWwxLAlBIdQaKZMm
UUAnftVypLwpZWMam3esn4zVvsWbqFd6u6o9wGmGMEmZcbNlqWu1/ONTyW670aT60u8e3F2+zsVZ
7owsDME7sxl5DVFaHz3DyrQ+SwWVJy0qobaQYyprnp/50msOdMyd2HdTxciShCHHmtVZGSkXdzzG
7xAm7Ivm/LF7rG8aae2yZESJkgQEvuOruUJ3fzh/x8G0xAqobI8hcGtuIjE85R1UVItDDS4Metp3
UMQGqrN02LDTQ2ZhKumacz20BfyZef9xt7BnrPq0KT+/mbVPPVhtDA7k/EmibpvF7CBusTdthCDw
FY2IsCl7shrKUvBSH4gJS9s5mlMD0eKqqnok0BVPElgHJCQhvsyJVXtBiZwXJvCpy9N6c7HL/wmH
DlbUE4k3v7+wwOgiTYU+3obpMY717633d486IO19Od6RHkuZX52XBoUEavTHyCnQujr76zWz6l4A
7haQLfdcOmdoo5oCEjmCFcYBm4Bfxq5KgrMmg3XQQl9j0V9qKKuBebqxVZjj+XV3IOjatHS9Fs3s
qxPh8O0jYolOcJDwFcUGMUggCtb32r4EALevJELiyLE4S8bBYtwH4z80VNqjcz25Jdqn4541yp4H
WlT9PcpOM4nHAHx8ZqHbqQwZGFwXdvkZPKseOkfU5Sc7EOf34z2bGlRgFMzWMSDO/p7To7DnNe7D
1s+mGQt80H4vNuD8topMxvs+bVk/k46Xio2jSXMkNbqGQ5V9Ekp7ukwtfDhHbaPh4PM1zAkbGuWp
k8J1/o+5uPNdEvQSf/mD7CONHc8DAMlR0un0cvWDj4ECFk3zMJqgsdNBYDMxZzIyJHgd9EIZfvBL
GCN79yHeXPEWHpQt0symgx46sYE5mjJerMipb1S1709Ph12gb3SKI7hV93GdTT4E9ioFHsrllZKB
0iAxBiXhr8J3wulOjt0yKTs+MDxaOz+14wYyYAm5HrvpMMZXK1aA/MmaFdv4HBQ53nUUvFllaml7
MjQC7u/GrdVPfN209lKnmQfirAq8ru3F9xyytWj9BjstxcqxlFJlhnUDVPStErN5n0Z8vc68pUhI
ZEmXbCExxxmhQs2frnikbswp62vPdztPANmgIJKVUNTVAMkAfuRX0KAGLxBTdsGABsYzimnvzVdq
OfXz++4guEZxDBr2FcPSzz5HuOVorqRl6baqfzLZ+Ml/z3SNN/WWVG07TNoe1dlLUgdLcZPiPOuo
CCb0ERFN2lhSpP3CE3G4bS+FNW0GMBa1n2eZUV4y7pJH/p0CF5SZ9sdzSPyZp22dS2Yv6GXa7ZFY
SsK1DVEnABesK1Oo/rhSSb4gIIj/mZ6ZY6vZ16zI8GR9vQOhjEDDjEsLjYmdfKZwSh8WybKbByRr
1moQG6OXdKEHsaxzYYnHkyBb8qDA6svk482dSSL4OVbNJ2J4XXBmaRsDIGTxtA+k2/vlAcr2eaI+
bZfoidyyt6/WUFqtVONP9278W/0SQeETaIJJjCIOIyVGDxcxIT0XntFW4kiA0OjQxNPdD7JeJPnO
8vyWSfq15V1ooD4ozkRsRBjzNJWkgG7Fs9IuzbSFX8ufgIyLYlbAJoDOSsmiAVPaifXzRu4CcxkE
r0ZsRYDRBGQbNBwT1qWU7wY4NnvWHnhHUXyIzu8vD/z2go4eLXBjSEH03mmvpk7mTOF449VEGGis
b0oiF1iVMkE+3t8sZ7yxGNYoCCRTfA7qagL913ALzdssPATAHULVsxzM6EQfjGvenXJYbXY58H71
nCInbSMkIDQS3nFLfoYOOP9BqmlhnIN0xDAstdWugYh74Oe6rzvFMZIf+a0jHmVGcSuLq1XRGMvW
co/7ZLrdssuxKhehSMee8tNxuyrXEfGaODyC6+Izx7Pf485IdWEX6auQevn99HhjMQel6SmX+VHW
aRtgPuIyPFu2EKDRBZHaGAMIw4l4KLzwUisiXg9zqa2I1Z/fNfCXasy1+Rfw8VkjBFjcE++gIe84
3s9fwHRO3QmNI+rjzmvxBJwj8DNb+fMKubTwD8R5115/qajOug+LF1EPdm5F8uSWOm2/pMB4S4/w
qwOpik2s2C8mCX+QzZILt83MyNvQgrkcKn/RUh8PxLUBHOdONNSljXTZ9/rrKUb/gqiJr/sfee1Y
T+BgesMlTtSQQdFtvRZ0CvuxETHuCBjYPc8eN4f7cmOfvqo76FNlpe3Gal+Mjl6dr4s29f8wEi4r
lZItLiwHI17/OnVj4Ie+zqRfOLwvhx9HVB9bwHrlzXeLgrUXGwxzmWXYt/3ty/uDaNnEV3c21+Pg
ZkQUQWO+b5pITMwgzDazmV0sJBvlkKkXfvPZ37fvOfaP8eOEWLj5xKoqQANISQ1oIhHw0k0nHJmk
fE0PgCvivjaw/+qz4WehiJxKcScgV5MQL+9auVBSf5crVVI0LX7S7Dr76S5HM977qwck2F+Ws40A
P2RC07yc59KL2SoNtIAj2/R/MqigZwBfl/aeal8pT2g8ihdKen7TsGRBkugO/x9AkHBxZyCghGO+
mX9VHXQaKWMKnM1ewEhhMhELWQpwDdgt/YDHgAZ/52YtvV/SeEaZTVmaml6dClCIwlyyq52UERgJ
3/+8IOKxrz4WT7Wbgmt6KkUHMPs2jQTz+L8PTIFW77qRgrog7Hku5C5bie2p+a5ZI3GC/NnBINij
AwzK3N6A2V+kRjk4W+yKWJLoPeWplfzkbC8a4Hoy53dHnkgpH2Yr10cEVpF1YTLmRhjOSccFlraW
UI31mbzcGtOj9lKK0Bt80SK3IZH+LrWZkc10gN3L887WAwy8HCHepEpotagRQI/XnLeMdkijbajK
f5n/mOhJkwEBcTqVvQmstiI7Ms56NVTP4Te1GmVVUMFh160QkMLkaLYPgycsTCvXYyoNbvokg6IX
n5e3JXGj51JqdGId+GdNOB6azDimCIB7VZOxuWznGjVaNRx0EwJ2xMmAr0AsAhjDzBjNWLePpSJM
tt+6xENwfPntr8G6qbG02sGbEPQYWZowQL89rsWdD4X8VpfiFSSAE9nq9pSnJOCfV42U+MeZCb/A
C5g+LRO3Hr2sGn7RkIFWUExEZG4+h7QbTf+PQ/6fS3tLJpyoRSGx2qmFQY8rmIe1647ZXc63Afnf
/mT72gCe7BwFHhPVc+h0HJJkUctrYwTJKeaC5qg8FomTxNp4I4saccKMHEGRqbW/3lZCPH93CEWr
kDQM/fKXmaU48A7JTtH5dQmZUNFIs9APTG+rQ2zRgbZP+0FokIq7KGCtxKihCUHARvXQz8FX70Si
EBert0JuNd+J5R/oSe66SCq4XCUa7uyATcvn8yfu54l9Yyq+mLQHaK7hcvfmdovmSq+imYYhUe6F
1334WegHZuPl/t0CX8+6+JVPKeDv80wY1wFBVHEtVC23nNvFRCK7k0NF2pwCMLsLcWmaa50aBNzm
xKsGjmOyd258pQVPxjDlkt6nPqOGLO4F8O9P2Cfc4KRYOgnvPKYavTqp+CVcEe8SdTdu19wpefev
OSe1vzR/qs4pf6V4j04gID426xOqpYnyjzn1JLemUm1IOMhVisFlxoJcT/NW69DLo2q6PUwIcWrL
hPwU/ZmcO+8IsjT5sQjrg9gyizHjZxdpvSlOfaiN2d9N0cWYealhyr7CJhkT9dBf1/tuUlr8u2nW
w3XQI8oG5B59uSVaU3tQ79WVgnekzQBxen7bqPRWmONoQtRHQRT0IdyDypuNwADV1IBX3E7CfymR
SL31vYnamP81oecdSbMJyenFNo/dg5dvCZM0GOOTj0mFR7JGlppLkj913bpnPCis4kBv5b7NLCh5
16Q2TE1mj3Lx38fdEazYOuiSAwG8KeMR9T5dDZr4oI70IlFBIbp8EstzlBl/aNqvqSYqSD265Xer
j9N0j6WbnZIkOD1VFYIZ3otoOOWXK0kHDmjYL/rhOl7hme28FDA3OuoLDueq4SWny/vgT0WWHvaG
WX9Psold7KmNS+ibI8KODEoCPMdGXurnYBARiWlHS6u65lPh51rOStg+GvjOaN/tz8Qjiy1BtrLr
UDFk3Ve0hC4JKn3FmyRqYUmYh9ktLSHX5ktH/L+lZQq0hMNKTBDUTc9dtjZsbhcqXyhxuty3qlTg
PoZRqUBXt1Hw1pImlngxw6MHHpNXp3I0pC0a3/8tEmEbU6ufjn+Fp6MPSyX5680TzII/N4fX29ST
4vRNYiL86b+Tby44jFIGeqGn/+lnIu7cQue6E0EDXXSUaZRHgytV1NMgOwx/Gc/nYf75VLnAF5g0
dJjUtgt+DcnCpy7PjWIKzqPEWDmtu6lhk0gqTrlQhzz3smJxdu4V3QrbBkoRcFBYU9CxB3mXaW53
dON/1VKyJ0eg+9ybuSBrXxsR/PkntwFp4eK2I+6nRBBHCLfbLarxQTynqACTp3Dgz8H62FMnKrXE
nhrEFr7QrzZ/i1zXkniAz0I7RTwm/5RIHbrQLTI5osTIiUB6J9C+1+emhfz4yDH4YS4HTUGw/FGb
k6PXblR6L8dLazRVlonhcnf7HSxaHwhtUV5TvOqBW0TqPG6766TYPxituqjYYZILqirfI0RO8ZQQ
4bVu8lzqXt4aeWtKHM8X93Y3M4KzuAmtxnneA4AC6gtAVMMwqcWgnNuaRRkRVHm1J79WMYM2ublQ
cYG1nXeYiXWNf306pBeqn3WfSSRDEi6J3HiSm6U8Drw8wCjdo91Yv2uyXXXN1hy602q1DtKzEt98
/wd23/6hbnu2xSW0Lt3llncqIN5g+GC9wTtGm3IYupBqacp7Prrp9IPPDvs2p/QTZ1GlsgNBgWRA
KDgB+D+5TksyjYU5P8vHr8ZlJU+yHsKZbDOagelgzv/fYM5HPRPv5RxMJoZOhQZqn72DqoI4j6si
aU5L0c00Q1acJtCyhhrlaeyDgDZph6h9ttGJlJZuRd2n74Olpip3foP2nXek3wwBSVjgP0G8oWtY
hKFlS8CQexz99pcehJtSsADP+rQjxDE0u2wGk82jfl67YN0Nfroar8pUOjQivL8LWskp3shAskEJ
dGe1XV9Hr06QIr0HDiAbY4lq/Qd0ZrCe0KKp98DIcXKesyAWAWOaDq5FPNQy90sc556rMoljgeEJ
uY3pOEfBwiy1zRsY6GjxdxPWZ4sixhxlwnj4HDnjgaemTK2uGmZ9DzyhUGwn/qDRcPVW8IDHLjaq
pLOdONrrhGpFcj8+Ep8wasbwIIABTd4i4Pp6X0ZqI2tSwguObGqeh1Bj14mlG7zmu+t8FE+ibQdj
MJr6pwGMzsOQHlq4+rDW6W5eFLS1OeJa4wNkC7LL5su+3pWEEr+3A81E3vKhCWx3hcRwk+tEbzR/
28subaIdqWspj9P1Iv+l6HOZwA1Ex3dPuDPAbNqJE4BXnecV/FFLhWB7cNKHwObeDqo74LKpbI9D
TytLHJhk4U+kWWA4zmNXPicsx+FEys2Fsmi+QlR27eOhpqEr1MCcrZcD/C40kom8lbbbcCgyAcHa
jaXpffzJWx8MvWqUMElxYK7cmQ7xJc5NOUi68P8KllIFUPbwwWjsTLkKvX0sIqgy6IR8/Y8St+xP
JJl2nCVYzz2hTGF+Qi1nEhbqLuplaIofpoU0HvVK57jsAAXhC8IJtkH+FAQjf9DLMl1CF21T1ctj
oBjn01WarcGDtKo3ksJacsPe65EiVH1rxTqNrB4JhifUvOfQpLthSM6gR7/thGpHQwLBTY2LmjVp
aP5Lq4QAjKWInVxLcnWDZ4aUlcgGil2vw8w63tNnml1VNQrObV+nN3mzDIVUzSm7YFjLK9d3pKkZ
Svw9bYIf8OyFZjknIrjvvyk1BzjE63n1lJulqI7QIJ6v+xevK5cyCmbv6DIRSdTkOUhIpq+mP8ze
ju8pM9HyNXKlH7OfghT8NPMwHlPGqSZBMZKP3w7QLmFj/t3LpfuzMbhO0BiDj+7hbp+ejJ1AxEB/
pyUcAqrnJjYjeAud8spJYRxkeaiktGR9Une6wkPA1N/MaavrmUtJQyBViZzd/qMbMG/faKlESBBP
5NAMJFIhju/TpiB7egeMEqe7CPg9H7bF31VvteK0Pv/uNuWLoHStIGv3b19W1BgGwzJEvcnUNZpr
CQjRz3U7EiCPCDtoRiQG1/KqtPz/J05lL5K3NjSNJPPLlWTaRokJavmLDIAxdCT/n2nqcOMs2fZQ
ew2rPV9fsJi2Crq5Gz5K7OqCqoBMiWcy8JeIgrqfH0KVDpH77QPxQOCTNcZrJbwb8EskTIdnIy3z
uTUM0UMKrZHeYAeNcA2qf17M0rbgO+ZQSofWD+pXHciGj8pDt4gL0htCKvcuZVYoI7IPvPpbhKTL
TN85WUJUg3H9yUfONCeY9KP+JH4aQlK3qskqOuaEKmgpknNSnogjE3BC7NJFVUx93X6xLRDtjrij
5CQOlB8lAotzUDrbWtEyuRAwlpSWKjkcHrQu6uCX3wkdFrBhKovUdOGQDaKFiWZJvDRoBpr8FYti
KZJzLkrE06HA1R379kxi5qwrWmta/ryPzc8u5mnGyH4iw1vZlLSnob+mbXmwBXz8R2hfl8myFk0a
WTU2Hp3mVNY6yNB1sPsB0IkSVUfh7pRUSy7iqGsfmFvhLu28jZC3ht1iRraqTz8iCAIvcBTNN+VU
x3ZnAaHH+B1zCkJgjVM5AjpK2raTm4wWGdWFOCCsE9/S4IdaMVuOjFrFpMZe9L2QhfHqbhyyCXPW
b+N+oBbEzcgtizIE+Cu0daYYgkob5qgnerg79hZzcB//LRe4jG6QWsPjb3LT4+HuyIYN6g5auh/z
SlvB+Osto98Y/lyrg1CjcvXSBoWjS5WP5AfgVIOG8Hl+/V7nivqOoWHPSUH+8QWEIIaGIDCOBBBY
jckGDaDDAzwX5+JbVAgaA9yb/El2Rj3RWyhgvw9GaVQke8h6Y4YHAeEOGuzGh1lc283wSU5v/dfl
ub+vCptaqUCz57/KgEhQ8KWYG8dpzrRuEOmlyWujxdytbcTAdJzEm8FpkG0F2XmPjRfVaqA3I70q
GNs1fUpd6NAZJQkhqy8YF6oVth4K/rVzIxQQDoHfe0gwCU/l/pQWMJXkfjhmJqqNrfirn4M2kPwQ
MzTliRfDWkfzdGqnUTv+leg6vIjb/h37vkJTw6gSOEYhcIyWZUywHndIBbMSJ5Io6oyMe+esNEbU
p5AU8GxVRRnlrtFlbExjj64slSaWeZYreChz+4gjItYjbDUj9ISeDQYNQHTRjog6xXMn4Hlh5+XT
EziRw2v4H4Wc+gPYO8BEtVQvd53+YS4lK0DKPUO3prstlRZAQMHw8U9JAQJkhq09Pm8heThoJjtd
eTTByxgutKNvLhEPV5ex2ykcfaezIPhjjg2cUqIAQDR6aEodY9mOErIO3LmnJr1oCMnirRvk582F
0fJwgiJhn4ksLvZJ4P9Gh26p5S5sGNOYItPTSkrDnLFRuWsTG5ux2hta9WxyPZXjTsUgxMb3eAWK
uHLbxveNiXvQmyC4OD2Pz9M/nA8Cruaaps/1wgWa23+30ave0ypACb5UVyh8yoUxW+RxDpox3sc9
V8domWeEmjJWiuIuKhqs8Rb0JdRX9uCC7kwnDOHEceG0kc1xN4hw/QhOA+V+Q+L7Jl3Dsv13nxeT
37eakpZq6KPiQpqRi7U5xnIkPM6nc+ifpvTAgikyuQOvCQDuFocLmUetdxPJmEd++Qdih18KBjsL
dh6XgMX7kofQc2S/fOTkPCwpVoz9FABCmAIE3Ywj85T0b7bHbPQrYkdGABI2+7YUybnPJb3l9jQo
+C/mEA5zaQlFjwN1pD5eRKfVOdRbs3aisEBogcQEKYi2lU3Bz7+XGkJCW9spJX5vukwxg3d0rBRj
8yicnC2UD0N4LF5ATsgJGFCBIGEdGYvBxk6zFYkO9IpC2rjHmMFNrfovpy/JVIeucwVj8fytqE6a
Fm8CnzR9FodoQ72DJwrz3bgUAJSOskMToHG/vWjgEoShsIXUXsQ55kkTcMQgXCDmcvgf+lwMFjy5
7g5qAmIrYD0Tz+KAvGNLz+Vplu93RY4w/1U7+/6x1vskMv3cizwqf3MLuSC3XSIEKKB/yK34KrEB
HeSQhFZq1UughVbaKWOaRj390ed59bJhLCor8VnKjYrDcZbyWKqqPAAV3pB8XgTCyx4fe7d1BNaX
4BHV9MFOtyxCXE8qP5ehKzWR/Byk08VF6FPLGXJfWRkbheVvLHyOcXeDqOoN31hBTjyVLTcydrhS
bllYmBIa5CESLnIbY1oxXiZq6Ve5WSlW5k94xv/5PRmrqBrxfr51Pv4OG4YZdamUMIuoLcW0WAjL
J+u69rBSbD80PQzN8jJKiD9I4+vRNt82g+ABABvrlpVdCrag7xlOP5NTjS2NTvL4Yuso5Zsg7ckO
5b5eRrJxshV/gJE0FSHhnVRo7tr8YxZk05amZvl1GoeSzNUzuaWZrONvj4aacSI815hMBi02yzNU
oqbp6SSYK8MYEsomSaZlD5S8r5w9a7Ie106TdKDzdJzzEgetenPZTl2zgVhk5T6gHh6YvLA2DWi7
GvR0f4c9MZ9W3/MNTUR0OMUZ6MqKA5N9ChoEHHUtG47M5kFZuIIuA0LHid+7vZ88ivqziMv5dtU7
XAeepYuQH/RF/z60q5o2QRVlXqybh1AfwJvtdgZLg0WyEZzxUDLzqFnu1Z4jUUO+GrzTZBYlUihO
szwCYrWR7MIvhWJC0CQe3w8Y9gtbdKWhTHkwyKyDe1mTB1Z9p3Fh6geAxMB9mc46yZmrqd7bjlMQ
oQijDafU29W/sFbZkWrrI8yBebdq5r7IFi8sPVts5qtAUEaSs/SHiQh+U/Oo37aFU1p8h1EneFyD
jPL55eBDkFI/wLLqOJxu5uqHsMSD+RHAc/YMQfsc3Wyv57LLdOUXkDP7Ely7U6GsNyvvTnYdry6B
X9eTUT3xZ0wAOY4VZH+KiFSGeyivd2+ZZacj5NlhYSsD5k92vMWKl413T0e5xjbSJcvXPpFdcSM5
75N0wPvbXSLrg8dnQG6JkYAig42uvftJAlSd691lMlQ8jkMiYH/rD3PDalT4MR9e9Xgv+F/pMYDo
qmIT1/ApHeo/7Q2Dmw8670i9/+AbvK1E/wRTIDqf39OG3DnX2KsPT+y0dF5INqSNAtKneoTFvMnJ
6lQe4jaNWeNlAGwD6lxAYXvqim6EcnSSQ2KrZqGjL8Km+58WtwM+Bjt47EysrFoVu8DZ5XaHY1i5
CHqzQjTr3eRry8xkRJVKUs+jEqrLKTNoiTKjBlr1qYYqwRP6OdWaqPoZIsoJakPwzOWdgVrP9QMj
HkYMvnnrdpdPCgZRdiSrVoi44P9VUM02jfBP1BTm0IcUPhvHOEjGx/I62ZjOeTD9x0PGVzYClEpY
h41tGsjlcY55bsXlCvw1ejA8XxqWrHUASwSwdO+qnWvfHzEyLHY4xN/fRze2mL82lpezDUISZwI3
j0S3639K6l4pIzGhxRP2NsV/wTEa5h7tex7erPXb0MdapMwI69YT6hkXaPoB/oo8TpBwkOq64ml3
nKVgnwpgW6UA2DD8anTbvS0hWO8HSGt4M9UE+uP9P80s/YkraQse5kUlmYbg+FZc2ogZIqgqLQAt
MrQlF36Jwp2LAmAYK30Ga98z0ge/qQbPwIz4o1m/OmAQUh7/UDUxh0JaMix/CugXP4tZTc2u/hHn
Yyki7Q4XgVs+hQVrLvaJOEXuI4Am2KSVCnnSve1WSJ4mOiQKuybHZ3pZqSlanhwHc7mtbOQstQs5
6QlaufrFnTcOgQUrElK0QLeZ197aQWUVjuyzlSNBawWvZRoaALq2M2ZAIoqNKp0DqLZK2w+19nQl
LcUQCaZ6/u4vNo5AYW2FfdYosd3B9P1bQ+6hrYRS+uTTlDddy52hf1qv/pYYmo0+7pCmkNYOHh2/
bLFT4tUy0iPd9hUiBAnBw9ve6+EiHSAxZHk2uoW3NiJGWN2J2xJSwuo6AGCTESCFdDjhuKvCe/rc
bZ/xE4XNCfYtPmgA5OE7uCr0VYfJsGyWXoV/cp35DdZnA/6l7gyGSrjYsIV+3cCHxV+pSUdfbrPi
mQ3tRgZfKrloiRv7D65XgqqA1jKiPHt8O5SecBfPQ9yuNyvNNi/UHE7tnA8bxqp7aNI/X1EKWpsf
xiDITGtRd/XmBdF5+nL3E8bwk4+xCBC2s7C66wS/Hei7qOHjhOZxLVTJ5il1/pdWxomQaHuSrDpp
L/dlgd0BJ00P+xl9HjuSbg1VoTnbmDiE4Ddn0FIyK1q4Mbg1uTm4DDIF13iCfG5Mp2vt8SvWji8q
+F+nR35C1Wiv+NIW9stmGoXMqppPoOzeCZTiApLDQ0voQUU1VLt9wkKq1f2m+E7zrheDa8Rcr1Sm
Bk672a9jPt+ojgMsDp4IdRwH3kNVG9V8nW4zgDiL8FO3IPXEQB1lKVZeA3uwfiDAFTd3kIenUEH6
2HJTVEpNsdPMpQBbv6u38TCxvatBBLOxh4NpVkfaer9n1o7ZVfu2rEyIX++d1ypsesYqxdUBGug2
511nu4uvPHo5WB3bw5bP4EpHVGpA4YKJcMOKYiVYFUAoPnPvyzjssKUKpPIZ1JAQxDvCLuWQNart
ItqwDgXHJmt/opuXp0gceIvjSo8MH3oBKWVUfZv8fbw9xHd3zPgJrMB67Fngk+xwG+ZWcdyWegTh
ED5s/SxAQ7g/HQlMJiAzNncIo40tSTgxlmGyWE4YI6xf+NnUP0I8XJX4xh+ldPTEvv03a3ogsN60
2j/lWz3U39NvG4iZA26lVx0vSSf2gXjWoUFjXl0jeE7li7BEAvYmPsWJbvI6e9ctBNhunWRodsmf
1dzvfFp+V7HnIITY1oo6esvR34c9LIma7nnIB0Q5DKb5Z/fYzaLcFFy7tXhm8JvenSvwiA1Noh9q
uVbvKPkw0Xoi8dH2RFltymEJhO/NcZYnVqeU2zCoNiDrZHZcasSEM5FdaXyN/mk4euqo5bRraZSc
IZ2lU/63YD+4nukzF6Xbil1++pOt7Eh0TYDiDPeDVisTJwovG/Oc0DMNtYdvotTdKqkKD6FujjyF
zova3BIo1DIZm1786ahbuoVvvF2vLOH1hTvc8/TRmFhrNX/zdGXGy9u1wvxq75o4cCsDhp1r78o3
PjhyVSM03C7LKTsL3EoYSksG4TDHV9MUa8mgG/HsiQqibiuqinraWigvmhilNgugYGqWXRa7DLQX
khPrSaoFROuwMvy2QVOEfz3+valmZ7c/ZcbMbs4QOLpRNP1Uq/CGyH99j5PDxBGbm3dt/INuRmtd
gSibvNnxwEKon8+qGTxCPHNbU8/1QK9Nfp0kVQe8sw4zQRBZWNA/GCUnUSJXQgos7fejDsvEXYUa
SFqKdzHxfG3MdP502MEIkAMzyODkB+a/1s7+6P1zQIQsrMWwqZYtOwM5Yr/MVOEPlCf50p4dDaWR
TknNYJaw9BUY6Keh0uaCZRmRx61f2p8PJVJ1VdbTi6s1ypZ2hRoukd3cSqJdVESKYkHUbzSKO2vC
oKWsm2tkYXFPzw7ROv73Cuf9eruMVWuOHqwshOs7siD4gv+du4IxPviBflabxhENrLDdHtD8KDLx
aPcqQUBeUQ3YeCnWGKktoErI36riQvkG69VV9N4Kk6Fe4J5blI17vjT3GFubFW0Il0QbOgeUP3ta
sK41/OCcFvQ7DBOIVPAEPXzCzFrSZs9K4e729lhVtSwCpmuR2qHi/+1qsuq1ztnVubc/+tnS7ldk
WldU4UHvK+OhRmxXpLtlB046Zi7e/6pemDQaP7Xniat4QqSM8SGnudBSAZg80JzPIe/UAZDp/8mq
N6vepfHoNEAdB0V1LqgfvWYJxCHMtmlt/4tMxkk1GCwAl/ERlqr3+Mu1fqocAhCA34XVKpAUUCnV
8GcUCcR3iUxUpJYkShVGHHjCBgDNRmGJ8fAjPZr61SIaJ01ne0ZI7cQThiO2t1t5Y8TT3oRz2E0X
GbbwhyABt6QYQNXRsGRbyciHYhY+0vpGkckwsqPYRzIGsFPeMUzzUV7fWHF5PAggJzAICM/nzPrz
Q6fB8WnKxTYlpd74FGECLEhRJhn0KzzcpPDN/FTYMb8uj1EGbrC6rdDzWwvukbJJn+ssElVoqU7U
mQ7Trq8TyBI/a7NDIev+0znXw7phGqRUhg81w0IsZ5aC3Ehdv6vY2k4sm9YcLHPxvyimphoUI8/N
5hoXOWU13GAeFangk5OIO47uB+o7Ro/UyDyWssBQShyGN05FpsHbSQ594+ansypuQ64IZ+Io79Ag
02o/Bp/NIlt4N+EmKQiW6l012mI7DjBXimWYaS8SUFPv8PfGvgS0bVNuBDNXf8cfQXsqJEOS0COB
8l+SmKOmeFp0/aFaDg7FMPhj0JhTD0KtQqzz9hFYnu5g3HdsUx7aOk5BCa8k3zAn3j5C7JmQGtCd
ulRC0tOMDG/6S1g8CwDX61XxkMZe2Fc7U1CKRlR3w4JlF3FB8KQT/blpp4rp6v7cPCWh0GXF0WIg
0ew4PrdXp4QTT3QRm31XuNKC8feqinKHAf897m/xk5kqgSnImFP1kjRzI8H0E1uEpDgB9RqlC3W3
J20gh8rBaRhGRNjxnxqdGnTExOdgPBVZRzv6aglz6s2d2YRaZrusFICSjxLAmIBxUHC5hdTUbkEE
W8Sqg+P6DPN2eJEQ96H4D06FSra+CwI3M3Oehr5gk/EkHFy063S8kjJ6HA2mifN+GpvgyH/023Xa
L+r7g4aRzJemsf0n7ALypnUdLa72edPeVxn3WCzvaUBH+dqsVfCemtkK5n/kYTWsh9FsMDw6QxUY
hhdzNyftFoB/d6GVlyb06D+8K/hrbQXO5EdxJo2mdrIbnlzvN361+hQNRMVJerATyH7iPjf/vcHy
h0eLqk9W4ZsZIGEUnisRYD5eYyTnx8ovPB2ihOPo6CkVoARh+FHZ8t+DLWO5w621O6HGUV7NoyAp
rBAZWsTC055Q/1M8yL6wYwCK+ewGe6WrA8HrbZCX33xblj0MI4FRUpnCA8e4OzPsCd1tbFsmb48v
DDK80nId0iFW/wO5so6ngY26NRyn9UlrZmAXRCdM+FiIB7se106JdZ7/KNo5B58kJy5QHLSgX2XI
WnVYR5lUR5pYSWAoBkT3CFSOOhAfaVAyUDZDZCIjtyHl/6gjwXC0jZ5eQZCxeIHPeGoFHY5PbrL8
VvcCuIGMvCQD/yh6zCbyJf4CzDRmLN804wnDT7aqa5znhdStKnmbaVjPzxYoxdAPJPWMLmKSynUd
g+VMcDGJWw5tjmbROQp4TnTK/S0EDXdJymTRbdS3FndMTsC4jmvpIhCylxQX2XG5RLCdcH8Ue/Vo
XBNs7p4AyHoGDbYoo8ZkG4rPsqanvA5BEBf1cCw9VwxpWsRMj694UzbY/MN/NBbzFB0DkmzEetNT
aJ/YXu3h9ccz/WQhkzo1rNm5tIFWkLmc4XrHwY1tAKU1yionrUMlubzZiWzN1NCLzlwccnz5S+M+
eioc9lYtU7yuvLgtcqEEzGxx07uqI/tSfnGxMU0OoPt5VTYVEt4OL8UbJ70q0ZGSwIHfvN63QXDh
uoGXxC5McNMRI0zsyVWQ2EXEWIe9i18a0aNINu6TQbQWV3+LkELS5/AE1nd+MacOaHM/bM2BOIkz
FeahiWg2rEY37l/gMpJe77PBYr72cCO8lJtt9VJnzd58x2cgQSOZZ1nXjlAQmHJkudyp1lrrlJXY
h0vyh4jgOqyCkJSvNdIAfhNyCidWUmCbzVPM/o65d16LjFkwGVa3b6nzsi9GCs3dMM4GsZQEwbO1
8nVdBqU9+YJWBJz2pRIW4KgkByuKidH5o9hQKcoakq8ndzO0xTviTB8GwH0tAMYfIny85ieNC1S6
UwWR3+/r025BLkwvoqrK/eGa246oqbriDhNScDXiR7XJTLCqj44Y8FH/S9+eNDo0Y6AOY5y8Gm+W
glbRqr6wvyKdhbY4Ui/6pFvo2IlkcEIJxFEIpV1Ix3PnCFIeJ5t7Mrwr714/CffG5jTM6y/Y9LIm
0DeJ+WCeRjVBv70ldJr75FynFcPp6f9wHxQuG8bxxFbYh4CgtBttBPv2tOfrTtdZVne6KiqMgDe4
uA/9WNGyqGNAMMMi72tWk/OwSkQP4lSwgTanJIHGjXiG4AZKLUSg4+oGeBqc2DpUgvsKXaKYYLDe
4WgtLzNuQfnbKO3PcwGG8ahWIl4KZEMp2Kj/xENATtPAWSDv8I9F7ZC94+t3cI/ER7jUJYf/K1Wm
/pQiE492bClIqu/DvVibwLSH5XTePxOU5i7e++TLz7LDrsEfBmPvqSwRuh2LBTQv/dG4hNK0uF3d
B8BYa+AFVGjNqrSiAfEb8UDwuJlO9k5BcbZDFcGEHhbyRgTBE2OoivWnam6Y1OFCYDEs29ajeGz9
2B6LE+XTft9PoCbKrQXEsez8ZSmb6KnvBFmQRj8ZBlokb7CYkfmR5eNhuNtYkIZIY4E9vGRBcfqj
vYwAek6tSJeY6XxuXlApbLPNNzwTFmYE9ES0vzvThuNcF2TuMwcMgVW5drl6IUbqPpLr/xRy+TKi
0I0mm2Kb6K7oFbO9/lQA0seCYU/HezJsoq6F+0apr5omUaudquP217PnXZ6qPDOSxS7CZ4r1laTE
hDw3LPBQGMW8wAYybuXKfkXUjt+o32X6HScSCldytnKnFfDHFRi3Ct782N0iyR2e7IeISTtRphLJ
XEYq1+5gPHzC1Q2udOj+6Oe4STLNaNOx5XHYw62N0EGR7pNcWzVOuMN2hL9hJ40c4gemxObQ+eXC
IkNpXAGoF+HI3wBhO22otfHClVDVGvRbIJoWoXotJqnf9FeCPvfTsb8CQzfBFpMrJbYH2omt0uC1
RkIR1DsxFAxLNGIgvd9I/00ncsq3Ba59AnoY09lqxMGRi4/29HDXdpRktMpXJUDX29wa1XkiPwJf
KRZj5/QKupzCKUUNPF+qSbZ8kwDe90JKA1ICRzf3iqNomViOSyhCFFn502i8DgPbiZRNdeAGhcbO
DqKvGMLvj7MdC8LGvT3IiqDayZySxzVoqAaMM5wNISJ6IV+0zKlkbyMRdUY0LJxYmTlH2XutzUrC
AqyfXh5Xu3RikLWQMxZ5Ogt7ObWNH6uoZqdQ9viqgZoe1e8Uo7AvzLEgi5NwDFQgaDQ5kjw3kU2g
LPRhta5nl3WZjx4tD1m2ESx5cALpovRXZ+0hF5SvshJTH0AG4Ibw8KFfUGdIpJRNr0BRNWNWzmNX
U5nUmzu0tq4w6d3VKesWLT2TkxaO8eQerQcAJXvG3YbGc3PlPyTvr4otSfojiCCToObVbjgDFwD9
BM4wywyrDnWDb+2oX61Pgi2pW8DjMnqWwwIN7i4wdMUpV1vfBVwtAcMFGKrWrvmg8RHcakVWH26G
+eMBhwL5L9ZVWOaUlPd//t/OZtpH+khCAqkbykTv/Ra3czTavzBbpF8kseDbNuXZdcDRKFP74WWP
F3aze1aUu+VcuaRDWynqyAGUlDhnmJwCpfZUNrSpsax0kOEQPuVRbMIlBLNbs+Bw0cBHPlb8bSTC
Gx2cdOnU4p0NeNE8HzImhRxFZf+KoXG1rqO54fYB4G8XgwXQO/nvSsSOcfKcNEFyKLp1/OZ7u1cP
x7gEJNkEbpS9WFKH2ifbiRfC2jA51qrhmVxee9JgbLYydCmhdfxeL9l35FIPbxbXKWK7VEhBvLXJ
dxW4UvcR0Bc2wsS1COtlYVJ1okTjJEjBgce4QKL8zvIJY57BU2UdXUD1bb0C1qALa1UXmzraxmbA
sBSvh7lSMiWOWAYKARIEM1cebWmnLXzCeEHlHJZjkAi53r/NdvNrwN+19ULXXTixGLj0VI91j0Vz
CfUP6pPEUuR6RqSd5InOo2idOCZtG0OyD4YjPtB+0u73HTy84LK90jnUwt6X8trCO80uCDkbaWO1
oP9Mvt3iXocCcAiDPbi6gIxS/DV7ObHOZK+Wpb/fPhoDhyJ/Ojur8RwUE0fdLYGvOYaeeXye+aCF
lWslGKJ0ycs7Gl250xZkb6168+VW9IzhLX25DzwHrAGLeOR8jKkZ1oKafmNnW9Eu1hzZz0UMQe8Z
9U4pe9GB+ZiMlwqVi+0fP/Jeja7hmEV/JSEcjmeATmUhNoJFABGLb7bneB/YayR7tiJfLhpS4VKG
Fpoj/GgFnJlH9mkh2vJsFA+h0J0ZlPvWaRY5IbhE9wdDH3FCo5K0a7bwnoCXoy+N+ivHj0/WIZB6
KtCx1v/LwhPLHiynrv7pXazPwtzYSD8gmTZNNJyeAihJOMAaCB+wR8F49eXiWbqMXbavHtWouUym
c3OTnncolEvtc6CMBw/TL1EZXKygzl/6bmhgqGy+1K22RrgTOxPoNdYeR4iAjUcCqWOUCSXYSBEu
707vfkTGTPTWgCuJFzwoqX+4yJPnHnv/LWq6vsUmNhDRNzp+t3alFrIjmgiqSoxEZbZk9kT+6PRa
/2Qmc4JtD9lFUE6MLKenyxCxPWAQfyAVda2nFCQZc8vD2QjQGnjdmD5mk6egBP9pC11Q5q60CW8l
TomiGCLE81fDguRhCOYFe6RBM9w2vwZtd9IDshSZ1b4rGuzI3GZm2GExuHXulrEahXoH2lT760VZ
9oIyU+WlNEbV87R0AASi9INWpmuYIsgEid7EO25+hJ04f42vTwZWMMi09hZlvX8+s1DlJeoLIVvg
Cb2mmXGh5P14FAIdiHtSNoJ3S8V5qPN0IYUu92WILIjahx4jn+cI63p4V9yZgjDaUjV56ON6PYyg
1r1rgWa70RxgNA/FBiSTDipp3uCyXw+x3qllgFH0TaR7EJbfK+JggOs5U6j7Sw7ssh6wvVnjA4/k
q+VNQlkCqNw2i+rO0ilw4FlbIsvfPCkA7nlTWTDSKci9ObDINimsh8F4XGCB6UONQxYQRKBi3lRe
Uexiabxj6AkOT+E3jwCrOCOyOJNa+HNCad8yI9w/zH/YtPIHIJ5r84lpISwkErvQQYhvpOvLMZud
0IlaAz9Yrf+1Eeruw8CZQ+UGax9eIGt3ouURLUdu3r6/mI9yzsUWcH7qqZ7HdEbxO/GQ9zw8Cvk/
y7U49/kKl/+X4BETYg5CORGMauq0OOBDbgaTGI1/Z4PxgNkBmywAFT9XPFJ3XZ4KjPvJWKG4+z5W
40gI5l2Y2my8mX+hns9LmFtNe4V3f/+g9/hDDecCIvFU2u/P9DeLDmXfP0sr93XDkIqF9PcYGeKS
K9ViQsftU771lOMfiUY1o9ZH+lwCN/sCtNy6JPh7cEH+Xb6v9uf9d+oMCPoOaHNNvVNYbR+lScCT
7WVgY01euccHGiGj8xJgbk9PbtoEiL7I5YlMV1eGjpaQLUaqcZc8foKTTQpQDP/lb4cH/BpOoj6g
UJvrTlDe1Z2k8w9xc9W/AB9zvlutkAwF/3CuxwLDsRInEk0ELadvHsLdSS99BTCTh1LoS+AT39ua
vEDUWYlUZZ9/9e4L2sYTi07MU5h7J/p3wNHKrZUCplE76J+eE/trhKe0jz/VJGlGSw3Vf6x1uXjT
x2csXRpSkpmmcteJMjo8iyKwR23Ik7+1WHr+VJe8vSFQT6cWdyhggZT+TN5xtOWn6lPc0E3yd8DP
xq0Ylqk2NcRYCl0cI9HLQ5Gl29j8uHdVnBG1TQxdjSvXMAPPqSHavTxqEJNYER6b9mJ9PsWYj5j8
Z0mOEelmOeX7m0/4JRrowSck539cemyDYKikn15Q/pgkG6WoSXJKa0EdeUYcVmE9X1VdAMZUGHP3
JqPTBRkV2ke6uj5fKbus30k7rOqziEp0+7pKx7MX2I3mJDli+9An8pzKyy6Zd4V9VqxKmzddc478
txzCv0s5dy/zrNhGKCHKUxaRknNEHJVNQJxCk42CRY0VnUn7tgaryg/fWELG0V+7ZMg6KjY0WmAn
+RGIIploXXi8OXOODQGca0wKeaYrA6KbUF32qOHIXa+x8cHsaO8L6oCVWKRB+PTLzQAaZkOXM1xi
t+g//Rb7GezZmIADLC0PFHfNutqQGK8IA3zeW1GyCWu7tgGg9SCRXiD8QlGGHF2HoBq0Be77o8K0
8a/qUcv9O2bm5m9wsvStMs+SnXym0AUkoZxY8+gx4zt7YNwss7TTuEkexEuckBuRFkKUJn7EuyF5
rw3NwwtQridtzsBqgJsWbIOR1GbZRFzJoMBouhd1KSFBf/WpmoWnOoaAcT60/B2zwwyMvPNulnWl
s++R5kadosaruVR5+utpihLfsOw/Olj3rxfUGIxrruMJgnDOvOw1PYTkrXtVnR6BLM2X/y3NSnJS
ZiCC4K7ghHAmFRLrs3tO7wf7Dyb5hvXWdeeuSVKBB3Sl1XTMyPyKd/LRPs9dB6PBTDWb3K0Po+Z4
K28JVU/Om6JG0OdF1BUuO4smmts0uYvdS+rLz+x8OtHql2qB/zofFz4pzQWD31QiKDQnG9odA6qp
S2MOILZ9eG9ATfg4+ZkydAUMjWrGsicQ81XzEXMrZBcapv5F2kbJlVi83dpLw3t4CPKg/BCWGpI1
9s+wihUKo60eaaIO2qX1fB9CFjiJT303vZlxWwyOjBc8N1QYeRREUqyEm5zCMPm1ZIbia4cQiLpA
S+IvcAGPkuP4XlHKHmSSbGMOgVF44efOtIsjvGsWpPln+A7FzOuKvcR3znIkyR2sy1Og7wtD7rDv
b3ViLG1s0vhPTCFqynMABg40s7PZfFoDnFR7Ho+WzTfacvzhSBJF2Ooumv8a/s5v/LfQpRLu0C0v
iflcSpRr+2A9sCZ2gS7xiHEPfAjB9np56BhOd3sG3Wg6skKe/vNH1tkGtqiaR0AmBcRJVPCJmnJ7
l24G3t6NkqbbP9d13F7Wn62aZdOfoW3JF38Wzet51FnRDgciHDzC6R32GDPETF6vwelxipOpHRmj
U22bEhXW3nJPZFc6bCVU//LnP+nULXyOPRMuO55wJzLuTymueMnne0UymfUqQ1R8Cf1eMfpZNbd0
kkuO7ayMBtdni9Fh480R1eLhPMKNqI4XmpORjdC2ikrSmGLzgwJ59p7kLPllsomzNPCFUUe7ysF+
uRkMl6kqg+AK6DGafQZnbkeg/LKS6qBtl9st6HX75sXKjhSXHPS4VV7BaxsEqLCjI4+RS+sv2gFB
DFcXo7dX5Qrju3GsiGDF9jbZEnXggwRlIMQMfxzA14CzPVAN5+ZfqperiXHf+Tt457ugk3Rl2p6T
7/b2UZ52tz0FWNLn9ifXjRjxVLWmchbSaSVWibDfYisJ7+1Xgp7kBJHl9HOxDKt/FeIHWmguALlC
5yo+5p4zsXJWvO05fmMC4oEJmM5LJWMPf7P4+zinSbzCAu1NbH1kcgCBsMHR2Qbn3z4A5nWtHZ42
utcnyhmRy0bprJB3n4Nkx0sBjga9Ou9Qtn1FyfjSZmEAdIph1A+QahfI5EJZdkrAsdH8KwrZMQvc
xcRum7eYeW40AbavB03B2I/qREnuzM2o633Op+cJrtGW3Z2qvqIjIawIzeZqrSiN7x4CUbw5LkCx
KTE84kIjLVxhsuIDBvZ5rdSmm6QM/FKKpjlHkjDzBCQZcnpHe5cD9TDGYHSVfmvcYn8X+/8nHkjM
uKpOch7symK4FXwO/CezbzIIxSy/kJaTHPn+1YWL/cimAW43yNqbZaMNE12BeV0tzCOfvpNLl0sG
RyaITFwHx0TKhz+S+2mdU+jy/xaaAaXJPOFJ1TvzwIX508T6vQk9KkISNW4PLaBZi/0ytAkX726R
olzzRzbMrU4h6baHwBm8Kw1HYznjwYRaykqZQWIqcRXk2k2XiW7lDZs+v68WEVsoIwm6nL3Hpp2F
POQoVjtGq3GwPCQDXvExb3RN950kk7L/uvXNvwpYjcDB7+BIAuDpxsYsXbA1uPj8JXS0xWETU1mX
ZL/7QKJQ9KLGWiMeNlM8nrRP4s5BHmWhzHdhaae2jG/7ZIdbDcTHqZ6ehgVmWJ54jAxGJic3gTJy
evtkyd5WkX6IDmTmw8BeF7h5COv82v6Og6PAsQG52dVHLxY/yQFLKK1rsbQ+Z8wSTmh10mSmYoEA
fx/Y7OSk+zwaKgQUOkFIExriGr2HqqEmYannnU7Pef4A4hIoldryYYa2LQ3V03cF/7JVNQo2cz7J
YP3dEkwQz9SXuT8RfK6eDzFhTRYWDKLp/juYTaObs1r9R/dQV78B/hBa5Mf/MMVfX0md8fxF5I0J
wyvd3ilRgl4vrgKQOM9f9PtrWrhnTDrA9DzuSPvyHSkO1WHj3aWjkMNuUcS0eTNANdnunj/cAz/2
Tgat6bMCCLgl9HZdGr2d7ksX/quvmg2a8RDhMN2il+c48/ZeQN0LKasoBRsSTEjlwTls0MhOHI+8
T3EXvkbux14ZbcdJzoheBTMvGzy71q35/f0tn9p/enmSPjaaz01/D6b5qJUe8AwCYQGyXbUaLb3A
38eSKS/gBFe2TDotxdQH+nmFEL1HUcRgKmzz5+JmVmhTDX6Rk0wJXLDQrxpvI/hjhr1VEXDZ3CKL
I/ejKEmH8tzl9cbb5wFcAvW+o+4DwRwe/xBer3FgU6kr/U/lE8ykvTFMeD88/JfieWgiK9no9d9G
zRs3OU0g8pcHs6c+AyHfWEXs38RFMSzJwA+rW22FkFevbtvNUhYWN6jfHXcBjGMGpVzj6wHBuo9S
2OOS+1gloaN5x5INaN3EmMjuXRSd5bIHQpJePyKo7Rn900+22wOfXNonFRa716/KYoJqAu7lznyp
BiSOM74rT8lozJKtE/0Olp/K7QMSZqOzfodUL8yGhZjc1bf5UavgNZBctN0jg0e7ahZoS1RZWoCZ
vyUI39NmiPkda2ZiEQswv/4TcaTMPEYAdrI6YQZ22gFv048QXHDJuLYxSQn8FFwFpGnnNknt22LB
cyVocRyqgv8gx7YBpyl9ZulnKWtY6aWzUu86VCCTio7RCqqabSbA9DOmdP9UvaPlsCX4ghhxHqRr
KmhfgrwxMUwNLXoHL752ajsHa4P+9Rc14+vxX1PZFEilU5ZuZuW8CyMrknGtAyxti7tG3mWdxyqm
CyrHoF8spWYlVVVdMe/F3Ys49BaxRKeWn0YR/Sh59oo8cgOIRYGxEWhUyAmmGg0OAtf+SsFo8PIz
UedJTcuwQ8fBO0qXNRDWpV8EOB8oT4sGt34rr9d1XLvtHLJUbCovOlR4I70EGUaWi9SE9HZNrBEo
ExPzc/TZevKashTlbfRPCCGfQiZpxA/Rc0FpIs/FT5HU2izhlD8dSqXdGvqPrNazlOJjNX0zvJRl
odqGQI0DmIMehePS7rUUQ/isBCtl+erkc+TK/wlR28+xBPjM/++WaKQcICeWwKnsYns36VsFryeP
367zIhZY+g+3EKfpbCy6ms6ev/QloajBmRgsgAMtrLv0ZedcInwtRHIwjUxbvm/39YrvD2Dq6Jb1
W6KLJoYESm8eMVv6ymZRX04Ry9D+bU99D3nSIuVp0YLPuUQfe+YHCFl56yxfGEUaK32DQa3VplMt
MknEN1hB5vytomCRDeF5Rv+9hpxkntzGSbZoOEclWHiCowV2gxjCdkRjmn67ANj/ijX3zJdNxa0A
lNsTWFRi0/E29SwqWnRzTVdPNdcxHtN0I/qTXjwePJeWy52e8oIEoW9/j5pvwCBNsjkBEQR/OKor
yCjAbjUgcF/69CECOxWelVGMltBtmkuH1e+FxhMJwmTmvKTRll9BDtC+oo6Ua+J8hERAHwwgT+9o
/CEl/ixruUCN3iqiHifvN7rv6dR1O/lQ84s0QbRyW2I4VHFqy1IgSD7Cbf1a3WaWH705yfmp2CQq
wITNgTZKE07AiYAmBoLtfUMUyXzkZ0l/8cu0mKOLrbbzHFvTkk4wDV5StIFLjLvjSHK0JFEexe5d
TnnGWNBLnNLA8s/KaNwbK7VHsc4KfW8ET4bAuoj5dfOuBubgsOc/w2PMpfyAhUD3b79F8SQeuY3X
YzKm+5Us2AhFuZelHRwjZFiQFf49Mo/RCKf2wJqeBVnxU6wwOR3Maudew3X7+9LrYxncXKK4GnCz
zoF+anJPhvLGKdd2wcWJoJmABUv/BtSuziiU3KXhw7pWwfPxbT68UXOCrUMmpz5M/mITk4V1cyDA
9f8oGwAJdbCJYf4tPRwD/PrC8RfeHZGljRXN6F1lwH6DIDIuF+tHORemLoOXhzgfSSEO/ePPsBtS
zs2m2b71PDBv0RkHeAOQ0Pxv+KwU3/6IC79F3zjL9CTOWHcuI1OTQt360tTo+N7TfuXdKBQprRyw
bBK2dDK4+cyn50IAt/PY8RhFo7Irby09qs6arQDCrWVlexNqtEsCjJB0ZokcRoXBwKnpcgciStbF
8ar9vPq4bAIR6o2ZOfjmjRFWhrexfYRXT7pkgmJlUdHM3HqXhLTzcoV9TlaDBblGRstII1+TPueO
OpUj0s3z/rvJrOUi5+65xrtryXGBLiqQb5Oq2hizFdiV12JpcHOCro4RvB9hQpz+jHNaAmN2qIkW
YceS/U5zndjgkSPnuSYWDDWzKgLkHsx2Wu6M3OMd6bd3zpNq9xJmt1EYu8xzeMs88zmMXWrz+7rr
y/iHMBBLlNU7QSIVIR7h9PJ6xyyQG214opdj0S9A4nmZRZsgeqXz+vmc9Hmvwyc/hwq8wxpywN26
hSswP5pWpsAKwMEkTdWrocqf1X6c+mHmpnL+/mFexgm15gLXxfIoCCGjFpfx0SKFIoQkqSTy+CA7
1V8VZIQiQGxvgGfUZ5zE1nczBTbsqJhbFXcIooxuaI+op9W1lbB+TXTbFuzgHqb3T2KL7JF8eH8M
mCvmo0t+LIASChicO/8Qpx7dLIpVLwRB5IkTcNwQp5WsXbTCASrORKbJEhUwG+CZO8wg00jrFJFP
pti7z4Zli1sIQAdFb+DOR3Gf/DTl3GfBOuBc2QXH8U4iqmDQ7/QPoS7VhUC2g8di2wdZvsNb2CJI
uEHC5CRo4o+/iQoPocKLEQ0N3FTeCrDGGame4MCGGFo7rCfSxmE7wm9t/5t/3+z5LGJhVBBZoo9D
V09JKUcNovBU3HgcGod0pRtJgl8d4h3WGDD4CcLzrpWx/r9eyAIklusCeELzTJwXvYopPV/ET9/U
8PSu8mJ2Zq6qQKDaSTcukiwJwJtvs0G5kc5ERjSBETtAEA9iXuUnThcsoVSpZ5xvk/L7nRPNW6tZ
w7bSTnai5mdSBOa/WhVi8Yff5kXqYb5bk9pu4olKojNJR/zpaiwiR0xiyi8ZC9QlWnCP3oNGcQ6h
CM9zum87ArlnSqYWEArPI8wAl7kQ4bFtUc2hooCUnByUueCg52d+hIfPKbV6dqIkIe9DN4mhM2oq
uFREge+HmdOWw1z94r6tZwvab8iPcxAfn2wSficvNz7LuE4z/AVcH4K2pjhr5rpiw84IuMlH7QDY
/reVkcaTYe4G/FX1XYl3OBOWDlJD2n6cXMvdv+b1JewKTgxqVxAPhy0Y6aQVpJZ98YIMCOqGFTUj
Yb83D4QTPfnPZc935jZXykyZ9/VTnQWwIuUdJkik5nJgr4wtfffPke19Apym3o3hGpL2pzvHsdm8
r1nBrx2NSUCvXF4eLPHcJ2dAcJXj7IVQpWeAebOOA2p5nm8/ESbMevNApsYrYmTC9ebnnH8GNncZ
lcEcGSq52tYliPozavbdRt4ZwNcd+4m0FEDK6E2/Iwgzv1eSLmYRo/xrLeq+cJLpOvM76CHq1nuk
O3WI+GANCXy6aePh6rln8BYSRGDyZx1QgzjOQsKM/MeDAsSZEdvACqbzAhrEvLvrGjfyCTw/4jPu
2PT+QfKpSj1bm1KExbOIxkNJMvnnuLxyNWx16bYh2tylU2dpXqK3ShU5tLLhV06wW3Q1LKQGVLhs
HLbtoemf0pKg5SoMFoJ9CdrBMY2sL8y3WOTXW93Yxl4/stoOCaG1U52v5LuRUJzYQBcJwW7NUObC
51k0yaMPJrE6fnBfUysgrrulQd03/gFH9KQWtUPs1WqTnjB9O9/tQf47sSgEsv4l+ckMF4stSAjC
3CxyxmiHGtIV3ehmsFRDHLdT4SKEI8CxsFUn314j4InqUUZ0EuYEl8p8J5PhyqJo+w6sNPLeSiIl
nSOpl7AxIKvN1i95e+mWEVmiOMeEDgONUIdoJW0zAJ58T6noYm5Kpzol5JuEwZw0aleAmawqVi0+
Maeaf06VacpgWsNvQHBDtXr6Szh+BWyjeoUYokg7oHmchWKsWzW2nOz98yEGfIm9IeQbKQTp/5qt
P6PLHpycgFczhEb48o8CUu/HAsol0xSzHrjqpcSfz5knui6xkgvL5n+fiSEEMLa6U1nuxTVXiLwr
/IMUSmVaiXWGTbJC7H+ZGqf6lm52O2uEDLuaZXVbFVg4aG/cQbwKn9RnrDtYwLTpWkz0Wf23yDmS
n6aB7BuL8pFBU9MRp+OkCSeRgt6bj3SL8o15+zJwBs6Y3ngWfAyZghZBXB2OQYCI0dlF7shk3z1k
r6PMjaEhT9i588eGJpfHbYvs70VjjsA7+XuN7/P9KgJF6XMBvF/e+kHKtzcWHYjdLf3epZU2ltj5
gnYxw1PqaRSQol74YzFGVQiz7U+S0bIUL1ZpgAO9nERBlEZAtoK3X5yUk6JCryuhMZ+GYKOJEVr0
Tb3AdVkUQHCchvXYfCUVxKiPyDqQbwzK6Fv+vzDZi54Jm45zASK+PKieYUJkJLn+lryxYb20SNbW
5S/W2dUSRFcAtiCagB23F+g3tNiDOvGASnZ6TpcuiynCNjIKycaLNob/orN6pXQeGqTqEUaPZVHN
oINcl5+OtDG9MADU5WsUHB/p3EYlfA4jJk0ROwi7tD1ahr3/mwxo6JrTt2g6AGEHg+YVWRQq5EDe
lOXwZbnGm5jq/mR9NLF1+lgJule7u4A6raHfNqi9F58SjrXCslRjTQ6d0ITvHpjpvX6J9pwsodj5
scYacla8UlEF6Jt6S5C5shPqywRJE0IIcCL3vxNP+RUyycMSja+oPNewRsrX3K8vlhPOZS9RgRyW
KNWD0DPHjaZfWUcEv9evnf3WJKMbZ3Rt9cRzL4KCt/MahIyn4E/7c97Kj8VKxlSv3ZB9ghWM6B77
KYHtNAsjChKNv8Xv48f0KTfx/7MLGm/rHkNbMa34Po/ZPDSfv46bXKtjJnGIvIOJJjI8gqMXMzS1
LF5yRVpKMJQxOHnK/wawAGPmRh9kaHCp/R8yTH2XI0oKm5ecMMQxRIGCbn7xeCSkHrDT1SsDAbsw
i7/svYy6TKBGjZuovfsN6zRNx/CkPxUQW/04VbohhhSVekoyhlKrChtUGadgKp004HlYMO0XM5rR
5oekXP2sx6l5cCSYKKLa3qH1q8S+FG2U4BmWaMHwWt57/zX4LDZrQ1l6P5cO8eoCVUwC9ll9PpzJ
p+RJ4BMhwjFNpyDsG6XTWkvewLVxdsN8w+O4y/Up/tUhnXfD5m/vFFiqHMBTAiSPnvH2t/M02vC7
q3bjVOgtvTQ7/Bnkv/9GQlVwDtvRa8QxBtAU6c2vKBsxTAifGsoq9iDSb5IuZVCMHnMgRaXcR7WS
NZhFElo9jV48hhnaAPfsmJ9XbtnjCxHZi9Bww3FbPSLGRQqZHjMdaJb/8yc4sqcD6jnO4smP9b2r
HHHACAtUZFwgUPZ1DAVVhKAXP56saBBoggpOvNN7kc74KJeIMul5Y+JAjfjlLAW8Cm1RZUiD7YAS
gVF4mVln2cEbSXyXZXj1VIwYE66NhkwTZR4VL0HANDpbE/jGsqO6EFxXVBMSIaO63j1kslH1E+8Z
zwkL6OHKT+uOVSYm2QpgxvB8+sfNyuTxaRksAyw8qRriOKBM6b/3W2I4efxUiFQ5VTfxv+ZZ/OHA
Xm16w7RG+udpKhQ5lbWoSagldAZE1h3vlhaDShI+0woqJiMs3/0hYBc00CuAnTfB6cGE0UbiqH6L
pVsIbiDaLuVkYkAaZtQ8BRkF2tqUcqXoxkdhAlZc8VB70vySc8ticL1jhQNEtjjE6fbihY5q3fdm
cDppR2soROqEGYZbaenVFH4U1nnGWlF/r+Nc4ofk7l0MGTIX2A4mQX3am7nacJZzCWiuRb0HX46S
P0qDa0LRI+GrrLQu8YvKB3wZ/n2KVQKGqt1BSiEz7INYDLbcrRG4MZ6qwNMpsxrTgtKJ5waZeH7s
Fw9xNcqOoS911crRK6AqZqugDFD6yEtRaKZjTQLPJK0meFCoCXwcx0rP0rNRwkfj0gEnOVVWMRsx
De5l6/CL5gLn2TXgWwWzV5ALjgbUO6TN649kWl11UuzmeksSYg34KRbda7rrgi0hquOUR7mk50dr
1aurMTre3mHfOy+wpI8UDRhFeworQwUilvzVRjxLk6iYUhx4F2NPXinpW1S1VtsUlaEMd09TapvR
icgSx/tWMMFuAjsMC4c0u02OQwlpEyFgKaylkPngDBzuQR+HjSMNbfOUUuEbZeADDT0AqPkqeykw
vSRsIOJA0UxH/2opfx8cxauspVpPWXwqfof4HpzVXDOZ0HjJI3rR88+v2v22tWuXt5I2bS17aV4q
C6loexCsDalqY2sz33F7QS8T1+qaqP4eZYzhcpT/YfiexSDcEcjR6ES68D6Blx9N0b14dFpjYN9O
rhElbHqYMlLxwOrVP2cDTpVNdk82hzn1AD24WAI9PbT7DD+Z1kFmjKAJ7P3zpDcY2Q+Ii/Ob9UVS
gtC9CBnOAGA+pSeGtjXnyyPmqGRmSZ6G0R0aXK3Rtc0kr/AcjgzY1znzHtSZvgYeC7qzhpXOTrr+
c0N98v/bZrfnPKfMtSCwAsiSvJdxTZPAR7J9nK7QXbEsZUHZVmQGE8UVGCCADWJTeZS3LeQ5AC+n
DBBOUqtf6Pbi/aHThGoG42K/ohGj2BuvFGgjoJlokjImYutaXpdWjKIIABJMoe34Lx/b7ELFv0Zy
ROURDDEHt8JsygsYoFbkFhj74CJ5Ck0FO1kgrKtPNYF/yGca0s8y+jluzb3sEgJe05sqvSLfu99B
KljD5x6IYmhuFpzl1yVLtOwymITNnPQWgorHJTVgls7MRhMqtXUJhPiI2i8VhdJS6j10btf6quqa
B0x4P2qBAcadgaYtdw+XZgk7zT3QmsXdP4Oo0we4lNFhNWUi1NSOT9PCk0h88Bd319aX6OmDzybR
zWybgt5USDFGiDTcPEFR6f9OZKyYnov36iO4l6ZbKvJlp/bMvaPBniZuZz69YMIkmq/oThlX1STF
LhXeZk/zRMEzNkDb4cZ4z72Y36JlpOWkrxoZBMhFl7cEa8bUi8FocRW9fqlxRU+ptLeX23VIAHKK
mhVCFX+T/bbpUGhKi5LroiVamSlb6Z4QkCgbVDomlxoZs+XOx6DWr3PSn4mUpTn75CFNZr3bel5P
JjP7/zgpr9FDVbtgH++LZNwBFCy5c/8SRamXbmZb9temB1PB3iE3nt3lBaz2kTyNPZdmjIS0rdZK
UjAKHHeBKhdRfWoufkJc7+iO7v5kj4NTF0vZxswIfVvvQsNZcTkyhzWg2UxoG8duQUSllnvX/uI8
D4vZLlfYtJ6g3pULE7oJ7cgpIe1yQXa5aJR+SPmoXxsRY8RckgQdAdvbV9PTjKjbqgu+yt2bTAgO
FGZ1VbjyZtKMmNMNoiK2ydex2s696SJd8rmkj0Ty+qFb+s4967hLMHBLg+wm23q3edKqKWFiRm2v
LcZtgSaaGR+VcxarDc5CBnqF31zrcv2P37IbvFWgLWxnK0B3/z8xPTSKrKNTEohdj26bFkyoNrvB
ivC2eZoPFdKO+XaM07fgV20dd2M5slr2osg2utRBCEucyLgW4YwMFlED3VHHy7rQC2oHbv3UN7qf
sjC+deUr/BwENUjDg936EPfzZpg4NESaYvae+WFCO1jGLUVvGPz84e7k9xiHDSamEI0GGtbdgtQG
xBTofxshhiAoFtsajVYZcD14/kEVN9X9CxyeMhk74M2ZmFwg4UrhcrAyBqqJ/KmNivteadU3PIOA
C9cXkWkte4HiX9EBUpra77ZfonEBRTXvxDVoPOR50sDznMshEqSzGaed4UNODlEUR4ML682fX2FR
BtHQZAJPDQgINHTJrWZnOSIRxa5I5r7Lm/3KfQemrwvhWxuGD+mbmISm10cFgqwLamcLuZAa+C+s
bLzEiBtQ8AuzqQkryhz6LxE36d0bWD4XI+3eQzenNl5c+16PQlgzwSZZMdov7VXjnp72sUu2YF3U
TzR8Gd3NFvy1BL4QIa3gpaXElULqet5Yx1gRCDFubD/wYz0CPxW1muHmMvGYTE3qx67SpaylTUL5
7b4zh00Lm4k8E8hTJtH6Dwkto84z576eqnn0Q10BKfRdAFgrZpZHiy84a3bJwAMRcZk7NNVqLeZN
mlpsCSMcKzYViCNuYW8Q3lJoBiS5D/+/2EyykVrTfKFWQp2cIq76nP5foMf27HlfWY6a8OisGDzR
mYnpX8KqSR+4bKwHgxkBk6M2zFDVB8tyGHvkPvhuPn4LW++MgAUoL5Il/r5m1DNSBC3Is6whrhbB
L84409pzJxrMwXohyITTvgQ4sqSeja09j8PIOip+L3vV3+TJu9wYu9W550UVZd8KHTcHU5P+u7LS
zf6ON6RV2T820q6m6dSJAGBFTlcVtxoryUZZBQKnw7ayoDOKM5j2VAG+wnFjFoqVQQUYUc9/2Z2p
9b35cDPBeRyYsCDoUZuuzPuh6fmXMprBLkb4dpboYNQl15SQtUBijEAJFqvJmfYsN/wY2auQAPX9
JI+AXy+ehsDqonxOTwqaecLGyZ1a6D3TWHFe7hQExHtmUScad3Q2fVjWvfuSZy4gZXMj84K/eWvU
jMQVHDQukM5uWtZMZiEtt+TN5Nq8YcWM60moOPOhQ8H5Vb76uFjOmPc+W+j1kIe+nevlbqYwYp9c
DyQ/y6M0uGfg0RFzOcXqurNCO7P3vqp52c2Dbkd8znnTTFmvBIYkW8LRL/7bdBG23/q4MC4ubBr8
a6BdqTNUXBruZ4fxBoxLbyB9PtbxqfukinMPOh+SwWHJmOKmAJPzovTVGbK88JWhNE13o7WHSIOY
FTG2U3pqwp1JPMmQigdIoO9HTBuFnx0FQs5MKunegQAXFNv9i0jgZvsfbsC/ChlNaY6ww3EQyHCM
SynobjQXy+KS9zktWdcQRQ7a0qsWzg0zJlBYzkMMLwiAxnVsP719xqkeWkHcvKuwlhEPKdcpIwp4
K4JJ4CnInuLjS/ZNgxKX6Xnmus8mRg80+UAaHVx7DU56TX70XCn994S19eJM8a1/jUX5BcU+Fbpk
rcraSwb6UM85rbP18EsaGEID086jyA7Xye67ITW92C2NAn6EpvILbKsL9l3eLuY7mjqKP2h7GFpY
n+FOZyxSHChI6StcHa8LnY3zAScQZkSV7tw/mjSmfArc3tUt5gCjGv7174Ovii8FUh0QN7+gUelk
40Dxq1fmtapZNwd8RJRJE7+Wa6OWyY4SRvCYRDCrPVDGOa2HoWaAjWcL1MVuj3ZQPr//0C2u4IHt
9kSdiyVZKewWdzE16Op5/Csq+mK/EtYTliZiWNZx6nLkOTaz4kML4Jbdq0eW9w0ddCD/fm/2BZot
kNMhmb2yVKR2CViffzCLY96qlQ8G380X2zTwIYW6V1YE5vwbSZ8VJTEK4LQ+Vt7mO/jUFCeKR/j4
e/22AxwqeYjpm0E2yYuTHKx6ZHPcKl/YAqHplFiy8eqP/cBSWSEjd1os/e0h7vwHHYrGUXFYJNj4
2GodHpSvkP6nUxTjlQxtybilHQJmbo3p+5va6lNdy9hBY+0egHBWeSGQRgGgjNPVADU7sWBpH7DQ
iCYi7mRo8dm4F+Ndj/IoVWobllsov0pMTJLzELg8ydQ5CsB2Di90pcR/W1rhXXRBrSVStxVpzJ8k
910kn6Hzv2/dkljUivUGcVe94kVSNA9aSAjfJlA/cGzSuItn3HN0ib7ZS3HioEOqt+6GyPqYEYqH
2hJ/f5/DzkueHbgqpnqrI+8bBX474DwjmLQXWk4A7FcO42uyykvmSoK2l3vlY8x49QfFqRMeK2tp
Tun0V2vfoebHrGi83ts2VYMn1iu3OjKZSIAP23O2fyA0N9Ia2UG5v3aALcPDgFUBaso0I8wmwumL
xjBDKM+LFqQ8D+TIrXlOmqKjEeYzztFeo/5UpFaA82KKkeazfkpuzJNbS4ZA7QagLB1FRpQ9nNtf
SYV+eUumQckNRXQyRMMJqrQQBzE44jWUzW1XHnYnUrUGyGTJ6f7wpIHsJ+WF6AtRD/kfwP3Zqywm
B3rEqeGYzoeeBL9pJ6pmqz82t1nHI7/9VQcs9u7vWnKyZmJgK6LTL9xIvU16BZnsg+rgcaX9Hs8S
Oedgy6REZS+5vg+yyhMFPf0CVhIwFkq+SRDoYRzBnFOmrwnP9eU2LegZ3if9pQzZWgg+TUTkwsbz
18aBEHx9eK2WqxV/PjVk7DDPQmevrCvJ2LWC5POGSvGHw0AUdeIQW7jpOJlaTSXQxrykxCQq9e12
tPWwtxBgu4DMFowsxAlX5FknuqjkuX/8d/+7Q99U7s5jNrPdwFRzPNGqH7mVuPdVLQ8CeHvl1t1h
ZR9KicUdC4H5h0YzFOFBChJqQ/7XN4rEWnpI4mIqVutZsUzmpDm+fmGZQhPLFGDm648kYYBOvNme
oRH1t9GNmozQvP4L60uaqGs9/kfAOA8TYsbbNwe2nVSjqwZVKAmUSNeEeF+biEiyNXI4ArjSr+K2
HUUIBBDn68r5EvjRIf3OuCzZvECsjxjxH1VDN0i942mBxUYm94KKwg3cg0TkMqWlAl0pwNyq+RkY
hNKcY1v7llYfGP4pVqRzkAk57dUT2CIBRepMphXMIIxgHhlUcYk1sh/rj++RUmCDzle5KQJOWHC/
thPWoPvzBOSd8fzivBSe7IqFZkq+nXHpTEYFrbXbTz6iK77Gk5daZXN3F8xjBWDvJWcLNk9fqySn
jSuxu3twZf5MDFsyy00XC5DvZ28KXKSTtF7M5EzXQSYyNo7vaItn+5W+9Xbm/l6JE76OwGsrWCEF
RFr2ajqaUXmxa4dt0hGlOQ/PfHLmP55CsuU0dkDZCTT0nkJOhEk8j45jerLOCIV4fazoVMVwf5YY
l3B1MSodSDsdj2I/JzYXTbS21pWQTwtIhbxLzKL0xJAi8iz98Hs3IlG96bBcMI6fE0t5ew8t7QlG
Z+k0+/J5CljFgMzww6ASXjsvyubX9MlsozOaip9BBrXfyN1hgH7kVT4hhReBjhX0hnz94CUNOYV1
HT6W5969vBck+3Tb9j1EPQHd/JLNXs9Gdki+lW86YbKKEpEeXRzMD39gg+v545S5eriO4iAR7xOz
nmZsoRLQLX9FN5wix5/p4bhARtaKwxshpJa18Ds/b3oWaRG/oeoGgdH+dZ/9Zpl/VhyUKdmmQpmW
JoS8mkPk8Qly3jq3Yx6sFQf1dz7vowwjEddFYHanrvFTFwrMyhrjyE66Xn4FXwUAA9j4wn3UlzYD
xjljJkLKvbyQb7qFyvbE7pXTxYtMYeVvmqfKZurQX1OM8dJ2EPxu5/JsRGRnLxg3MPTKFYswOCOU
6JHokY7cxfKwTVoH8E+UQ+YuyW1YeE5GMgFw3uWum7F+Mqk0FrOkesGiCR/VfLcYMZghunmX+24S
XoCIQj+lO5dFRp5SdiKvF5Zkdh6/wgwZheCqfwptZSyZyuk8SBaBUHTxGM/HL4ymbyqA4ox1cd18
WKPDtFtLUGmILLNFOudMnmRbF7AN67hVz0/O58N0czqburrMS40PtrihCyM52iZZPdAfUFQ43nGr
MthLx8uKI1Hg1wZTKYDB87PI9gjeeDrcwR3yb6CF6ypYjPaHtbjSE2IztEcYkGrKuggbkgbwFstl
7s+oaYx1UCF7VoL4AicNT7zc2gZLhViQlHYfd/hNwYt7isaPwft9ojd4slxlnoWoPX4uWh5SS959
eh9Q6aYTFT4ePet9dOGzywE1i1fBpqGpIwJvctERG4fjDmfex/1Sbct4WZG5fejjNmAdInNZ41CA
E6HZhpORVC0tUqWTqblrKS4OE8mwTzVK8hSCcU/gFaUjvz2UNfrNLyIjuRP6O8NS3K+8Le0DS4d1
iPssA/XUAGKR9vtz4i3t9DANiqgnON7zBBy6OCZT8VMCmOBQVcE/lBxu/VYGQs9SD51m9GZ+ySa8
p6pkwpDrCz4fRY80sAr90Zo/5JU5OZBX0q02pNVNMpdsieqnBWlW+C5p2uQHkMwLy08K5X0Qp7Jn
bP2NLpw/ImAzwjZy7fslHbgRJMFdq9cI/uAWaobA7MpP4bCU5tX2wDBcMnyJISimsL80OLQU4iSB
+TxeSWu0T/3cHMI8GNBB2AzW0T65SI4FM0NMbkdXxJaHM3gAjkh/CD+uJORYDdLWkMJgWO0k1vJN
QQy8NEV1emYYJXicS75oP/pTaEtB3yD+A4O2nYcfYgAZMVpNfAiRzL4Jys0Xs5Hgr0LajPfgC8Ia
FEuokFiOdiuBdtCPhbgBeDpQFNF0fUzR4aWQYP7exzGfJe2YmMP+SNZiYdxi9GpUmK2ip2Fjw5On
hbFhhKQEbt4kM64+LWPUGtoGyCcCffFjw78v7drVqGkXYWxS3MPl+n76B8gtIhPHQv+gD4n2VsDt
gzj6ylLiTPtjQ4zlc14EfrESJ4ashELBc+IuM1+NtVmCuOvtIERC1yrPfUGuyJ14KC7xToc0QHIq
yr6DwSUrSVvgVrI6aSZll0Lem5R4bBT/uggwAI57u+SvdfQQnIMevuU4xU9hf4xswAAvcoCzkqRi
rFB6Z/fu3N/6oHkFxOEeIT2XGgbvO2X8ZT+WTiOaJLfsA5kgdIlMGbZ0GKdGwxy76chdVNMIQxcz
fCYblMLHYu7xpHmU91DIEcuZ3+BpO3ZzKY9jR+lQicWIiLLUyGw44JaeXPQwRrTY6lEMgHLKh+25
yFmWYmvsht3ONOUts5Inhfq3Feuhepj/q/AhlIGCg/fxg6JjSMAlp1M5IA3jCbrYofZyh3KRzBoc
eRyV9KbesWhhHyyXDwW3XrA2ZaD5Rc5xHmRKLonOIhWEDF986V2GKPUdAsneE5ztAk20s6NmE4wn
6k815Z5hdru9UzmRk88aCl9sGjkQHpgUl6X/26Gp0exJKlW03l2BCk5Vlc1BPzZcSOPQkh1ggE/b
m0uqnmMbVG95Tn8zPVsbpPllABD+jxc9kZmCmjVUZ/jIRDfYNPUQ/mAjcdFPwZaQ9KcOxvCD6QyE
3qEbgwfVCgGxM6ZJsS9ThjVHo6rAl1wk/vDg/478Ze+xRPqrvgrQPayr+AQ8HzktOxHb3uoRdAd6
LbSoyCFolb0JojvfdXTJhG9p0JSFvsqI+eNFNPSkwH3igLuuRMYsa7s2Tg1BSgYzc1+aF+Hdlc8q
/jWl4Ou3eoZq2lETf8JAG/XRuogHm2mSGCE5Dk/X6F2t4QTKuEbfUfYTvoeW5LQolMG8G9t6gm52
Ba9BowDMCWXh3ZtBhsSl/pehBtYAu2kEy3xIDsSKvLhcouIpRkjqPQTQ92+csyjDY6wjWTsYU/00
ylBq42bDINFiyUSHPZQErBWJ2luOUX7EzG4xCWtg3DphsJJaQjuqlgLAvI72TuoufPQICC+0qmhr
788zgKzOG5XYm1JlNrfam+n9VgLHfDG/W53WpYq7p1Vqf34uG+1UwGZogYdXpSKUDdTiVqT31lgC
z26NHuLqACFeL3ZdDeU+3Q/P0FEhi0JO+ovRVV3rSEdI03vWhVAOY0l6i3LCdILMemfQXBRAirb0
7p20YTNP9T8cJ0KGPPQJev9akrPd/nbRooMXuyZGminzuvgv51p11557FYVROkNh6ysYjkrHT00Y
OEFuER/i5QbFF0mFJq1cFf0eXRNnleCnr2rl1UQPx1DlDQP5NLuXKZDNsgRQdr47NL7cs+USbc5Y
/+2OP2ERqYPJSGZp9SH1fz0XSsY9P+QlaCEhR13aEnNN6m+Rvf0tkOi3hbcgOu02/m5yEXhU0/PP
oYrqIxjequ1VJ7O26Ov8x1lCqt9tjs4O2ww6z687jHfNukUJIv5T9nMnE2qzAkMZKEzHgmWqZPIh
mX8I8fAhQEAXg3CylMoK2QAYDqXOGHCr4DiJYrHQnn4bCU1od5Qg864YrO0UhO+sBUwWKm4FSC8x
VlNecEK9Sg3VzgMBWIMQRrOOlbt2YVrk6+Y93q+Vy9CfR0xHaZhVeh1FBjliMr1aAoFh1jtXd8kz
JgK9PnWrhDZOXsHlz4yIx3yqw5y7p/INrwhGD8nZWxKcTVPTaIc4M/Vo2h4/Hl0vOQFNIkA4aZaY
SgP1wkkBMLrUtJrFfYKIjKnr2ZsHSp+0AGW0g8OBIK8NVBZ4uHdVBFWOQ+pljPYbNEUB1C9tlfi7
RsozFgEhXjcVScKhj6MSTlkuKwzOSe+MK4tpFP3zvRpJ0/mE0jwvgcZt1llbBnlrtKVHpc/0Q0FV
vsHu8MyvhX6rfqW1tnBrnZbNWjFyRSCVzU97DEGGq43DCcZZEO2MoAzM7oKvORjsLL7N3T6syAY0
SWjdKBT9jkOfBsmuZViT1ykndyWi/xubeEiDNyYie8aoeBv9oNW6mj6VVbR/dwADsM53AYqGp9qO
nmjCwVy/N7vtu022motQ4YTwanEzrrDI6HKRJDXBl9QvlMVbbmLzrlc+VrTLgNuhLGJx70qASvmh
rPJj+d6Rs08aFuBBA4yqcpTNPgl0RvAnyzwf7+MGnb8J/7E/+bE4gGj/fjOXHl3a+19Fnl/huc6P
B7VcamW3OMfe5WCoEQ8Ht3reYKBsNVAWV42ermLVmou2Pp3Kt9mzxBjrrcLdYpInEtRUIMOzmUBi
PcNwcnqx/eNwRmVTHF5Oe0MQ7EcR+qxvKQRvai8HA3XCCFWa5goCczQQF7bydMbC6somc/IQf8I9
2sNZuGQqRrWj1ltaXJzMUlp9N8R/HhHhRAMcM9zw/6lC9qUcWc9WDnhEHYz1ARDo5e5ik6C7jw/W
aq7BbQQocOgPkVeor+Z2/BwdOLrMeqyrkvV+pcj/4TvfetJ4ohof2aVhL2qflr1BoO/TJ0hs5GYr
sUy62sO/nSUlplUnjLLIkZ+W+gKda+xHUdFjzytVFhJBElwUerB/SRqhyNodhNadJfB46MERGM+Z
uwcFNPLwQKHrxs6X45A4N1jpMAlUYoOrMl9nVLvrYSjPZV29LTbSu4808pxG19B/Ub5XoDtsJ3Du
WRtd8//99+QU/EKUN+xxi0Me/fLLTuV7Mi6n3lClDGlwinxLZqix3CMrx6Oll55YjtWDs3cGg3AN
eKE8AvdHEEwuh9QVBlgNCzR8tsKk3t1HQ+sudSfsj6hdhM10+8GfwuCJbXIk+ujMU8vuDt6oUAdB
usSCHq++OOM+Lp/YP4yw2N9S3C910yJDoU2zxWVOSXFoOzVIQ8w0dw4Fr89Nl4bngCTpzj5lNdG6
yV3iVRpdOPCVXkEypwBLDKuBu+MyIbBReaqzUbattiqYl5u7CeYJ5J+EqDNPlqAjZntQyh6s1MJM
i3sSAgCe7Ood7rUBwkYrEQ0P36Jw7TxpCf30NKh7osZwN/GAoKoNKz+33BUY/odLwr+k6e879JiH
P+wHiVxjRUJNcYRSvPAZU+uvsBSzxaHJVgYKkhPCQM56+SeYYsfVOF/cxhv/WCfZDOtun2L5H0u1
KlkWNrq9Qh6f9HN5JzRgZ/3uhydYfHKtxodlllFOLrQRfKZnR4Wa3dachT+SGJ/lB66Mu27V5Hle
gOQbm0QSP012uTcobk1ejpdczP0hKcOw0kfYpY4WxZW3XjsneP4SNFsE5rAHRDtlehcrP0bRP2z/
p/rBqswfCpCR9u8blkakqg9fcPsIPFs0L2gb3+0gPqFsaba1hjBKPTMRr0eHneDnFTfDoDqwH+m3
+quo9ajMnRfDyVlf0t2rsY8IoSkYfTPzNqgX9xU1+O5OEj4EUxLgbgBD+pGJhOYQ6lSSqVGnz7ze
siWDE3+6766upyODJI4W1AZsEppkT9FQMiqn3OfvVBNM9f5077Fs8oadVB5RbR4KcsUK4xFuHNZA
p7bRtORQF1O+CcxCIts0ACi04+eLeLS8SldOMkxghz/ozHYH6LcGHyGicEzYxK3ynSF1u+15hcnn
NOBxRd2aieGUOPFY/wql0iiG+l1gxXb3A26sajr3n31Ms+hNPJm2Rv0zUFJ9v5tasvTcjTV4Gi6w
QRAQICgLwmZsCGouF7WX40k4GSI7D62jXmeZCaMpdNt7kjd9cVV/NexteYiRGmwsdmHwjkZVdG+o
N7uOPVNNqYsumHh5JCFrTDMIw+tiRbXWZ7LOVlFcGxzoM+dZreyF4QUYIDhlyOWyY8uxp5yJO58W
JX0CL/9Efimav8hQNhfgSFihtO1wy74tZHkkF/vTJU+LJ2opo3IHOA+8+2jRBTTDQ0y9Caz/4ZAJ
IDcEic8hIaBx3MTbEa9WORNj3UUl19ZWrQrNC5G6V7OKeoaGb6bzW3/v+hsyjv4X2EemO3w9Yy98
O8L4X/gVVPfGoYat6sedRYUMseXgTPnAa2RAmLesI2mi6YDL0wR/WZOC0Ss8tcNBhw17BYxtiXwJ
Dhm4KtWJ4UVBBxywVCosUHwjkvAtHM/6xflT6bSwmlhzj7TkM/LF/du2bl0XS8x/fuEjTz7dAlsI
0ePl/2vcnyqkniOKxNAKstwnv/ParCxp1jUTnHB08Nd5LDCnSxKM8ZdIx6DpUPmmaLh86Dt+Xm76
1IMeEEC22OJZ9EvB+7Gbu+WeNpdQaO9epzGZxP3E2+no+FSBoudDve+RKYVN5t40mNnlgVDDcyjH
inAUmD7u0rYKsqCfW9GXONe3gG7+Z6owX/eekwMWZC73m3ek/Jv7gpt9u8zhK7jaclSk+6tDkDXP
xUHET22rBv4fEFIW484JXBPDim+X+688AWKJD4zkJUYc6B7HbGh3qpQfqlVDEN78Dolba31PkrR2
QZFVWD8ePx6YQisJAKzcvM6fVKiOBaZEfPzmWt6qvubA2p90Zs5qcEJmninZTvoshjI6jwM5GK77
JxD8pJXSdehHIraxbqNd3yhMdTNUHApmqviVw9cTSsKEEtJEwR2V7dZ/e6rDbrRu3JVFGQQePIQa
0iM2+kudZCOYj/PR3vECIVUhnHIf502eeWPhS+TG/Dbe1BLCLfKwHejdFvnuJdRG67joc9WKAIL8
DOnKg6V2oV/Fscu1G7/IFfMHkceHbncEYhqQ9GJOn9Qgy5WNHbbCyfMFlRoExGzAoB2Lx22PYB4e
uUnIyuEmmGHhGmmFl9X5mNMeZgldfGQ3MBybl31Wl7OJbeiva3qKC/IN8FdhCVQS6arhKBM/olkx
ZTL4oGThuvd0Lbls9BQd+7yzwp6gWwcXc8gEgrErtJP1JAcc5mT6oBwbcS4l5TY0U7X3Oj/+Ii2E
ivDsv6/EveaRAsTDbU2KiN6d23ungt5BUEGzNyKE+PJyiq5iFnSr8D4f8R94tJT/QVzeVkv052LZ
0Reggx/qf6RkyeJMrIc2VB/gPhfqQaF99z2Pe8aOclXinq3JoDvsCBf//yJ32QmlZeaHCAvBECxu
qk/XIHeexoEn5CIYc/3G5EuL0xriMshwU4mbLHg+5urjKcJCXEV0wcfFbge1L1Og0JPgTGGMaXk8
o/Kte5G/fiX5fl5iu3U+WCmJUKAON19MKnGMQFaLOajG+rlwXqVUX3QiHJa2GBH868iD1NkOquTb
UPkQ8eCe11f8a88Ns7lpjLEdD37eY2UinYV1UDeoYMtd2YD8fIybjSIoXl8BFnHTTXLRm5AuXikT
Y7BwLHmssFC6AubK5SuI6dY4jWgnQaeDDqQ3aeUgeepbXSgZkZcibVzqhXHjevhgeLBMLlKPpx0P
fkr9rE8SVVuVAugLEheMDyfBdp2l/9acZ8QeI5RCsYU1LjCsTqYCRSHBSh1Wd2sJPpuWZlHUNQ/3
HQFGK04FAv+yttQFCj9HOACrYj4dwuN7XttIIAdTmvsp+OeaCaDsDfy3GEIr547HaaqgUNafmZlc
/qbvi/wHHVBZ6J0U/OLs2YcI8GkTKS3/LFC83mWWaU+FNyoFiZstdZcxgOXtErmh4t99I8t87um9
i+p5QqzGBEyoY18isIjYvvhAtSEqZi9YqfH3XnF6pY0h8H4sDv4wMq/Pp0NymSR4k1B1v72caM0f
WZg99Ri8RB6vgk9jFJ8UWx6DL+pj98SeRgbC42jKhpsttqbyXXVgPzoRL9GNn0B88sYRI+c+H6eB
h3L4apKyX4X3AGxS0UlNGfgRKJ/0Jgx5fwOuu/Ix8afO0Hwrc2DzgPx0AlTG+R8cwQtlOyKd4kXm
Ai7qjZoVMJHVTK5+Wa6P28ADLjfO2pgBix75E2tAjqATpYvPVz1wh0fAFZgRHaYzMYRYyq8C0o7k
5McgdmCqrHUq2ICMcFyPD8MgUGfVkATRaFqgcREib4Fg3qnaqx+gzj3V9QcJK6xtxX3dtyg3MAjN
K1ZgWV7oRRMN3IprTBY6eT2WDhIr8Ajd3HeqynE0zP3WXOdXfG8+P/kpelScRq8lbha6OO/s8fry
+3jzq9IKtbTirDJi6SJK27SarFRJS93lIVvZ4qosQPL/lozpiHw9b4mAoa1oWsed/2lU6w2gaYb/
BO5p3RxNCxoti8uvBTS3lm9/q/bcn9sz5FDYSgMpYri121dh71F+GxceFSuWQD63QIqCbcp6GsAh
+jIYW4iJ8VTv3Xuvv1LNjwObGTblKU1t7efaXEr4Ja6rEUWpO5cJVrpaAJ6OunazjVTANbWMwFM3
WDpKotil0pX1yX5rejnyWDvjpWJz5qmD+c/JP/IcCr7xbFO/o3tlEutX3gI3iI0FGpRP7L91FwOf
lKQ2s8L05ylbF4B6LN5UlA4Rey4wHzyJdz3lYSgJZwL9dYOvTze6Ae/zfOlj5MLWaeg89cU0q6Rv
WEXg/Ai5NqrYOTkZWuNV21+nhNtI7pT86QYl0Z954jrfGBDXIH7v2pkvkKzbgFpOLXTVjKlsGq36
8IkJvpGgMsa17LsKR6b8zqGUhY70b/wZxnzjEngl+aXuqZZUjneorUpnfNm5MMETpgIQklADDmDX
TLnv4sB+ytvNeVIlsgRH6n7o/Q9UBk80JB4TwrScalkBNnd6ezeWg+XBVZQQ1Sj9dicH0G/jI4kV
mTrpUmbczleoyy8Q6fLCP7d4y/M3m1w0pe7NAV6YxUNiHwJMTQULjsOF/i+Hjs2cLVPYKCoovPH1
m2yt96cnhr7LCrgfni2cpGGbJGJdKizZL2JVZMjwWSfxWJlysWKbFlyP+x9A3jX6ijZv2UW1UFdo
n8F0LUwC07aVxsplcFQ15eAhdE17pFATuMfUCJ3SHnaqiK9THBgfxadNWTP0aC7zSXNywvZofROC
CNvD0C/uTPPPDKdttVrqQpHp4spNKl0k6Kn8nSmSjAypgvB1KwPyOpdILgVEDXXRPRwhE3Aqx5Yq
+al5tgro7jPsMRkGu3JY5ULKq2B5c9Bo6eldrdkBRL0CmxJpIzEh7P4pRPu6VavSGgUN+TS020KP
yGXbnZZyrRcgGXjZQtBkT16Fy6ZKgElxRIBXly4dgZPbCTHrDMKiwX0twJUWUjmIl2Z1QI6ayAeX
FHUvvz+xt8ugjdhatF8NR2ZYZaGCRgT7lfZ7zO/TPJVoJiOHXt/cPHzoojRMX2IvdhgY/o4XZzYe
7dmW7RqdYUhdPdZ9m+GLQVh+fNjoEVYeqpR13c/UBPc92NGA4RfWQadI2CcxvE1TrWSUEWghCO6t
KDoPstyfQcOdq2SysikDt4TVj1LeFwbDLtfezsPY7CzHMBFQ8J1Fa2xhqX9yiCm8jd/HGHKLfvDP
LNU7V78oLjNYwgHxQLRN82bqOgfaiHNB2Krg6NURLy+GWw0t4qHsenWI8+8nrrwGnEvOPsXSyeQE
D7ViU9RWauGYPwZidc1EAiBazomGkNNny4YVio1h2Zwt8kamqoZIxvpI1FGBJmWpErHIoK4NpVcR
7k0mMZK9d7iClXFu4G5/kOfsxdWgXhpavRd61PoTS+PnX0RC28F72TRlCG3zUxooL2oOozxDPy2j
YTEv3Kc3VOrmGZAlFpecsxqwuyAzBFjj76YsHnokueRWPUlp4HT/5D3nCcvS+7r7dJxODNMQ2xe7
o9xESSXDVS5ifLOZoVXMroiVUyLTB4wCYaRv3LmAb7kJk2Zr4RlFWkjr4WjEmMFsOP6tU9737wc1
vpH1yjQPDRy6zcG0IZsIk6z2KgQorPR7U0SlkKk7drtOpyRQjC+6b22eLY6dRlJQq1YYHVb4ir6V
qk54ZlIVCT+bOobPnjEpYlTWaZirvxbbkvHM/lXg/P/z+z4jIaoC2p3aHANY5e7dDajNl3wrMnxf
Ge2WMDyoDLMgJWm6GJeAsEM42bPk+Et6nkYomvU9gefQFJ+a3UyF/8VBXp1gXGqFbH4TFhbuPBRq
bsly4eoE1ZB2WkruUbXD00tur8xzcQgkGQ6/M/PsrzE1ZsuWpGzPKNryPxgbSf0zXAWnhB5lJ1fl
vQCgfGoLB9dyaHJqpU9nb2s/ctywb8gL+5KTBf6QOoQhc4zp0eiHp2zGhbEAvImaMKtga5K0kmnd
BoL7PFryXAfpyI3gzKrtB+S3udybepcBEU9TVZZKc3D3ceMUDnHb6fEHsk5pS0hNvffMEdBu8qvx
baPdgAImyVX91LyyjDk/E6wKxyGtD/HqhyBM6PQZCoDR05H0oD8YknqdpZEUIBWqDlIJB/w8TVBZ
8PmFShzTpAlU/5s6UyF8hIaqXuV9ovTi3yHeKV2X9ao24VJyS+0OMKcW5Y2ySfRQgrwgW49mGgz7
i9gdWlgeN2B0rqLHwSKui0QCJAKZUpMYeKXWgIz+UawxojfQ1maOXse7dUXF/0D9zE7uBps6EtVb
qSseoD2QGoCwzZn+kxdeB1w6E90mY7uIcEJlWn4J73M8iS44UpTOQgNEs7jTtLAUaSJOowCr1i2s
U6B0EpY+6JdC7CABVHTp/voKklc3nYGeeUiGM2exvF03rjZSBghkLE7dN1HULD/s7OTiXk54XWvF
Y/ct3dFL8SIR8U+awo9Chnf53OuY2oHhrgd9AXPiwm4Uq7qcaYlDgQ6hTiuLq0BR4ovONXWjyEvI
+HcifHcXbLdfJuTZ9zWN0uYDHYPnDLO19D0lqlcucWew9/sWldBz2yv/r/Vs+Xqax7bZpM/Fn4hB
pwgg02e71GqipItLP56fYYQpvPIhdn8Tm5nnpk+OJcmeBoEvscTTCRsS3AXIA9KqYhljchyhb7Pj
YW9A4xlzPTqgCelxDmkpv1vyj2S8GJ34b2HWVSmzqmLrIuBsDbRVfHHIZPFr+pGFiujdc/4h9IZX
C7vPkhBcpjE+aKH5sK93+LxeIwm5PwfW5GcMZe/BDjYKAeUvGTesl8+tckeBjVgoxJ7yQM/I8iFR
8pDl2pqSw9C4IevZVYxBlwqjkSrUvl0HgZ+Wxyfdu3eyz7TPSSBWO2tyqnR/vEmMdljrWXeH2qDD
ZIgz0c6xsmf8tKAd+Z3wDeJqpQV2ZSJyMwqcwaW7GUkx+5O4hzbQ5P67GHpL8yYgvwbu9Fsu8YgI
C7G8k6CjoYDjmEgxIydWislre2JgOtSWMvSQOffop+arvV2WKN/yV5i2SbHWGTS9lUaNl6HEvJ4W
Y1vRN3gsnrdGIexVJj7cEP62D+5jGQytlqCrD0tKDEgJ//HKAANVP9CAT5Wv2pVlDLeTW94b4OxE
gPvxZ3bBGFZ9FuYxqfdZPVakPgcmxTCamc9rv7A/N3xuNGmFQss6g/wd7XeetmSeHtm0A2VOhm2Y
HNXRkt4yhNfSG805EeLelW4jC1Fj3imHqlIxM/Uoun1MI0nYqA/vL6FIY31PwHS/vOEw1r7mAT4z
mGwOKY899ND8opH0Bzl0UkKvDpS40da8BjcXoAu4m/iI8lP0LQkJPtBhtpHKeFoV0sdh4bhewuRn
UkZuAIxdAPOgjzzygQzUAgo46PXLQXSyMAdlsgNdatJhIuF1O3kncZ8EDtt+rjLK3i5SfcTIbShe
+SqSbReNm2vqL9ocTKw/VLlREdPR3HuEd8NvuT4WQYEivvrgEL5CXuyzDJSt1UoEC6y3NBy2T5Y2
/xle8fk/83pjztULfe9B0bxiPawuOolapVyPVz3kJE65M4DayTlgKqHQFR0lcymOYJ9xsAGu5IdR
CAFMbjAX9pbS5IS+TMLXsyYNxW6gdE9LLJW2CdY0yng6+wr2iYg+HnyKSU2SRVcncd9+obToWkTL
FsFh3FgcTfUSN461+bDEt59zb+bRM2hcaHQt8IpWgcj/u9G6XawrKQyOQU5F738cx2zMZZVQu4Ro
eoVesOdB9cbw1WjgYXP6BdgEFLwOv/Io0PxY+UuTEYZHlIJFvPP8GFJq0obYzqtnsxN2++XgDCmi
FAxr0CvgcI3+4zodZ4rAeTJNJWuEXHbN6ELHdJdxaI2Y9O4jWvobJ/DJcr7l3UKOLLE+vgStXf3k
NUeLd64VkYZhVhCPFdZTMetVrl5u71lo1JBGUqe+tigQrBbHyWSaup9lLw+yrTPiHxoYcP4OzXx5
Yszrdi40XRDulKzocSvFqqdkx1CPOashR5YQZ5bVszEiC5oryg7nMVbskRwo51VHzkWV4GzXxjsD
64aPoNI67/H877K44vQnD4KVo4rz2tqM5h3G5D+KqwpMOj4jF2k8fzP1gNFIuVVEvQB+jL/oT8Bt
6kdiMMt/ltcUG+frpsMhjQfhRFsR92sufOPYewr/F4kB0wMf759TcWChZUeMA5suQSrPGVVInF2N
BOQUAJhmmReCLjnbHvzBLw8VrY671QL5p/ToJi0R4WwgvuL8j7ukeXy7KXjiZNfd3yBTIq8ZdDu8
9vZOlFZf46G2l69ANEf+DhS2YUg8KLVuV0eNVF5vPxgg4caeJ4jwvZg8qff+6DNzlc11+rAv+o/c
L5LwpVTOjFsQbb/p3RfQH0IiMefsHikeS5gA9gZ6ok8rU3Cgf4HvGltJkV8Y2Nvq9vDNMxg3B/0v
GXKGvgsZfRu4kyiH5hb7TrfDGaiF8/TjGkS7cFjuAuZg4n3e4z7UrO+MxTeiy/LxJVhSo3NFTV3n
FKhZ34bCf7OQFip8k10hk7viae1WGPtAxqQknUIR21NINpdmJLhQYBhLEW/7YZSn9FBnD/lqu2zA
eus+CRqSzUkarX5UybOJTvHohJIGM32vUKOOpwbllmiO8vSY5XdTUcqw0vxKFv602FaELxl9OON4
KXom/Dx6UTUC/5ZviaOupTxFDwy5rGkRpWf5phz9+cjBTp67WE7F77pzdrbawZuE0OrBQW9tfG+4
WvEcsCWtc7do1YYTUPalWu2xvZK9tAtimt+bXeVYfgajiRqIw/gUsPbhPOI+ZcbrOkessacFH++l
sF63auxfSwGuV/NJYiAI540hm//04cAJEoeccjcLBo257DZ8SfZL/bpnpSdmX6C4DOpa+Tsqw+rz
M1XX5W+w4Ok1xH4JeRzhvclvU+LfPm/uYBmezg9gmb4hzljXil6QMCl7XWupUJlB3rMQzB7tFt20
DTuzn3yetAS9mdjdO9cv7wkRKiEXRhmsoCTixSQWm0ylvRyPc2H50qFLS3F5m+DCZw2oWc89B/my
TLIxSRNCZwrbVIsY4B43ZZCuekvc1hcBXKrO+e1+aUuO6mw9SN3HS9UfVcuFVj7Zvcm0jWd9ABWP
/RyhpBeuTTjxH9OvG8q7xOuOubuh4DVwjDaV04qP3H5ZgnOi4+ZyiJOKekS2ouqt5kcylYvPo4eN
p5DAtzhu92I40r9leKXchd1xHQ21r2/3ZK1K477wr2Go4qAZl1AxRYqzyOCH1NQzSbhCmr7la5TC
IM60Xfny1+IDlEYQLQnCDoHgcqXk/EnWSeToNx0xam8iwRexR/HeeCJqoJR0hA7nZ9amupG6vbP4
vdTmNBlto4U1oiwHOIZqWX+bYFH6G0Bou0G6TdSq/kB7k10n89E3cpF66W42ZN/O8KHqMefAakqa
N8YoyEQxZxFq4G7mvHyAGqDaBJDQ2G4qUxFjEdT1spLLbEFUPa60K13jo/+Lbt07ZfWT3/w6WWQe
jOHAXg4Vommp7zqeEUxJqbdQe0MB+FjFkc+aZcKxQiQsoiZa0MQqMUVdPkngA+vLXpdmztd3qs5n
OZz4GgbVqcTRHPuRhKm6xFSOOdWV5lEH67VWZtHkFMcHHzyTcxmpuP4Ch7lsORRegCI5zsT/C21R
NzeYchSwdEQeJrDPuzHX36VPoEW3eyWRmNkVmAu0Yrz8JdKihx+kmnhMmy2AFXb43Ymi3UxcWJyG
sWBHhqiXxADBIPLgwDuzYhgTxLFVelnoDg8mmnQV7/ImgmwEhcov2hSE20kZZzT31BzPQuzuvra+
oroAx36ivmHW5lRetYy5wfIWQhKuhHPpONUnNUGxnnE1bqrzq6Eh4Ol2CTHTlUu6JQAH10o2rBW5
+Ze35dq8SObPX1k9hVEMw+9qax03A4So6k/fSbzsU1tmwSxl753JffbMPKORh4j4pPDXwlFJAyQ+
/EnL3H/uNJYqE3aQWPBcMhtVD6RT34bRh0Xb/rkDMUxJTGve6wvuAKJ8llVfEuJXplDYEpDezJYj
vDajv0o1kPBigqvYEpuNB8IKiGi0ITq02c6HgSEusCqaIP1dJJkEeW+1QlYGEdIfBO37QUKU0ofn
shjbJmMBfqNs2cGU0qyCQFETdJmv8gyeNHo6dH1u+7UdN9lJHNRPVB15UA24t39ZJIZNGTc1qTxq
vwF/GFzS1d4SJwf6zDizH0jlMKxwIM5F54YIUp6mzNzzY8beMv5xiQyjPtKhEQEgaAvrsn3LPHTP
MKvHsvqKpyAzumDfSpvCuJDrVhQljxGl8ZVjou3pzQxHMuLcxt+EWC1ChUA/EMF3GNPNmMQ1QaiE
s9nLJdqZptYxyY5OrLwq6Qjfw8JWIAAyzOBxXVQPxplrTJnQiW2yUSapMDGdNV6iCURDgb5LpLL5
VB4j43FWVfdHAk2XO1n4tvOA3F/REPi0JhfvbhaCeBlfSH9YyrAV9iVv8C0OP58FlZB5ub1onUfh
KWJj3KZXsQuZcLBFdRhDpPY+tsFnO7Qp3yclprC9Y2zUbs4VWtntXDA2nRowZAuO8pZieM1aYEwZ
nTOUA0eRnw5tNCRGnDdbdGb+esP9TACTNpa4+vrdRG4KWt6C52EJ6VKSB0XBJYDdHfqkRpnITLat
FgthdYc17/00jzEsCqQ032/TTtJ0qBLiOoX3l7MNN2Q8+/Aw5zf7L3TgIngJba8RIeLZ9bMjE17q
RlR5n+UDoW1fqJiVp9o+jHUn1Ngt4te/NxyKWfgv2YOPdWMN3Knl94kde+ZiZWDZ8zvSm/Mup0SZ
7HKu+9oAkKCGP4P4rfMZML9QEJqKsRrUwLZdPll8ElbzwiffeXT70brhTrfHiJBtQxx4VOZ4oG28
1WeXuSs6Yu/GpJZWT7NJpevPnfVFhDKy9fl0LIb1MxHa5Eiz8Pubjlis29MP5+NYKGlcCNzjO4Na
iLM5je2ab+WtC/vEED1oInz2XINOWkQ/rYP8RR/q8s89nQXGSoloRXNODIqAeLNXGjXdIxMSiDAj
uOf2khrc5rMQmZ8XpqfNch8kTTcsnOLC6Bapj5AKapfOMh92+OB3zZVIzKMfJgCNB9xUgBUyPShf
nJ7uhHq8a4tMPxmaYpIvDyyfuxBcS67MypM+pfKEsPK/h49mwvAJ8RAPm9YaFkoFAKtOdJYRBERP
BYJHQgJ6seF2zVJXhhyKZxqhJjYtVqZRVwJ9ykFwHhTExspQXxT2LNgWapOWcj+0cOClpUlS6+r7
qqLPd0ucltzDADOFf15AAS7XnWR2CUm0mSo2gEqvbDintSf/aIxqA2sXB6ZrNoRdy+uEHoZXHhKz
79fenPcZrHTbL72jmOEPtM2mzsaOQ8Tq10pbwXEfoK4q2Xm16l2McorRRsTBYXiM8CkczZl5rFu6
oGJS17B5RGzDaLgTmTTTHB8v7CBvB71Uumt6eO7z07v+nCHI2DTSQABk0MNQ4mr2nTOM7At+TZNl
uSddh/LYwTCjhy/QzUU8CXwHeoIJt12ksCbE7jZlL3IS7c/Jg6cPtK+MUajcBJXc3JWMJj2HVanS
P0OSjGXdif1fwqyBVt95Ta9wlQObtI0XzNZT84ZbnhDWiB8WxA2oAgPZFyv4RTi23lsivcVzi70Z
G8u0g11fyvskEsiKubgnkK6RoXQRCDa4x1KMmWp0kGzJS068SGfdDdlBEayeGNLA/Q9C8m6EbgvU
00782Mi8pDJVNuOQHXV2h9ab7kGLkcsHkXzZcsXrm79gYJRdjQiqQZmuHI863hzJFf9dH4dmqsgZ
z02zQSTwW4ZgDKn55kYWwcgXF2dpmrToUOEQ52OqM3116z210HburDjFQpQg4Qhj9LahwouXJBfh
cIVN+k9HYkutlWNLkcLK+lAExB3jXKkmi1KKBx5EMU2V95l6PKWvWIcH59xl6Vv+HW+ZqzoB0NjC
K/QPEFcsMoZb8OQAi3hYjXfSNhOt7yqx7K3igMwwDbH2pSxxjH3pyjeJdiaWikdWx3si4pLUURTF
13VmKIC4kv1JzkqDdycIO9HAK18EOfLdd0zxdMgLrGKj7Np5CfyLLtTobKHBu2igK2iSWW73iisX
pId9geM2IPLCd2/Pu6hUDiAzjAbiWrxHO6jrycpxtrMnQcXo0k+ZvCMQUT3OaUUozWZ0H26f0YZk
80YjOg5yeBymplw+15O4tkYQFDYt9sGgVhO+Qlz/br/5/vONau+8DK+U0Q2paBj5z6lKF2Z6esVK
g2Q1BwANyZuocO1WpEFwM5q1yG3EbZgW58NA7T4EdxEleYtUkFiCxMkICO/5diDaw2Ks/7QitOe2
dLy9xdmcOX+4cLhhzWn5vqGsmsMxCjW9HSoQweKEJkXf9AVSxuV8SB+IyuN26adOT+lI20MGg1sN
AE13gx4NaFTRERpnb56roqHNGfyT2bBoNt0k+2YVNcdOek8TfIZWum2YODPaoUolFWLxmjg1Lntg
yBlr3YC67IqyrMKFXmN0eRYl2tJ8FP7HmI4LOl9eyk+IzbrlkxJimQIzbXPD4WyW0xtV6dO29TnV
AzY+PCCrlBDLYr2zLKmtLiOf9Zq1A5VJ2s7JZi4skq7aNv2sxByKKlaXMKbpxjlDopPvBjQ4Ipdx
9rjTgltNo2n6WmVeMMb/+i6XESlScA0ch9vwH/sQsBLWcqhMbXoMHt6ojnqQoiGIvEe8zmjd1x6/
d2Wofk0IZqc4hhmCKcHkwYLK/Eu17yCD5rgcLoLgcsLwLtmE0p/h0Kj3sFPl71gnLoayZQtxYnCn
THMYoRQ1xWoffEEw44nhpHHuHopyT6nlQiOCXbzyNXUIBuesKumbccEtWcWKTp8F3RbUwgjgJ55G
Gwghi32MJabSHqaUbky+kHOZFtNlyTHFVQMagJsTyLMb9j54M+F5y16/2FEbol2VcndBlBhSUYP4
qr7CGRBhBUTC6lu5uZa2iIeAy9a7aDIuBqIDuyVpKwEv/UiwsZKrZsVQJ7rvz6Yi/qDWYPSVMnJD
I/jpXuEMbkKyKh/QqxA1UycObnk87aVHrOMYuYP+Mr3Rs0btkWPyCUyHd4zOQpbbP3MztntXTQRN
K4+BsIRyinooXCU/72cNSX0IXIHmYupAgLtkxFn0Gw9WH69AVFnNLz+j4WgiiNEORyYGQt4adPd3
HhVqc+JE7R6ZAmLy4bB3eucyA3ZatLIciJ2J0UBbiCYBu9GNglnhtC8edpEdJYygvHirnw+pEQ6K
YRMtDKkth9F0a1oLhXfv2ySOUS6HqhDy1Rj7V9gNrcqbrKWJ0IKotJPzCES7gErzPDW6mcQ8b4OD
Fc3Rd+kXJHlKvWMysShtU/QB4ic4c3t0Otmc7ba9750/mjjFdGriG0fcAa8OlH8GBSA/FUA2ZY4r
Iw4K+jBkHIBx5kx3yyBpLgOL5TuzigqFXygbpb/T1keyqtCdJDoBfQz0cy+BBVdhHrUH4AdGB+Xr
R/6/slq21gj91WzPfcRv0c/N8WgoVmBXI2IojhNfO+92M+i3aHdxh04U/Z0+9L2M5DJSPsd8v2pi
8seByt+WJM4Hmwc6jGAFvZitmlB7YY9S1A13j3COVwMO0llNZIk7sNhnvOlruG5fikawgJmW0CxO
JaJs7LxtQUEkoDixYfGROhw2X2UsX9dgRxJxVTqRDnGUAO00aJibBXtbpltCMI3b9xRBMnjTiSD/
NOA/wTQadPKxe2qEAhO/XGttiMIrLjtihZkvpyJzUVwcFHeGS1+r35EcK2JA5VzjAeanEb9ldje8
sXmoJf+gxPI3XZOH6o/KCnNVWWjh69D5O0HBM6mDCPOvmfz8XnkVDalNGPyguFewyZD8znermn0Q
FUt75pVXn52OcQVDCGGdmq/Uxr+zAJ+UECcCLWlffD8kZfP8/02+s6aCyovGuC2J2VIrjN8tResR
+kx0i7EasurGxkdMRWiWwAHIoYqUP9HhdUDNPnVt9bUhq2HJl0DffRXWDfI6oB6OuvTa+6lWfyIN
hrKtVTyIB4Fc2DcAjKuEeEf2Ig/vpIodvwRp23T8Ffq/Cl7y/Oo7cYMEerirtFs/VgWttfmvUH0y
l6DUTzzsKfQ3EljIe5I5BDA+dElyqeKNKpqvxOnqawmVZrBXYYqjrdk1goFO9GA2iZQi6RBk/d6j
eGqQgCgbEWyqZbtpUJ2CdjeZLbzVz+FqnckeaOM6AMPbVdA3k3AGmht80Ez8rZTgz6w3XcmxuyHN
y+zNE/6Fp2WDexxeGpUK9FcKYlYQhOTR3isKfg0Lddy20oGK6hqZY81aSamovbmE0NbbUKWbTJvr
ePiYXUBahxp1xAVXZ0aZsdKwHMqSR6+bR9M+0DsedGISYS/6oY8xu6rtfe8bYt7C7AVIvPvWc4CX
jYYx5nqiy9f0gkPIdVVH0+TETUXd23AJkG4u+BFI0AdxKYE1iZnZuD2mcOW/YTlsondhtKWqHlHz
uQO7swNedj0lr19N68eEazhrBn7tNjBvPAo8F6rdS3Ui+86KlG2+fV030EZJ0SiBmfKGB/GCNRdt
eLCeW800+5J+b1P4LkahUJQlubRuvvlEVDkG302DKF3ZCja2rJdp9NM2YEiekfmn7gxh9m0eEkuF
IrxfONHGj5npgf4AcJC3KF+B7Eo1sgAoJlXA9ALjIgTakmdFrIpdOJ3notvmxJ4QVAiA1qo74pWB
DrWNIlhRe4kImM6r93F9jsKtKyjC2Bkys7vWNWDyTgsJvrPoq48s+bExOQ1tYi3crJyMXC7C55yz
u/iEcyw/V0CoIl6OJuQW/8QKDa1f4dG0Zco/gUA3UFfljD55zh+g6TWkXnMfo6P4nCac16ztlRfB
Bsrbn0rEb/2npjk5Ik7ni3lTjMH/5oUM7Rx6xmzb57is8tNgRUC8o3CSsBve5Ms+HUOF8PyfWeBU
13gNw3HL5cJkTNVfjp2E3EaBxWgHxgCOflOOobaCwMJYJx62yu1TT4+8W10avusqCl+TvFCWCEfX
+ABbT2uPRC1QmwiPmYRBl1LApYajgUQmCJwieNXp3JwrCS1jnf/Dfr8beuM7DineW69ORDVQuyMd
/OoA35RMul8C43wuIEE3csuY1KC7VWWwFzGpt1ER0RTYXEh7M7ygioAd7m0blOEaAy+NgV5gN6eB
LPZ3t7KRWJ4KlAvmREsna8VKPG2TGVxP7i9UI2pJtENk8xuFlFPEzyMFrQUItlcr4M8J3rjP7PM9
iznL6ghwFQQmCdERQC8/DciHBPATX4GJwuASYBlT37c/qQwHGujGrwwyPqayViTVeQiJNj/1kK8x
y329W9d8vASw3codxxJdjaiYx4eRmAeYwip16NpJ0Aly3EPFmxbs5HoaFt9PAG9aPf/PEZCPFJWO
H+xhn/eqafmInOnQ2GaH/gSf1Xl1e7TCYOYUZa+zPdWve5w8XG9bq/o6PjPGOxgL0K3osWbRQ2XH
/Nq2g9YVML2d7A4boa5LdHUIuLbsXDbqoWhCiEOSMZAVhrtp0pm4SNEVXuM0Y2b+ozG/hWDxG9k6
f/bVGyE2PPNfAWtPK7yRNSF0nVvwAbp7VKBxxXgX0Ty69uQuzMftJpbEoIBOPt2iJnIJi2GpA56g
hHIda4nNg32v/iBxek9tXcqShM23vnLrcRZAufnR/FgOEg7zy8jD224dSA6HaGD1lpPjYGMcA7EF
AXvfHEYn3DaYXMplGv5l9sFq2GOIJ2OjqezdJP367KULGYRHKR1336j0JM7lshHw9HL/IYpFB9GW
iJVskKUDj/c9/8fslczFi8kK9d4aFfSGDXFPiU33+ay7UlXvF3X5TZUr4o4tVTa0BhWLihzioadI
hvvsdizgqUgQF07Ug73hC1rWyS5YecC5l7MMEAn2a+Ow2gN+vJ0viO5o3HmaZ9+1AjoOFo9ecO5X
lfgR7dgm39AsqmH3QXaXajeEWcbzxFOpSeKWcu6SQwD28OH1HXw0Rm9xSA1zquOsp3g4tpaMzJB/
XcH67sxNP9KQmXq9D1MOuRCNeIPPda09Ge4YZ+Hf1uX9ljf4iCakRaUGiI49y4Hmw1R+FNREEUYl
j4gm7+zQTqbXcdGhDF6osF/E+XEBzRB776wWfzdV819F2nM34OA6tOvesfSJ4lfnsIl4mue2bj0S
hDSKtvIcPYikvnX9OCkGUdN74v7EwJdME3++GRi+0YnX8BU785Tk2X6SnhM+9CQ3thFs/L/QhVna
Nt//Dqdmq02pQM716JSDWfPHTdgrEh3mulGU55O5zUTqWLmgGqTkJUv89PD28J7aLsQle7lJ9Nif
PnJ2tWyw9/h3k4SbB7n/7Nq8o/6IXaDNqCHrdOjTSeugZwYph0N5n+xpsA1cjlnthmx9R4C7q1Sd
fLJttHfvUik112/s+v/r7Zq0kHcvUUVjUlR1xruPg/jNG9xNEAOzKzCZkjL0Vq4lw4kKMjK0ZPR1
981cAsvYAaNVEX2dowKEnifjoT4t3yHcschcrr5Pi+MGiRACI/Jhh17irW7cCYWTNu8uSqZrMmM2
lDSgs2eKPZ98HwCOhk/FmmYXcv12rmn2Ra1QTLiANCemOSMyO6TUYBCgxmi4qGBN26ULA9/LIWwk
B4zCUcllMVEWRWR7M9qHwxB8DUxZ4B7ksf2xI3vxz0VdbjCPiXVs7367ZjS5/GDu0zBNmdfNYLoF
EEQlhkZnAui7wVfEP9vZ92deARa0mvhIWAglP47/RcPzgbM3bAzrLusBcH/JylngKATjUKm8zk+u
r36KUfN/Or4m034Kq37A8wM1XGIjwZ7vJf6xOLJ3h1ohRLS64bJveL74qg2+ozOIibnhLgv6Rnjb
jeeF51NTANOzaaoHb0ELxWfadODM1yxyFpz3OZicATXrhPzemQdfygVhK096oiO90ntyMt5loswF
G/Fd1vUWRLLdZ+qwRuMzM9H5PZ5DgGbV9yVp2jm5I1lT3z/OQWgOGmPKyMS4MMi4PQPq3fe7DMS5
hZCaxU9nrt0ND7kovvbEduERP+kLea+lTRXDXXcBtfZq9YsOMAjMpOhx4jr2rVZoucI+/2ZTxvB4
kjAvJayDXVl6gyIV1klInlTsObG+N/U6Gs85fwNMNUrU1ijUEbE5V5a23VKCyGfluzmtGz+6gNpj
BGbujerqDT255FsqXQBHSLZtyc9k88vUTC8TfWmOngp2PZpUSbjExlpELkBVnPq3h7+F+t0Q3EOg
WB+LFQdjO1SzeFgZeZij3TUaM3Mf7DgEISrpxhnKLYO+oUWHiDmI2/BMJXOZDs+0avXGkel4FEyf
Sk2Z2RtRAGOTZL0RDLnSMCIsnxVNVQW6pHEMgMvoSnisF6ENEsvzxUdsHfXipg5vIv62mY7qYk5F
vy4ZF56vTMqi25Bbgw0qPjbSYYN0FYpa7kxPf0G/k89SqsuL63+HKLrSt7wBSisNV5Glaw++RSSF
/gGbWnPI1kFJN2GfMCswV8iBHfr8kniQQfdfl4BwOdnXCT11AtA6MNmBvirjsr1sgfB0NCWBnaE6
IsbmX1sTO7P9XzihMZA7e6Fz6Z2GIzarARIUWHJaEfrPuI+PWKRWQkRGxXnFt8tr46PM+OEkotsk
ccAYuuqRLCzac8iH5Xf/A1oyX/02jGiFEg4s2N/5/elYkpnHEMsfhkaMPf0IhkNJ3izN2POEFuNw
5BiebWa53qxGqJV+EUKdSEJC1J8aW8qfIbOr0tPCSRyuTHl1RFJ4Laax5yK68Njl1sXPuuCJJv54
h2Qmd0+EBDn410T8tDKX9oGYbQdCyBlSlR8YN61NOYKsMZqecLY61h7DnLHMR0XI088f34oDbJRN
WVTfTaCYcAOVSGIJlhiVqUCKfFjc1aQMlDYhkNCYDTNvnmqd5B7bdYHVmZsS946+gQuF3t1X9wXR
Uyk9jUShUmoeypQtuO+yNhXGYi+rZZF4DuU0nF92APSRvuk5HN1dwUPmgwEiEb4GR3ANGBDkaJ7/
1piSYt7RCBghARtKum/OhzaEYEfFnRQjPOzSOmGXIL/ob7AJSBJe5g9V8VhVmPNXy9VdLskrdtzU
0Rgeytf7mvyDxbjEx+yBjH0bwGz3ymlGABB3c1/2SlZAJ/a315fA8NR71dzGSbxBhgJ9ixcuNKH+
FKWDPBgiH3Obr0GRTaXDFesV6Y0z+91rsSXtv+Tb7Lf5H165muk0a8MGFdBv64F3LBa+H7oHFg/6
xdvpz9umUVXKsn/TIK3a0EubMhKSF7b4m+SqywPmNjNzSQK4FflWfTRVxkuQasnj8ckTZ1J7hAz+
aMEyUYq6Tczgqr71377EN0njP3J9zYGRkt7kDa1iCQ009A4WPKDxtwN5wcAdJuZHiRum9NqDyAKd
v25pboJdAZeEA7F9bsv7/EHR0mTERG9E2iup03nx37M9J6aV124JOj2lpdinVVUwjeTdOKiXNGI/
ezFio6W2VaQGrdKWBO6itdQK1LJjrVo9G12xlQ271mdSk+zGPmbs/lAypz4+TnJ9NzL+PNMVlixy
rYkRsc9fUqZjfQLQmdH4o1l080pdwf15/s1wy+H79b2Lsx8ViUJF9DimXF+2a8jDZQ/7fyEsi/jl
PwU670EZs2hhU9hC+XNh5qBFO/mPDfjaVP3xqNTQEbvGMBQQbMc5EXmTo6saF9cnC4Q4PT8y+P+u
prlHQpM1PKUSjI6Enn5LQmMQga1NLR8c1A7ZZd50Dht0vOhWn5cHi3nRK5Tkv2UTQTMuIklfU2oz
vWxs2MzV1mmyR60BH+xkajFgCfbO6m1Xa4r+6t4KNkgBK6blZk6eumUERmvqkDV2HBbvARR5WzfH
V/8xnGgV7hqZa8qJvkZwzud4PPFlu6XcsZWoZ/fN/3ERX4Yn1p/dbT88NiuHkd/4Pu8joF87/wmT
o4cFhS6zPTHlBkrITCs6B1wo4T++8uaookKDPeJb+wj1gqxAS+uTlDzS6VjXa5Fu7oHJNDOPXq0p
Y7CJdsV37qYRSTjUH5QMJWJZ0Z9AAaRdImsAngaHj0IJFYv8E2Ibc6i5ImvmWXK2Ga/WiPX+xSnc
/JbXioZD8pYkmuNTmRZFEFzO+ExL7KsDE9oILwiVKj1vlc6RkefbqNGFHuo4rdMWO6RNnzgcCO11
qQY0T6FZI1aEv4r/p+18VFKkEaaX7OgXpgRJHo6cTEav/YaKVMVK7uTLozACJPeMlI4dTeXAeSzJ
HeV+x/PRRNvOyvmJa9F+tgfow3UhDpj7pBST8AWkOKVSJT3qPixquMjANhC/vnrjnX2rTre8PwA9
rIXmEnc2X/Xfcz4JmREOSTns1vy9CVbCZMujdxHo4/hoonpSoJUreOAo0DK4PAPuH4AS+uaoO36k
hr1zipCgpOOYNRCeR+MjiCVR/bdeqMgRqXKy4VCEvK3JSi0QduN7ZHe8gzukye7RuXCORrTXb0aA
Wu1z4SfgNs09SUjZE1Sb1k/V/mTwe7IKgM0lPxMdH28HDVzDDD9Dw5CRzQSSoTysryMBekCKUgd2
AYXVR2sAJjw3bj/cLVtSzeldQPfIYF1GdhZwmAd0ONesmG96OG7oQ0ugHF9JNk704iahChyAVal/
KKXivic0wrzBThOcabFG7EG8gTkgnlKRMBH8r+e8wzcTpg9y4OxI/cw2uyjX4Cw6DSB0vOpE7U84
TZWX/n70mNrgrEziS70/sJNEhLmEATRdL0TrgWaohj+st7GhOJEuwtjEsWwAartolQIJ2lav1eRR
mmcu7CV578gwiRmXoVxlJr1ph6BI7+Nw7Pcf2PdxuhtdlJb7mIr0lnRqnuCAe8pOrJUv+YylMFPI
RhakNTAgKuLX2bvBSJLzY4Pr6t1gkG+XsqdT22URKiZ4nczppgFouAomqrPDKHXqJHbI9XsNdGkO
DN/QyMytpuu8HZKnYZe8kH4y+yeVFFsNnssoijGZVYUm2SJce17b6WZtal8USWUhR8G7PDY/a19m
FV4o+5fWe5avv2AP8Q58aCktkqx5VkMOv7/BatsdRwN85xZKO0cfHHNjBtsFhYvqopNxV/ITCTYi
QrEFHEkhNk0+zJviWaK6AnmdHktn/nYjEL64X2aLogeIW4fe9hOd4c0Tce6xZpVM4dVxwcEP+Qll
42vspF497n6EN3RuWXiOUFd1qWYpR90qmr75pLwlgsPNLAKbNtY+nJAAb5eJxVyJGWUxFGZBvM4N
by3qB7vNWLORmnKXv77ZZdJiRCER2X6YBCCBTBrrgEg1UBI3XiQlI17EneV4jOsg7ue9j0+cXN85
FBBvcwaCQD3e7jWugWauoSK98gmJX/tOsHquuCPEt2/qhRGLXZK7HKA+YxdMlL+YubW4pkQI5wr/
JbMALw5dgwE7MDzxcb8TSHAwNmYXh/y64wqfhB+xsP7+p2szGgX3OeZQC1bNwxafqYQ7ZzwaLoiP
DpRACQwyRkcYBvvPJ9WzBM6ebKtGAr4UPh+D/UPok5ycj9XkwDjrVIOBsAI5lQuERXpHQcX5tzPi
QLW3c4ZBPtpmKT26OwWd6hbIYNUvL8LvFNVlSYzqcNg5x7mkbXn8ZvgTi1LXPjpicdlbkFo4/muk
Bujwck8YZ7CIo9s8fmp1FxpH4ejD8AstN1fqFStU7PsAGXXNGtyajpeT9dV8hpvBxiGVZN/Ody1w
7AYfcL+1AXUINPO95E1bAg4XOO0CvhBkj019Z/8T/xDmUhETneL8faIWnWr8y6HL24+vWllvdzJn
eE3yfLs15oPDH0nL9j+2lcIYvfGT116aZu1Tmo1ia3VDHfcjllfZeDFZ2cnGzO2EYvFM65l6RReU
s4LcRJHf4sclqqkh/tmbpNy9EPTTRZcMDbfphI0cZ2ZOG9uJ/TOXCQ4uECfVzvJBrqv6kIIjQrYW
+4uT/f1YxFUtVjl3rBUXlT/s/TXXA+1kMiuzPelmkk2fBFqQzy1c+ruhuXZS1VoQsYtNyBDm6+v4
DIMdP1mgbUgnIeKgAwfNlE34XeBu3ASXt663IFmjJVht/bo1EmOherIImR9oAYRN2BXvVBK8rNZP
ltUDE+zMXIOfiCZnUEWIzlOy4RTFed6t2Zmi+CxeeCp7tdUHslh7/oZl19nVPHeRHIHr0iOXAZFd
thb/28/VlF8p67hDPfV4/RB7UXV4pMce01TuKAyBs+2iWIBPUIbH/gtA7RbkJcLN4fDra/PfSz8y
PLPw/pJb6bfL2SuyA1f+Byx9v3bty8f8OjvlC+yhNTbyKdAG5frK/txzCnWK686xyeBL2ciofXJU
vdgpuLegCeAFMMJIRwRAO9CzhnDd7BDdavSus3Av4kVrwKIPJDavy3BcNDz1qjGR1rBd0LDcG2ga
6xou2FyW2qSmIS01eaBA6FPNbj3PYMHv5bJO3qZ7FN+aaWoYR5pq0Qxdde6feU9hT2hxuIvpg5E/
Rsiy2GACM+FHrshbsoNjxcstQzJjymbFZi5fQUMaCIKC/PLcArAFVyT+ssQS/eMAlLSKZJr2vckw
ATmon7SK1Pmd/h1UZTUHKKNttPjl15Of6nlqjU3Y57NqSvIWmSo2FU0pSyTAWByDSHhHKFVHAPyD
+PvbBs0/JzF7reP9m7z++wWY4QtkX7VCPxQZ+otutX+gCunDMe53bQFTfty1UOCRxPMPpEuucaWe
ogp/V52RgJoF67erNstixQHPNX1bFYMzZ3IzXHT2nr85GB/6G/SVujqu7AsmiUiUFbRkhJRNynYh
LCbTgCnCnsTuG4WotrTPRxXsNJliHhr2hHrZcg+b20gzTzDCpPXkqvCftw8vHQeXWZKVyOlc9eZM
UC8cd3kOJyqAfTPIb5EG2INKw/E6KC0L2dXDFoz9APscvPNPOck/p3Y8xYDHz1jpd/t7hJDr4vGg
C5SE9TQNzh4tNQsq7OqEgioTfrSSWBEYRNN+2wL5oo54vXqNNg+qZe7uKbROFZBK59Irtn4TaahS
Mm9fq45DgDU+ZlPhyD3idoxlUXWjdzHS9ovfyuwdCNiiYCO5ie31Km7fVV3JEjuPukTpYcFkm/WF
iMd/Vhdj2Unxyx7w9B0nfnzDo+LBQ3s+qZUtKVwZK+4XvRGUDJiOY0JoXETesgRAvpHcyYs+qPff
ao7URT+sQK8ixzVSHTDjsO4Yw6/UVXv8gepQSg0clx+/W7NFQbjePM5sM1IjJUziGS2fTnXZAxZC
wfVxo9ADWJ/hooTSzDSWPN4V048g4D81Iyvv8eg26t8XrMVKjrPw0yApc2wda1h0S0p4HGHY+6aG
Eyz/mT2mFrnj8HsDd0FIe50g4nXPPEZra7iS1XoEJos0WFBPvG+kqFAxTeSzLah3ff2pL/w7PtOP
rXzDB+pRK70VO7ukFSxa0YLUh668YLWtjFYP2gAqGeE78vK5+Sec27ol/c4Nx4GsDj0XHU0SSQLF
4oSzPbeS4KKlbr716TQpvzpUWFVa6UKloB1kDKfFAjeH0eimq3iakRbBNYOcr3Oz86L7KqYuKqLB
bQxvYCi+uZbCcL8a3HK3rjPH4GPscHkrYhc58sAydOp3SEadegg1y2nHr88jftSolaEAvDI7d6sk
2soODZposHSexV8viJsIZYYwLr/AIXLivvPya9SlSe6SDdAA/5DPLIHNABYGPFAgEj1W9tWRnE/b
geP23Yl/MIzTRY54XewM94Ilw0U9joHSOIUY0H9QSGVslJ8UbbKy9D+RRor7+qP6Re97b1vbHItO
NDGKRlX1Op35Hz8nQ2UjJgRNUGXMZG+Np1zJBuLrjlCUU/ckc2UCju9S/VuiP1uAcxib2YzwqX5H
qi9cUl37wpvd/ZnlfXJi3MvIKlRH/ju0hqE0Vr8kF4PUHQDU+ekHeziZbSrhqSEM7YfNMdNL/+sy
+6mvN1MUjNeSbJcYAyhmmBV8dMbO8jVMnlohMM6D+Xr6Js17IanxbgIokAc3cQHVZR022bkWMk1K
/dbzDeaYYRC6rL0fhsarkpRRtTPOxaFDupipGQ7xoTrdH9AGtxoFZTWMW8oJ3GdCVyML/uU6h1CW
g+yUdI2FHbCaxbxalQMg0yNOD1GkOUQREDGY9QY4AaSTPdbIdEKkiQFtB8b5NOc1eYzcSBa0ddfj
R3kYPLCqqQ+g9dcLoNhiADZS0vQCjrnS6YKPHoWk3tSYYxppoV1dQg2AcWbRI50SUyrYCyatbSTi
NPEdgZGYJ4AbNvKWxwOP4u8YGhDhwivZJsdnF+PhaSyWKbzUpgdB8uoGfIuNrvtSgqvmub+Lld5P
bYM74cL5C1+eU1owcVIuksrMno08LEQERT8dVoFKurj1/qg8a3aIVfx10489spPjPh+7/VI54yRn
3EAo29B+b/uw46v8LLqiTlePcGgi6V9NNFLSyp2+2u6NmROmorP2Y4tA6cejyNyArfhYTIjeY1GU
r9Ep2dyp0p1ZZGojZSS1r5EmrQuXasNmAm1urqftkBfZYK6oqDMVkolDUXNDxaSjTP5fFADxPPos
Mo3KxP386rpLeOs9WJ7hsKFLxFJdGqTwWQ06y2iPA/89jCvnXVC9ZLbPLFxpG8bKkddIRa4Hyqsi
QFQi2LOmYXa3iVKpYnsOM9zXQaKqKzSGoDpk1v3CWiagO9xjzpy+5OYLuAbzztVEC2BEcHZjJpPN
tRXxreF/gBYo3aB0+H6q7wR/8vabiqGyFC1dKTybAFDka4XtV50nRtKBpAMgVnXkwwxTE/GwTego
Xj9qzG3qDw3yA0W7VZWRJm/n7em3LGA+T3bzruVjqDxdSupvT35qZD+OydxlT4+1O10T5Dwi5m3G
c7euk88gmJNbYM+aV69rYtk8hA4HoLKotRtrQaqJsJIwhKnPCs3986Cs82SfViUme8MKzud2QP3P
WEsNGkCf0Tl2hYgqvy3rDL2+XE93ulgF4DbhNXyCwZu25WDmJ9uhFm3tZ0a9bu1xcQjTrhqX/djb
0VUH8rVCQvI7nHMdq+v3BhZeuNOkSJQs9V4QKbFOL6pWe49uRew38pzoGBwst7cDnnjxYT/oZw4r
Utxjgp7e72KhKvHhlccQ6278wXYAcbAn8SA1xAC0AePITzkpd3tjKCXZbujuoHvso9QoW+POysR2
20KK//fFZZ9CNxzHCMs37ZhEpQyAnghgua/9Utf8drAWB+FJM8E5BGJKWMRoTSpSd66nzRLmLpiV
fD5y707ZMcr7p79rNetPnRpaSjh47Im4ZXGEw8iry5RQZqra3ugYOqRTthTkFRDRwRS2fDNvi00U
vk65YUFJ62LjqIvvH/BKr/fCrleh0EI/bEFjQ11SabLj3G1BYzQ/VuAXquCq311NzJOJe4n5NWpe
ZnHa+vFmwFfQih86OpK2vJV0haFtWMbc57iYHtMZHyj9jwJY8u9O2RNqD/hJJuuOfx9uiJ6GjXWm
lq2dMZHQrBLbGOEYGnKDKrcf7V5/F2ayreyjDhwqES1Okh9X2uvAIU3azLSfqV4dJy7PSPD+l+xR
qW/kzQQDVCdCZQM+DgEYuC1KrkezPqTaXv4yROLP3p2p9lIiAFO4jR3my2rp52DOIZWd5mkhsLVa
ml6TRyt6xZdOpsTeCgn8ONzXABcsNQQASRAvfvCaZ1Bt+nBcU7k1u/qUbkd9J2908BBl67fCRNpv
EeI86bYVdyA2q1Ez+Tb448U7/gcQQ7SSqZa/BJD3Jn+CyZq1FrutrIpNw7sNKK7KKF9jqC3zp6RA
jMnS68e9P2/EYq34E6wrNJrhsaK1Tc3PRbYR1z77SMHX1ADgfOuquNAptWYW6zBVfGWJ8Yx+9lzs
DwEsAtEKIHWF/TXNjm3EpAhiU4q3XNJ9uFNpSzGM+fo80vf1+YKXh/F1pUar07sEdK6dFfHZnIwp
owZXnWX9LGynsOXZlJh8/77XvSGbdfT7uFH9lVIShCEA/o76bwgLJkrUNz6QexVcC9953gQjlpiK
4A2EGpNWXo7iX9Oaby3xgSe12UZTf97M7252/HmawHBAZHpB30ECcQQtc13RAkc98DFMiN0nqBsc
9hV2MU1fVx7/VIRP2SEnQxnSucQ2odaDjjwD2WDepVYqTCn41VpZ5RfpYgpKMDOM9/fEApMWL7O1
ipCTkIo8YziaOhanuhGrLVzWi319o8HLZbVc25/nrqjZ2m7gChLQk2x7nXgE0O1ZqVx6iX9lz5U8
dc4yvYAmjbAk9aSyIC6iD6+4sFUJZSrDdFsU/z3ta/LG1GqhGmHtSam28cQnOuhHTlgEl0f9ly0P
0+lEwAzOhg8/GHreLvXaSZbwCUAK7P5utmerwR6vBJvBP6hGUAKwE3W+R4YMS/ngOB25+b9dRFp9
YvXLkbvodBPoqOhXbNp8k3aqIfsWzV1vpR873P2GU7Op6pUq45sBkHwpXUQu3jCm56luhGVmk6D5
r+2H3bs/QlBoyKMXOyZhYuauttpxdpwn4NcnuFC29FqQ+q8Nlz0xG0uQdtyQioS47rt4ImHuL41V
O2SLidqh+dMdY8SMyuFCCNH7JANE/SIsMbMlDcUEqxrOBfH/kkOto5mkKBQb0l3ONdEErYmnGQDK
cnV7Br8WdDTTCcYpWBJz4pF5+vJuJCzLrR+d4Y0g0JZeNE7kNR1CConwkpc01YWt/v5KB25h70tI
mPVEnilEuUeI2l8rHUPOMha5FS41CC64dfUgfj8aPOeEjQYwvaR+dozHF33K+/CWDdyYlJcMJHzU
8hWHCbA0b1Vz9H8pQhBjowRdb6oT1cazgXy1ab4ERv3+0tXCa5nrraNL6wJRBtHt5ROScksEONuU
gcOEykv4U0WdMmO7mqKPtbFpYqQiWKvZOYmSflyTskgJK6uSWBYGb2awo8RZ6Bija4Ui/dIzUgNL
miE33fFZHgUoC5wo6pWWAgpW/+U4SDhfIHM+IwYLMwD9zKLMJVRiDRYsLhWXIomSDoOX1ckytkgA
hkDDNqvoNDG/uPkCHVwYtMBacZPsGof9lDp0NMfFRG4THaHElEtTfr9zBTZZ+DzGLH7dMcuF+hhh
9ypJc5Nt6fzRjvvQsPQerUlOK8odHLwb8aaRzf3trSqibGevxPBH+MeYJqI9THqoMnirsWwL5gtl
LPwmPfG41uVOBCVdzi7dGV+C4S/tTr6mPOyQ3Vix539hB6byJsqpoF4rA+7yQU8w9V2fBX7+AjjJ
Fve05zu5eZ/TdaOi3z4NUIn1s+x58rgnS8D3IxwgPZf56pVcu5RFV7VjmvhMZ1hT7v+b+chG+Zi5
uInwA44w7cjsJfcHYwRrSOB3ptx7pnxqprcLybh1Q9cybwt7dsA5VbfTSNO0yg2ehhEz4GdYnZA+
nSh/aGRtxl8hJ0lLKja3zweJnHJWoFunGMGtQERd5u8GFa1PYb7KP3iBjsu8eCulQG9vUfB2OnIW
VBJFXQZF8ZSbjjhmFZhKbfrR1b43NXsx++Ij9Bzk0OJsIN6GeN9bLAtVcJzRhfIqH/BtomuN6SCT
AcotPCIlDB2dQew6as/p00UIP6LFosnZWMNvd6GtFtRb6KYNnS03xMg/ksTn9gFdlCtkOrqhCVdL
sf/3FK0Vu6dim6YBzNtRit4yxXyexj0LRHKuVy30QdTL5/WZ89mzSWENro9UjIFvkJiM47Kxx4yv
KUYh2fDd4LP2M1jqadbm2/rnPRpkx2+ZX+AQ8iYyck739vda0Mb+3J1D6PytKChbbaskZjTMahl/
96MfhOB0IHSfBwPZY4w5KhZu1p4NMorgE043scKFGx6QU3tpQtfY4VvgvOhN4qsjD/64FGWBPUE4
AzzGYmpY8vZCyCLUO4gZwCrJomPxniDKVIEabNhWtQA/qd1VPGdWXDgQzpffq8ZT/5mnqRI6RYYx
OuIuXp860cDZ0SncXX1XOYxqzJzbc4Pv0Pz3+rMTeyHjvLHKwYLod1mM2ndRvMuo8/tymcGAipn5
H0M9CdkFbgNwpbmdmTKU8wRf6kX6KEIPLEh3pJDfFIRreRFZ3vaFG9w6ABzrlSydDxN43tjxEDnW
CeNtQGRIcLBKNJjp8ZFMRbDCbHe0cC0Fxgp1iXq9feHo01AkwnevHWUxAJvWtlcLTAlhQQ5uQpPU
GEnOR7XP3564nOniMor/EIy3wT0/xlsobGJh63B6wJffkcB0MIrOHRiIE3fAMfgnTIh7bbBTA4pt
QWgov0TqWn/xNGY1qYZGwXSESi29Faxl3dABlUnDggPpFjYhRRuELSwmyP2KLwpIBp3CS6UGjd/k
aWZOqlydahsbLEcJd5k3D2vywOPQNKj2M+x6it2oJDqMzmP0JhionlGRP08YX2qPy6+KGajxAlJq
NpsNUM6ktwRmYZUvOBY7G6bKw61aLqlaTQ0hdpDpp+8JpDh+y55gi9Czf4mQ/w6kyvdyIXY/3c9y
ghlWkLOUzlj8sRBtIyP+WouZnQs5+xnBgTIBl4Bm9OShAvJOvsElkJ/lBc1vb81kn1QPwO1x0uB9
lUk1tAsT47eI6mZKi+RE/uE3dehM0dD0jmSuOL3p5rnUKg1IsDUNCHewPFUo7dbpjDoR4l14trLR
4uIUHdNuvvyXnAd3Goy0MiXiz6nzgdVB/M9pqI6GzpN57u3WZu2r8OAr1qoq3dmmrDRj0/+Yb3hA
Xn1BDhmTbiJBrTApBOWa/A5OkHUK8qJIO1Z0EHdv5ArnlLUGwhJjx8/1S6qZLGUgDgrTVJx1/J13
xMlAV5atIHG+6yzp2H6pJ4ztvrP/opR0RSyl/6AtFslsqroiPvSq1mr2MD44z1MV9YfGWx9jTR2k
mguIeffAV1lb0ilERRVZvhVFiRKktN6pq71SoDD04Ob34NPXwrqmp1sfFKZNwDkReI1C7+RxNJae
O4xW00pM88DQGn1j8fhCP4nnI69sgEfoLdiX/LcMyyj5BnWuZX5+aZmzz/J9vNq55JhPGzOhCcxl
zYxqypmRZEIMnLOoPuOrXKRoi3jhsXB08JqEMuW2qCSTVdk9n9HuxTsJw4qbYNq5O80WfevFQTtZ
BfqtiElXUaGhgvGB3o8jg830DgkasALFlx1AbufteNMVxwfSsQAWs9Q++r4Kwcoi42lY8gOY8ABW
pmznNtFm2R/yh5mlqwOGrM7Dekhz5IEHM0/Q7JXCm+3hwFZmhbphoQM+WudjiI9xY9UGa/gwryjf
SDBCjqbHOIPkE5jcBjurpd7wsRzdRTocSO4A7D9ZFTK5HMM6bcv7C5C6MYf78vQ5L7hxZnJMcK9t
LrFNWnSAg/V/oG0HlCYEBH6gxQTOOPfV/HkvUbm2BIn4ZTC4ETpNaMYzr8Jm7/C04ZnPjMAy+jje
+HQPzy6JMIwD4A+970pdWVsedBus8W4o3F+C5W7q4c80SWyDqMop5IK/FDEKObssyR5YSIpFfPSM
FF7ep7iBPqwk2tRKC2g3ecrbgW114Lqe4zwCADOscSOf6UKLAwTc+jRYY0FUBRegTYQGzxyQJvHQ
wy4b356tWN3OB2PTsgWjPpB7gOiLvfQLhKnsaIiDfqz44JgOTc1wPb+o5NS2NLaZf/BAMqxZvakl
2SOui0mTyd88eKM66ngMSRKu8aCx+WHnVbdTvmESUXIiyx7ZEqIWvQdPWiXevqxf5Mz/scA5m8VB
95jK2PNn75gg3I6YsBSoAzvaqofZBxmn6GHx3gX3nPiJ+U2XmPGa6Tq1DgHSjtP5MA4NDnQJGHaK
02JkMhlivxg6BpKjPWOiCNM1bhBvTrllvlQwjtMGZ7JNT1cCSL0R2xmQpK1m9cFXupdDi9EQ3MKx
A1JI2MGxJbdSaVVZUq2dW0qf3xI6ftmhootx2exMQyQnXUzci1n3ourNwig8PRNrh181G1QAfxV3
gTlw+CQpo2RWTZDcGPmkee5E2G6I4Uujzorp6A4ViBVXDzyzXBRKvJFDn/HOk+Gl+21D4CsIY+so
UjUdKGzBPt2WSOg2CdhW+wbqvD7cw+gct/iUSKe0Cg//mYmdZ1VysMiCcfw/3V1we4+RsAW0Ttz1
1wJRY0ppkJu1fkGS6PY8UdJ8BItYHSKMu/vEeZ2QW3vsqLZThahk0GobHeAODLxOo82DaOhIBgbG
mXip4r6sUHX923D6Jc9fNg7zkIxGeQQbo88x/0ydRv8k0WQzkN+gST7UxCHB3ekgCV8TOAeQfaSf
ePYZgxx/UvEYQ37CM+zsHKWw9alGDUJQ8co1hNGJTW/XBuzmZW2gQ28HceqNKe9yOZVJoZOU7RDS
FaOupSrm8HVsae4wLFY9IFxklllPop7KnaSF55K/wC8ggxF1MzRl1Sd6auYJCY+hWDLX+xEe9E34
W+v58UMeHuuxY7ohfUWtphQDZqxbCyo4xDaYfGldS/OJp45wnkhW2qRPHCcvy/L9z4KPXXKt7QRj
TdI3loZO9c9v/v2B/ewBLhgeFR56CWJ8zUQpb7ASdGsogE/2/rLCQ9WPg/laj5hrgrqt28JpUx6/
cKt6Mj63EeyzCtsIahMzBTx5pLv5GT4pQtobzW7uDjq0GEwGBDFgUTKRpVEBr7rfjRf/hheqxfyb
LOMORHwL3aIneQRXjKy1ZYWrEG/oHgiQGC+TyeNEbHxCy6K3mr7pWHe2etHs2UY6gjd0BLi2eleN
7TSjTfmPm3XpmdQ23wxmIm1/7gHZuforlqqdvMU7kdwFro7k75i2ooYN63OVpXqOIEEFuS+3fFFV
m8KO3/v+qGZxVDmwj5MjBQoS8fu4RZNY+MU53L3ay51sA0LvLYE1loDdWWmjUE/XhQUZ3w4ZIt+s
j+E0j4cXVSoi8RCpsx51rNozCkI6xzZsb4jzOF2r6NGywRxi4Eic2dRJEvnEo4VtvkiiQU08p2TQ
HsLqIWGgvPoJEOOthtZeFfHn9mitYenu+4XlPO53acQd8rMo34XGiLLcl+EujxpzDyUpjEoPZex5
mRT1wBLYl2LcJeuuTCfHuwubM64s0c8RfX2kSddoqD9HeZvDRP/shBbM+ATGZaKuwKE10pmvYjBm
ivnvUth7RI+5lZyFfBfJz0qexV6JTec47bjSpKaeJ/nCSraKfCMOZMPBaSoSmlPecm/8jaUVGH+L
rSfP8r8x8/rBa82Byxgmb7h6weo7i+0bo9L/ieWKAegbIHSG3MW6t13GBInJ6WlmKZbRZNKzxAD1
wbIHCoDYMv7phNtjwPeT2XDGxd9MQnUwKyHQLk3KwxyyCvY6prYr++DiCk+2fEz2wN3tRiFkEBO+
kjRXJoAKUlX3ADPSq6fHqIxV57kxlbCmuv33xQE5JXDKo9EnCqpf9eGu0U4D4vnmrChbP8Jdk9Xj
No4ki35EdphUyByqWcNKLNAXJqlAn/WxsXiRG+FOXtpDXGBEko8tbbeO0KL9NCh9KVZvjCDO6Mww
nxBpUseQiBKrdzaWxPlSh6tVbW5nHVk7HHpNwAIfOYDJKhOExwNDaUwiWOUYYRsw36OIEQjL7zp3
P+H8XHKTc9s5guDfxNoPukgV3JH/gOlr7OUtgrzcPJWDh6YUEiV54JePQ5btZz5Ufvze/xlFQNkN
ZedigupCqAZFjdzLBz0BQtN+ryUDm5YOcXRQaWkDnMSj5Ml3Cf+LmyX86CFtTjNsXkVXLLZIsWrj
g2O8o9fdAfInf/UuGCKYsHTZj92K9NtpqQ6FjD2K5e7S2YA5MpIMSpIlnYYD+lOlO09sJ/BQuNVG
bpDT+ghhs/5ES+wnh/AKSNCvFv/V15Vwl0yG0NMDnuH+ZGuILZXbx09PqMrpVIik2wJqHni6PhEQ
CzIx1h34gz5DFv5wwwWi4WaxTB1fTzliiBz+XMu2wiv0sRysC0DKl71rpnkw4BlTuqTf3iO/38oR
3+unzSWH9F9GIzvWH6jLJSWqSQeSBbnlQ/lvzkAHV7ckmPXbvS554YGmB0+AtNGA9PrjcDSt3HR5
wnoLdyoI2QCCFiOZwVwjdhppWlMd4Ir4bTEd2dnLtgNUeRpdRCieaXz4Q6EO+u/4QTb5YGO7h7lp
GEqS62vz362g9/K7OblyVr654EXMvdAWs+zadRqVqnYyLIOaUIN1W/ETt2Xs3xS3xMIvML0YK5XX
9SoSZDomrJugwdhTgav7YcuQuekLwBHEvhXn2ZWkObncfGz6ZJMbh0El9BI4w+L/egWPmEzBiYFR
qHIcPb3XeUT8Odqu99AqvvVRKywVctgLB7ktLO5sOFQldP5eyuDhDw2ysm218J9wXiT6Q82g9ziQ
CnXAbU1WLuW9Hh2uerWskU5tgTA73vGLwCCMyqEjlYnVneG+I+RL8yURAZiHrgpbbtJeuHmlhtVo
pL5HGvjz/lngkH5svQ6ZQTa8aA5UGCDOyZR5fJ05Gjf7aMnmQqU/wXdHO6K3qifdzYCUq2hM7eoA
XsAFIicztrxzbM4KkH5GdGxzLjXnGEKN6GaSLxmg+BKAzpdNI2azla8ruhFocMbTbn2b0Dd4FG7h
j69o5S93h7GfbhKEpHy+SPqvSLoKmGXI+lrjAsU0PHCV8w/r8/4/M6zXQKKh5y1kCdJWjklwZj4N
BrLQU/N2DSuopwah4NR8zXTYH7Ng/+o9QnP83saHKNazEqE9Onp0m4uu4ra8Agb9EBbYw06wG3dO
g/eFETTtRVnMjgG0Hk+I2dauQsxT1b6iR4IwJhVaWP3VMVNFn4KenrxjvvkqgiUB6tkbfmgqo0l4
XTO8/QC2c87qO2fAQJnmH6BNZJgQ27jdwt5TDVRcJ35nq2IKkqAxzEPpp6fmkfnk9M6CBwR7Ykbv
NNGs3czQ18D5tweVymYZyxD2Hy1R5T7TaTmffN8guQvixFlUsh3uQeYBObZy0YbJbmV9u+4AVFvA
ewBBB1s0nSwAmJ8sMwHg5Oq/K7FMrZsRYfKotui/ky+o8bx171hxmH5LZ1KoSAwlLKqHoeQt/2lW
0ekd1/rscm4sJAbM2Ir+eYw0CRoOmJr7wssOFF9uIbu/Fttp7KIAO3nGofe0husT139e8/jFrxSk
gcuKQoD8RGrXkTn/EUQi203y/WdYQvXY+TGBVEpZ6D+pa2FSNeoTSFu99Ot7p2JjAa5XWsqmLLS6
voXcR+5aixef8YBrCQnQ06Nd7bECGFl7GexCv1a3xrEoC6ytbJQ5ecmHZtb6/YzSkJzRd3uIvI3Y
TINq4cYwPbCNNP6RaKooLWdZlTVZX2KDS1oxFkHTiVk3BW1ne2HGiYEDq1uPF9A3GauOxjtTteUy
js+9Z1pSh/AmKJ3b6zqdt7zVBfXNVEWrD3s8rm+tmvuCQQiVBEB7spo/m1XStQSbVxSxB8xcOF9u
Fo1zJZa4HjIBDsV0hA52+cHvV0Er/3TYuZ0mPCZdUhee2k71ylJPfcTf//NErdJPvrnmp1dTYuTt
viFTURZwDFXTik937MKKb+G/vZ1TcX8jF3Yj3CVqlEaVfbFjOUgPnkVqzdgizke9rZP8lMphW+qu
XysO5FpILs5TYQ7NQnecFfzxt1/ElCEpWzcIfdSz8/u6iSu6CdcFPw7AZiGmniq+UKYLx3Ln5hfx
rtIkIdpM2DSUYykxsGgezPEHCJg/2NZLdHFswTksU3v4/u5M+MqXY52B+Fwjd5Qdp8IHfhsJIUb7
eAt3tQ/gZNcN/rl1AXJtomCyJRLVuZPV+xKTrYNr3WT/UajqyRnEOI9M0qUcQJ/Pyo9S+qFezPvh
do+mHdVfQSnUBWTnf92cTVneHledSR3Y3L+dwhNYuWPXzfZmEreWzkmA0Dx1FgM4R3jFJ9ArbrEE
3121WiLO9RKu1bRbQvWXm6kFU1yZ/qtLzdt68OjY+AD8QgruC0B2kh0X/YzDCd1EDjACRmuWU3IY
/FT68RXHpbdiGE6ASc/05BqhXYujtMdQuvI5MYQVVbBJl70Q/TVofo0WvkpBRTmfauJLrpm0IuWl
Av/8iIB05HH3Zi9NgfqgvewO5DIevb6DsA+VokS6romcnIasuik5ZHTmoAZBM2pLkqNwAEy6aaL6
LhxdLfl1TH9G409F7nmOiPJPX+eccun4LRWIwecNvoU1HVabtbdkipilSoOciZ9ZWcx80+n+Xlrt
ofLLUMXVnm2vI9tstWYtzcpwjQ526tRduOAkBJmF7fLoLFFf3cVJy1x7rKmXNVinHUZmLoMAOKu8
cvDLEtzAadt6xOLe1NAg0WdUfOe7Q6IU+IRdY/oT4LSA+JeYRBEtkmTdtuvqHssF7/wtKY1033Wk
srswFGVE2ICICjlHO7TIJGZx7USQYaBzBx/AUbeTiCWcEl88Z1V1ZCNNZeyRk67GtCqHNFQb3luD
r2XwqIkqo38Pafddjs21PL0mwtB1LwNu0gHz2XRW3et7cN2kbqJkcWZIU8KL5zqw4yo5wlr4y9G/
H5LPFQ9Tt7Wgcn0UTQgG1XzSLsUtgvBTapYyWL4XgiER7UbvKjwhecsWGGVl29DrIIurghGUFxXS
nfw+ju2Oes7PVw3bW5wxH7lIDfWuFkqdjtsOKdKr3xglsfbnoEgtyxRdZHCssLEiwBbVbige8EVH
yF3g2LxmjxadA8CHRgGygj/vAqlMlmakoPQ2kEwvb8b88IA2tiOZ70kYamRQyPSL5UbEjJCH7g/9
3tD7JQJNmGFW6KQJzyO9KXBUhvcN+n9Om9AxI8/BPwA67PH/LmSVapkM5RB8Qy2GJe8C4VUFqhee
tdUirHG9adu00O5Y1llRnoPITGmmJaKhNIgUF5755oAkDCDRWoKERtQxu8IBopGUbXpTOaHssJU/
UY34eDFueAgQVLGhUlvxZv9Sjjd5nTxfLcxprpFIEHXXy+2oaOTDW2ejGdszg+zeht2HqeX3JPjW
pP+lEo+TbHnNjwf7iKqs/G2tDGLb1tjSHU7ZbW7Xg/KB6u4ra03kKDfeJrNWBm2BWTjgcx2gZVtE
ETFSaPsuM2kOBySawoJaqtDT0tVjZvpElBL5E5+1ZfVdQVkOoo0MFDmtAkK2BM40X0g9wtibkv0d
Wws3FxAeHjn6oD+AQ8vWJjsRsbjIOPlvcu+Ud8cY7fn4hbb6H3ohbxi41BWl/NN7derG9akIg8yB
be6xyaMJ/JF4DwV5zz488wTgtj5PxFC0/tV2vI6yetPKrCdEWbRb6B2lYLCzTWlj1pV9T4cU6F6o
wGWMum6ZoUOLLCIJEgTjbU64ecOm+dECZZ+hHWJY0mGqjeec/09bamDyTiWinl1OZTtAYDvP9OvT
BiY7n7oyTxUeNWOkhJUgcSApYPvt6aaDkUteaomMSRkULnl8j1Z6TjQLzMVv3rUtjvz+FXSe+OJ7
gSBxG8XvLmidwjIOLVOAqBcfOlLl9XlKcEKrFpO+DQ1jPJ7bOumXjkWwmhGWuG6hBx+XsBvWzXCE
2mZJC8PwvixdMRdhSBC/znx3zhNNPwoR++4sHN7YqJBngK0XMVXDJ6YyuCILRe4dyuKDVLfI5poY
D3XdqwrYowTazUA43V06rjSdkW2WOpNZ16DH0T8xfhs0nt11l1uFgeosXWsiVAnR5AFuJIYOfxPk
5JmxRdq7/dDhqahdDK0zOFtWkAi3EmPfUOf3Qcafkdvh7Gx0u5Zuw5tnqtI8nUAeMF1mowUgS+Cj
21zhAbdUZAmxzuWOFOh9z2COAS+ogYGLoQpXeKXc7tT/THrwws0ToQtOuF8T/4gjoagpbIE4JQTf
yH9NftF/R3VaFq886CKFXS03LFJmfekNEVIUccv9N4d3ZRHFtZvdtDj2ylEtm8jWCUtqIbvRAn0E
osYI3cYUbRlWbwdtKPc3p3C68H3/3POYGnXEtm2Rsyt1kctiHqfUGX4AFt71U6tcYpY8k/7ySmud
IO1yLIz2W7AOCjniqeptljzbBbz66aGe+8T2/wp+1BhVTzC5b3LZDN73RYS/gnMDOUl0u1u7xFw/
Drr3QNEsNiuC1KedRLbI/NAQjN9RTwatOf3+pCgqBufzu0bpOyryjs8HFJSlh/B+RsQAvewUszna
TR0t2FQZPqqccN5P0xhPzJEx2IY6njB0ZT8h/B5qiLBfCZkWGg6kudemRtEa8c06jRMzNp/BIaL+
Cy+nSCsNRDwv/Y9e4SmaPMKyXqZeSmgc6cZ+ErU6oNCiHJ6lfzhuOm3GIHHI15D5Anak/PYstfkE
5efCvzO3EC5tjoW0ZIkulJlmhgvOBExJ7wo4AdxzHEJu7sKV+2cqjQWcfigCBTQYYd10F502OapO
wcVQTTXUx7uds20N4ufESRyRGIy2Knla8ThAuD1fSGzowSwfRy5x17UqCcbpDv+ahd/IjnyICASs
gaQh66tRYQNVDUQ9qc8PIYbTiHAB8xx54rgn64mHY8vL1vYjg+/0qQbIMSkm/Uhx+zhcF9xrIPZo
6GzyapvyX+sJau9TwHvxWuYIPH7StgGO9PEn443OPLJU72mXWvA31rMBlxMfmfHju65AzyszY27d
7TuAKTEmchnLCbAz5EqI3Q+tI2T+9s+a3Vja34cHJolOjYKS6pf4MhJXH6RBaO3GSTpEhCQj5Su1
UzodcgR3qcawmSuzZ3mMz7lkY1lh6eldrUWKv2M4J4WTvpoWg7EUjPML0/mc+PM4l2DjN6qk+6Io
FgiZZtw4M4NM4Cvl9k2/DsRgFYf7HDgUHMKw6jyGzMJyEHnlFcEKViscYN1TCW2UcH9jGrEQS9VU
Yhlgvj9Q8xG7eJdp8+LWjBv4qu1zNTW/eu8W6V8q9HOqhfQTnDYWBGBLYblu73wVMoJo324F6jXS
aFXxBjxtUAQepo+A84H1Bp+88z3rQEqckgbDDt/wK2HKfuSXmD+CbxNBuF9MuEmdLvSx04XRbTb8
5eFoOtzmlcDX5kkPVivw1Oh4vaiUPpttswcdewr2EgTJUuRN36TVKee6oBp6HXDUt7s+twqb/l5z
vB2WtAZbEhQzYZhyDqTpjDTbdtp9t0SqGggcS0ZKhiOJY59t/uXQQmSbXP/ZSbII/sdWN/rkObqV
EJWf0v6uNPPxiUfE+LuapfWAoEJVo6tLlpPbsPT1qJXJfd/vwnPGtQJqbfAOWfmTAGHfYl98bJEo
LDNjT80P1Gzep9uzwDfkh/FnN0e2F45U97y4clC3RgXpzZPzp/cUHyggFiR2pKKhLNGGJpfEEIAN
QKIDHoS1SBQfyWCryotrYJuIMewjCbu8odedEXKW8d/UtOPNND07vzt6O7I3ULgqM9GFPEyOfolf
rleKMrMH490byduzQ1zxQONNRHNfObUsiwaTRmM2T0lqI8DDxWwz9ScyJ4vWFORM1+UrpC4ZJdbV
DAOgtiQ+yqx+iJRuKKQS2ea5RmKbcvkq5YDofuutrPqPykZDAZLmbghFvE1QhnVM2iYKOXxH2Ge8
lc9yFWp7Tx+rLGcvf6sQIGmoWsB+ffU2CP8p5XPj8NcU6J+VPbZvNBLzdPJXKVFm3IBg8Bg3iGwt
w/1iMPHwzfw0xrfecuj9Z4mS3rxNKwT08HsNOUcy0Tbbmru3rF44QubnLqxy8MBqoE02l+umsxyc
c2cxPVne6ZQjCKE4D6j0whJxzskyqAe9hq/UkMPmjggITFlbAw81yqDb8NUvDfaRMjt5S+TS9E2L
HV99wUdRRfHohlIk5PAn5mECgCJuTpQ9PG7GTb+AAgFTMend0W1oeybRa92TWfFNJjk10PIUgU1M
KGbV2N+/YuECuHsMf2iFIC1rQYow5qptM62Iw56qEDnSNhYwjmoYkbs2b7Y9YjYGtxSlsIlIKZXE
XEORCucZlz18E3SU1U03Cjjmy9hZiQdSVcb684d8l/2xTy/EPELJqYRhmSHYxT/xCbNmawCedoF7
OmaOdZQ1ekqUfvwKMBz8l50byBwfXJ1TazHxqfCQZzVWi/x8j6pTwXF088IG5Cz8trRMAKFRE1qv
nvRbBr2SyaIL/xMwO4vDFg3nu4iILz1U6cyHx0Jrp9QH5X4EbcQ/CLmZ5eavCTbj+rPH4Sr+wC2S
m4z2WvrL+ssIp+djlQbfa+1elPA7kkrZDVdeG90DgkdDDwmLXVHab9O6zwU76auzR4hHR6PNaF9T
kN6h+iaNPwQ34TOfiis8RUpNg0PqhqCg/Qr4eqEGI29ZoG1OuSCPUzP0ZNDR+RdjFCnt2gIMVdHy
GAa5hX1EzQ+d4I/Gt9ljCfG77x4jIAWO40v9OaPWhWsRdHygQt6YTGS8Q4kOFctTT/EgRJkai0c8
m2EXEkSDKJly2bfX17DBCIyI51srv3UvNW6rc8oFvf9gdilVJ57+jC5UZsI/3EEUvGYdZEI8YgHi
E7eagF9mS/usS1HOUUhX0Ucsag6uDn/lksrE/Kr+VJMhT8CqA6omAPRmY4z9tasU23eY+if16mGV
iNCFjFypWvftTIrePe+W4x4244Gn1BzA5ERwha1ypZax1PsOoBf0PEL/7hyDDswozIbE5kbmFrnU
V/j02KkQQ+1QD8tC9tm9FIcWe+QfEHAI8Tp3CE2m+beWJOYDOhJrS27s5PqCqJ99833nI1dPhtT1
nnMhg81bROkLZncwPvoixKeNURLHFAg2jffKEJn3z7lsqiBwjvVF+R4ghpoXCcXi5EzsSze1S7NL
Ht8osZoO045ZGPOlOOrnPS5nly3U8GMAvoU33gU5GPTdweeG8ULbFToVYxon7r47zhgI65l2Vscl
J0eWkL5SaytZUdWG0Nx9E2ThcDQlKDwH0uiRINd7jCaLRosayLYcYh5T2LQz+ywbWNFOgTrQkSdi
F0KgWcnuZUSu1YGqjumZj3T+O4MNqiMulm4QNrwsZKp3q6uZihOoUlhJ2y+y9V4k07YL6e/esFQp
1sr8WVjPSmt6HdMIDekXzKZzic89nAhrch9UMLD+sRx2+jo8toymBr4rGZP/frSf8WwQmHNMaMAS
qWUwz4nNrh/E2IVvsTe9pEVlxAPdFJZguloxfb/8EMno0KjCGel0r5bDOnL1VRWoOU3k0DTt5TEE
ClKDupkTNWN+Q3Ka/1S48TM4OtBr7ue8kZ/wbfIWMolqVWexMq2ipKuuzE3Zg9mgfOwDhsjSzs1x
2YAqAoLRP1fM4JRS5iRglAWHfDuK6ciQp+FBk/Z2ISFGddGV2NFatcZQTnTjYcBP6K4l3Io1+tL9
RE++3L7sArZlLtcr9mxQuV3QqxMdveVzXoAmMyRFu0K/tVhtNyauXDrW+X7mWVaFXujcqvpaWduB
k/wZzHg0y0NohihwahUNhm/J0hF6voBp2kGtzUR6IdtSO6fxs0GpchAv5NrPdnRTwTX5VzrgNGzm
nj1RytEyGfA6QxZs4uhH14vujGDrGhtJNuFx0CVDXeLya8sHTJnnkM91vPYxfkKJe8qOy0cyu9om
Xiwse4Sy9JhOFbh01VaNb5IJYMQ3kwr7tjkw69VtpPNBelYhJKxR5MMGwONugdl7J4oXSVEBi6Ih
u2y/cCPxn5sX35Ew7LZbZaQJPj2n6SiGhVaUdpjnkO7D3CBh5KEXtuSNmtgv4S+FcND9PE6wqKLz
19bCVIklKfWoFb6DrkDFkcqvAWW9s86J4WQta99kVUhgY3LLtQS5M0sh/1rWG7hqjexWUqect3I/
Jsq5crbJDpVSlG7RKDyptcFF6uma/6h1yc3fALun6F5ZhlDvg3SwwPJY9uop/5UhEQCZgiIRyeEg
vuCtlkL0DiFfHaJpo0f8HLVwTF89r/upfaFixxed8oVD0qYhLLzoWYxWhBj91jRF9mPoF/SQPMKG
GXCvUdAAG5chKo1VAFkg34NWKGowMYEjgCZJT9TqiFbHoOBV7m3v/N9Q6gHJNWfbbUqXJ7QGO0AV
VelPojdfVJ1yMVWsFvdSQcA0n5T1RKx+xaMFPIK8TcduESMqSvn/yi0jXs1JUoQ+VGzdPd7QgktV
dQ9eo+kcFk98UQGhTbFiNL4/Casty4Xluqf90Q0UEK+eevbbIBdjh1nQANHFG4gGZsTMYaVkyvXR
Pt8+fxhjm81Iokvl26ZgQwG5oxuDDkINqwstqDTEbFWRWJdl0lNZJgOIjOFHQQ1NQbOii4yf9jHY
Bb+sOZmsy+sTNAhvTFwukideCT6f6tow25aSre6UO87+15A1TX7+QSUBuk70VZpKFpLa9ACYGoqJ
EI1Pq+AbshPXh3jlhEJSgMvoJOW0K81JgoLkL09q6aHdQ8y7hpVi39ToONdVgntjPSkPaJl95uiz
kfAy8L1GtRtU6eZc8vecX2tpP7fX1Xs8MpT/ZevOMGO6M50TEM2Tmd20uwRbrEkHSJ3Ju9phD0vU
N3OwfCb+ElYiqEDdRofbkU2QOK4ngRdYdqKBPS+N25klS4QDYtnRc0FPjzNv8DBrNfTX/J3PQXXo
iYrYzuIC1S87eQhECX3wnlV0QMYiqn6hQN6PwXCC4V9qHTDuVOZsD+o4X0bE/3JuPe5+QMXZcRSz
1HscuIkKXdQaNTvuaZytOjfqDYfXv7FKhMJWUVJBkxUGM2rABJFX+DDFd9O1ZclD8yfjB8Nmn1Cp
SzwnHaed6u6ehipMrk5/P0V5GEGNei1KuMq/hGhJwQm1XbFKuZJLdAXENUAsMjIDFRtd4Pxoyobv
9WEbg2jCQSsT8Q1Cmm6gJr5O5vILzRWkDi7fpK7qCbsGbKeum/p6ilPxHFoPC2qcMfDEuGkr2hB/
DPo9dGuzvCZeLfx9D73CaRwETUI0qhMkSVd9XaQfZntATI1tdc4w6WulLzCrZWkbhBpE+iDmrVPK
NdHt/Yh0l01EBMybyZpGWtXPqLtVw7BaVl+qpXSikJskMbaLt+3H0orO4rwfO9ne57YHPX8THDJg
iOdawluO+9uk7mSuBYPF0Ttx1SSSRLJ97GnvPMtj+Tpk1V+W9uBVLLGOZ8E8uah2ToBvDCOpN8Zp
AFHVdGVlGVFJZf38sZpmDDWTDyOctiXwuSBpGrQhQ06ywBfxuy6r3yqFC6ePX8OqsPvxrRcKpRCQ
q0O/wSzOHGSRtr+XPM16XfJQUPtV16HZDhBUThPomAIx4Jr2NjssAOkc4LWmt3gU3g8HCR2p0c2u
1dtkt6Jm3li6GkSqlzdmNitC3iMQBkJMS3NuQMr2Q5vFxSFQdp17PVvp5fbhwuy/i5Weg1Y8oiwJ
Df3DUNIrngZ0D3cqEoVx9NS/SJvz68wT8hqjkBGgdZEXVOrzG1eJtfz62qiZHXVrb8gJXlmjbuA9
dJDsTCkigkRwxFLrxe2FGQjeUNCK6fZV4tbLH2WuklAcKX+eiXLMuPXjlRjDhwMUBhFq6nuXY2t3
Aji6Gofb9Y0VVL6bdy7/tsLAJvd1Fe8egmODQyTpch6jFKqkHUDeuv2vMjhl/IKqU8oA2zW47PYT
6hu6U/k8ZY0rOPxar9axA9LvTJit0/coNZk65nKZpzb9urmrIEO1piWkzZRsiHvUEyYdgOxbPL9G
O5NcexrDzB3XBxhaZddCCwiHA24tTWswE+p/Blx5jEKKNpnciTva0s9Fn4h4yFBW108A5QsIXtj/
AUpSl5TG3izHcK9yzQLf+0xoMxOEddUpz5AvK5Ply8p+PMJiLWTd6FR5cbnncvRXuxtxUfE1D4oI
koHY5x78UsBzRkIKCvM5nfSWREaJxohL5UDi1I9W5hqgvuWYcPmzno+b7kUKbFGrnp9VLzulwbGx
x2P0PhKvD460XfdI/8E27fQEwlHx8a/H+Dk8A4bYWSxSJKsgk6/jJT3Psy+qLI4uxXNF+aKAnaXf
I/jmKRdOUeeWnOXelJL+Tv+X8RzVu9BkV/u7zyzFM7UN1I2yeAEeXpweRfazHu/NExMn4X6bVnYH
LZWr3P0QRsN3uMB+RiwCKv7/8i3xJiBNJdGHiCFYBRG8XGJk2LRJu9UTyFv9lPC8C1U9FN4dynbt
NiQYqnNS4GQexb9rR98SzCKrwIlCVPQzddp0HxUPX1AtSRzxPdJKBfa5Ryx01Zjngx04d8V/Efv9
QyYPI9nAu6AiV+Hwxr5cniPumPdF3PguAVkh/9KD6xSfb6XKXGyiZLatLKDYlRZFIEFmpKmjISaT
eAQ6eHGrlZSYJmcneXy00GFLTUS7O/59/2AXzIYjCQVbDPC6N9zhWrTxqf/31mAVSROFlHXHnP/H
oYIHN81h7gB7AAQPGVZyFAcsOeCe7yZGmx4aueBUSsU7wGq6DYZknthB65T4QcUAo7S1nqm6V9G5
0fLYHauKhuGJ7rAg37K09G7fdHeSHomB9YLat4e+5Woqu4V5sJWoFE2Hx9SPOSgtWwGKgt5AsKRm
Vwf5Ys+yyJ3BMqjFOwvUfb+fTLP436efhndIAYImMhveNbpKEpRnXGVRYqjsFmDkViO7lN7c87Ms
t/anEqiep5hcp6wA3c2EQoGrxEkqRe+P8o4u5lzisBlAXh3/1D07SS67dH3CpLl7kyg9d+Ro4pG4
h5f9ga3kOsB7iJ+yjXct95rL5PzytNLSdRV3XrCt+N2VPgXlERr+jdKwuiGousBPDt//pLdP8Dss
u6v69D//hK7Bx4Xf+78pw3/QduKLVKCubvhJ75emLBW+RN3iuTpJcVdBnkaYigCuZD5U+aViBk5M
UbcuCuSAtVv7EZqo+cfIV3IF78uY/Ic+hc8TMfSYRrxsHmy05YRkSHRJXe3WH2JRmGPtqpo4L/UN
wgFjjH28sbMriT/JpO2z+OwVEC36vm9Z40jZP0e9oLx23cR4Ua79SU6vZrAgSqXiQiu4bKqqHKMB
tq0wDeOURDCn8oiufQu1Ev8uWN4HbxH4nUgDa63YQbRkqYQ2Moci06Z5VJjWCxr4VvgyTGdxErGS
y5dJ4bfwHyL6IdPRVhVBuAo5+pm5fHsARoB/avONxAO4u6MFeVRSMRHWedxSP+CRo0xZcpT1bn0x
MKBieQ+EvAbshDWHM/Vu6aVZKOp5wUenFkxiNM26WVpRdo6g9/rdlsVJL7tbbFkd/vBCGD01Tl3B
/qUOI3u0w0oF1n8xd66nnVpdCNUiDwIoblS4yUKFzBIm2f9Blc8c1VpdM1OcPBE2NrdpK4m76XMF
miXrq8WEHOTRMhuMj28QlYX9W3P+0xCHLfkCWKJHojzc32ahRHXMNuUGsplF9G+MQb89tjpOMFM7
fnIUJ4/0ZtvOoYPjBzf5MCMHAFpzLjPkOC4vPeJ74RQL7zrXWHb2gHwOHec6hwwsZTIvOhULsbNV
OfNO2nFV2Y7HKhKVzDKSS1DPyPOallVWOFC7oLvDE6E8TnbnOeVaipeC0Lui8Yt6wihJCGic179A
DnD1QNvjecOZG2W9rhaXgwhk61dopU+pv62OfcFReGxnGEf4KdKLjfgA/W0uz2tTR0IIvuKKKcUd
cAyOMNydbMQJAsRY7BykpgUUxvN3lr47XfCNh8rY6CidsttNlbdc3RZsBgQwwUIYace3/mk2oNeh
74zqHqPFpxfF5Y0nQG9tDATtYOaFWLV4oGZme2tKpVCVG+9lwz5d6iYTfyNovw5qM9JX2WfLj7kp
BjCUmnx2rCsdl87s54m9cRW2q5fw0lgyUQ2Yr3hG1QdUi0zKBMWOMO9wJmP1Ax1C9jjHp1vF9q3+
jGUbHcqSWkY+vj6eoU5XiLMicckT+QWI9iUeAvHEtcIWMSpRfIXAHETJ2x2QgLvGFNoaugN8dH7J
tPyYhrPVSiqNqrAzZTaoyfyufaZpUUWEpL6qfTkaENH6R+jxyV0peqAIzhPR9FVMll9haUO4bIfp
kxKm8vVOaWlMBj0xAPh0DusNWhuREKpQjT0MfDBd9wKX4ow3e5m3PxespK/8Kbn70WIWLIKKsv95
CVQIvs2ndb62agIzmSW1t0M2USv/iXFH/6ibqoyzrrjwoEo2Lg+GTrc6fTiPBBsdeFHsRe87jcZ9
+suv7XKrHOIVxLnjoMiMJIYTDd+wCX8LuVSkCfK6a28RK0DewY5HQWXyp8sOnvfJbWbuER57K6R+
U8WFi6fonn5Mh/ZSf6o7dVr43V6cZ7ulcwY7I/s53Uk55Sw507lVsG7iELQ/yaZcPUDVkfW7Si2i
c43d09creheQ2wXqpHDVlag2V/2nqfCsv3bPUAActV45tpWl7rf0wtnC+uXPx4X1hb9dlEogrvUz
fWEIt7Jxed2pj2DrlBh/yuPME+uQR6wwZG0F2/HZrgDExpDC6xwuJueukeNNvgyMqeuxAIs6LNEM
058EtQm6kppdlQLCTaFLpmRbS87QFbk7ZCDEAWblYTQYwsDgAOf90nVBOEygy00yIfXfVz0FFfbw
0TXwVmnP5osgcc7cYM8Ym7e3fhsgRvyHsbGU/Ia7giIEUSf1uGGVwTRij0IhdfLVA6eS8RGVdfGv
LrnSHe5kbqAXqyGyzW23jiyzGeXMPy25qA+d4AZOJCMFHAU0pI/qNppu3w0/McImZU5GFojxwYU/
9FSyNckg1KARnYhuIAeTWSC/AEHZbcau9X2NtgyEEsBCFlozfSbOEbg/bLRUWBkKbM5EDOIhZapu
hqFE4KEWggPoH1QpdZa5qWg6uqgRIcoZhpGk2gtxfBYy/QkxzvFWSY6vDMr8KAvAtDbHc1dUxe3w
diJNVV2S+VdGaAtdQx4h61g4E0h/DISTJVxAbeUp8ntn80c6AFQP7dkKUXgk5GBrLh2GwnOELK6j
jsNXB/fgMHucMhMkpPKF5lZF1Ps+1STbKwCzSbjh3QRW0TONYwvvSqvi23s5B783zWccBscNzdCo
9rfFjFySnNzqYg1a3Z6OS4wjs6HkY4dCaWLqU/Mr6sb5C+F1e4Lc6WikrfA2im4fgWNL04x88TKa
xD52iQq6xj9Hlf6yLANui9RfppYa6TvZQqdMrfmx4u8wSEpyJ4xVqLkkEaBIz8EdbgD7ux0VBGsJ
jB8cuT7323BxUvKncnVXnzNZXmxBbLBLbs3WxGKvpZWzrlGA8OvMoAB3sfsSmlB3oRqbJYgNEWEU
5Zlj/g404qqurPIeE8G8anHQ1+Bi4VBLHb0CT0QVQTumJ06PljSY7T6xwSdZESMNo7sRJqwhHaTI
opPaXjVltjLg+9hmc+mUdd4uW8pnpKukqS3nZaSjAl3jFuzELW9zGsdXimbUtOYHQ5GExamj1fpR
yGivBkh5t14xKfDP7UrkwI06gOpR8Je+8LuvUwt5A8xEe/JNrh7ssnQ+Le4jOmpuy+FYnnGwWi81
y5M9Y7/O1XLFfa1LE8M3o3wi8iMYDTiO4xmaiinAJIVyXBlKC9A3pfNoIVoasbzzdN3MsVXouEpY
ve8ZKnb6VRXlehdriBgF8rNSjpdtd95fnmygOKEsb79hoK0mxiiMFUV7/yJZOvNNWF6SlgQ8Lkpi
p/evafEhEgNoUZBNNcXzmmX2Lbnc+L1OwXSlcBGlEpfHHomznMom3D1wzrh3sgpPcwWeDNzt7Kwj
yoJvFJ+1ZkU8h4VEdh9hN3x7M8pfFmjmu7G3530saWCI77+yUt/HJUjbikoETfusgdkTZW4RbiAF
LJ2+G65GzTeDUKYTihYjGnsp1BsRaEYwqfNgxpxdpq2pYaGfwDDBgjBYoLmZ9ryHsMZF5LizNLkh
jK1kiZKhNhZsl2zALFBeYOxOLlrx36v2ABgy2Oxf+cj0DzUU0vEOeWLu8W5JsxcdtxkR3JokMoZf
7BGlg9qFTfy9zLnJ0c4sfGdvlE9PEJGPWnlayzWhx6qVySglf32Mrr1BalNRW8x9yAE0dQCglpdK
szMKzvAOuY8QtlOUznN6mmidT7tlqIGNDrSc1ehAqNyXS7ZpACaNt5AcUyKLfqS0QqvOTvOgDiJN
fsD43J8Klb9JRSq5eWdtDOt8WtmAUNXYxXIxRorhOQkPuJw6ajnIbrx1u1U5MM7JR+zGtgvukYOO
t0aMvT4p622ee32ZxZRnA/p6/4hAHaYS0+C4ULfn/1NJcyJ45p1A5fRYAHNleKjfI+AgNMQgbl9i
iwMQAgQzj0jF2OqlTA6a43QcrthguHYfKWkXNJpeUDT72lC5LHiDxX6hvTB7Brrwp4eAZq2FOpVP
QdAI7GgnI6ovyPyCR+457ZHqaFEzPldDkefDOQRLrR81DkRqx2ri/uOKr1yRqK9e88OM/AndCYhf
of6GY7BsnV9Eyldym+YeziuewHjaVLTseXjNXXQVY+9IifF2pHf/dSUDGkbkYgYVqvRU/5OLoi72
769SUI1D4Uoj8nhbVcEkF8k6vcYCX3cgSOaXGvCqurbC9qLI9EbBFBzuVBzGkhVFYO0Q8bfqOvqS
308nTr5/e4imqQevfZfU+jcWQuz7gZKqGn7GOOhAi0AckTO9J5LXjlJgptZKFB4fXvElPWp34OEt
RngqWcdEKnO0pEjPaE2S6h8+EjFhHktf6q8GR/q3tzADYhrO8A1FGMjYiTFIsZc6wbwIEd4WA+CU
KpxvfMawTnJBDKitjKukFrkQLpzGk4jK6ceYkSO0zb8e9EIGqA2GP1igdJd1rW6qXb9AW2h1J2Te
4vfyPmVjeWFELobgc/vYmvOk2du3I5H4DS2bnnQx9hZB0Be4Rx/tp6REyFjjuWdStc3JfBFfsxoZ
FyN/Dp22HVkBT8LtH4zB5XAfxwom7Wt7zQzd6lY1lAtKAFsw0g2FR2F4FNRc3T0sj3DDLbnyR0U/
ibiCd3l5fB7FZDGaKiLUo19/g98KUntmQ/V2s+gm8vl/YCLmIHZBePzQUpzKXr7go0nyrjJVPzm0
twHK39DNkIE48bgvsWT/q5XM1Hez+zlIdsCBcArzhnnlZPoMhm/8pW/YU+SZOKdxkRN7LVpRJb8j
z8fuxS7bCTIUGjCmjRB+8mZQ/qL5AGKVPxLBcKfxtyZrVpObqIxZ2nBaBOPRnFAL5s3+08pv738I
kVVIDwN+Ep4QQVd57kFcBhClusf6L/A9CTIi4IsPBCHngvsSdzYbqHFsABRetrpvVDiTqjlBtGL5
gPESMT4uNhgeFWnwk1hY0igyR+1fywO73Pkq5lkRzfKzPrvYcWxGmn4o3+lcsjSisZSyYZuPiCy1
/I3cn6G8cPRmqnAjb3StubXYRzV71U1x3d5Hn8wxaeS8lPF4GTMis7hplau6/PqYqL4POD+C8iEA
AoR3ClCCB2nHwnDutpuI2pW3nj/QSiWBhA/gdCYcK4PVf1KL/Kw8tFHnVcIGh9ddaFG7V6VcKCur
BZcg1u3kvPTmufIMvGY7JJsgc+7u+twRROOoA3vAXbJBgaMlvtGyfszet49dbpRIY7+pTlimEAnS
Fw++zW6f7BSy3KjP+a1ZzVrjkJf9sjU/Dl0YCxAtnIkpnBvYeAcmD4L6p7ujkMyCCAEYV1kIrFNj
heQM1jBI32jyU/xKIFdcsecC00S7UpTPsYHWgv4T5IUTWGO9l261gfeofvWmVeNfZsJlB3CjjJPI
7O0XknC+jph7j6S4WuKwNvw6ZWty/2XQ/4CJPd4lUbPfla5lJ2faQ1DU0wx0mnefwRC5eyi2u5kJ
W761t4rwqY2vnfpQVoF+EvbxIXwN7C/LMuPWYLgBEIBRFAfG2m/7hq9IrnFu9sK2J7UgAJZWHXMZ
MrVtKnJjoo5b3yWVAkOlrG+qqQIaUoZ2nErQS6U6o0SdyHLFPpQ9gSoYu+GZiiZBI0QRZ84YF/88
i0eXz0LVuijcuDlsNgn2747/W2PvipMrGunxiIRbTfeYOgmkMmh2laWTuCsDVM+JAgf7YXpOrMbt
hAHtYVXIXucrd/+XgaS5xgcdton31ojpby4Fln7SAoPwHTS1bVFrj8hLO7aNjpoMOJPilJKCs3hO
ft5wAuX83wkgvB+F74DyyPBgOEwuUHI3lTjzt7F6WO0ylvmdbyXuYRw5S1XJ5HqsDRCSVPZDo4sl
9xqICENt3KSNQHSGrMk3tvwrzi7Vi83rAomJJF1LWNx89V6TQ98c/9fUFEV+MprVAxX+TaXTRyt8
25ye+q45PiOsUrsJTXxFQ4ikMCF7WqtrwCa9Mf9FZFhmbjYiRgdcaB7zzt4pr9QaXWli2gFLZ6VG
6lw+jAlBN4dzYS0WNHuEbaRPG9D2KdkWqYwT9+0a7ILOecgj6c0x3toUCgPLFAz2OHQC80v5QyVI
4QD8PPicg//Tamoe15S3uF2P9eufc2e2rqsz7IA8x/SplBJaWw+ylLwrGPfmXkCUT4PJ/QnRHaYH
3kWfq3PQXISG7yNtHr1iGPGfH3p5XdsseRl2eOI5dW9/Qt0tZ3gyYOT+sLPWJcTXDMtE47OKZ4lF
m/55AVglAZPMIL1kXadNMM/+x2/kZGOLIANrhssQunMJqDIlc2Ks6jr2SrvfgyHmXkuYOz2ZuWiX
GqQ6xJW536CbxBmFyMPrgrm32WMXAnZjg1YMoqm/7iXV1TQIJjDRtCj2VVBi2jEUYf/fUbWhNe+p
qHch1M4AkO1x62dyMAIJPU/TVvJUkb0qMwD+Sf+/rAdwqc7pVY6UdxvEVn/ieEB8NOJdm2GtGPBq
z7a8rITkG0SG+cx1S20WfyACaPzas3Cyyb6p20FUSkjazOM6S/ogY2sW4jmCda7EVw4m7YUQkSoz
mKHTlTaMtHgY8HXb+Do7HjcOfaXCaXEaZNZ7SyOdiNGBM39wXx29SC1Z+2sGva3MH6VGWs9pvZsC
tu7aTshEOWrA2agSjBtwkrXqV/yKgayJ1H7OpUVHVPWyTMIlkERzJfb5otldzMN3AJFrALFJxj+w
/WIyTH1RcDI3C3I8hqKB++IuVQ1OjQ1IGVCCz3EDpNSJAd7HBf8PVikDrDglwvT1wQHJ225k937R
qBwJNA3da7P5AayBBdC56fZyqvfe1lHl5dzuUUj7UdFlTfYJZhhOGF4Ej9QL5JOhkdU9RsqVO0rG
c84PbkzB6kMvDjVDvANvCOQNTOZqvEzukBYmfzgO1SQt7Nc20Ke+TV1hMzl9z5YP9sPMAfB3c5R3
o6Kf1dX2G8+/oAXDNOyY+qj7pYYpg3rYEXwWCgga5haoTYjs53/JzQ99JgtzVIXFYGaFp15xK2K5
l0Ux/itd1Itru2LMIg7LK2SAwx8ccXeSKC3YWoSq/Qj04AGFj5CtIlzuW3x2I6WV84kk4ah5v7jB
87VYl7G60tbGCjmL4GX0KwBXWNMuEMAW2/2XKifPhCchAPlm2dhOIICZm6jj5vy14053RG00jXbB
FgBT8SEeWXxvcYh5BL6g6FN1eydq0rrEa+OpfFks6RbJxWjlaWs2CPywGnz3PAHHoftXlOSYLNTF
vyejYy/8EBGmRtdGYr1hVgDuEdg8SWAZHk8ca5WaWnWQsmeoS/zcN+XHHwKKB82Ky+8mhhq50FnT
U9BXuZpck1+/TCOGRYSYMpr/FX7WoDBhPJFLXNPn56M1JIOj/V7rvC1vLWiwyBEeY43Z8k4PAc7n
vWdS51rTcTAybJ8Gn0moZMUbtqR6XiErYbbVRfJezk6UhEkFE8FyabR2+bzLiHNNZJxoR6xiphQT
+hX+CJzzmRiDK66ZJjk/NPr+AWMov8m/ZOFyeDm+MqOhFPNQvUhFOki1IRVILWB3I5o6+ZOsf63Y
Jx2q3XZKnVp5Lwbl6+G5v0lRvfNaot6aD44eQMxLyw3U1cTxynIAr2k+za7sz5lh+z74U0btCSSn
p+uJ1fbebCMMYyFlo9sQgwRzJa+UFAvI+OCQIaZdWm6YH4Ua0woLpfVgRKJzUME5oHToOR4xehim
QTs2IgYqsKiepCqq4TKkH7Qx+PPAFxeqXN0qPRpWQfKOyUSekBKPii4PWc1c7pUmx3rgQSnCMeak
IBPkW4xnAo8vwArlRWIDW4buNr/l/sjgFVqkDKisMJ2wKZyskIlsmsSTEuPaBdq/hnKjZ7Khk5KJ
IzXo9Hs53+pj/HUUGDHAJTmSo3Tc2Fol8aYPUAwr9j8p1BiNATpuYxKw8ccl4TkmeZEqhDd4s4U0
ASHs5FbUwzB8kCPGNfB3WZf6eguS8k1OhCMQgOTsV5wKytjaZYDltqk0UU08YTpy7Yuxgdd6W65E
Ej1/oxmjEv1Yx7chfkQ82jl7DSGsgns/x5HxiTd3KEErPPbLKtdv1ka/b9xwj1J6pJB1pBS3Xl2Q
6mmKZpJ/gcZ/viMdXX3P8dA9KFjlHc4YXfGRfoe7IkyNui91tjC7/uvnAmg3O9C+AGJ441pTp4kP
sZQJXOJ2tHxR3EaXZ+y+kHkVDNs3mneELOX5HI44dDpUyjsLJt8JDQDeR0gx2cP0QDllxC2IJMLM
ku9hT2zIQrb4rCmcUd4jkClwCFp3Ry3GOyCbWrV7AoonkfgdmiyslQiROK09eI8WD8TtNI5Cg76W
Dkry4r9+px//cKsW2/ZY9uuKRq2HE7IcewZ85IyATBaZ0alZ7SgkG8q0b7oAipLTgS86NuCPYmzE
oJ6ekS6Uw+DtJaB29eQ7cTm+zZ3/+qXwUpeh0rJDRD+JnGtnnBOcdjgURh4sigeBhgDiOesVCwyH
WeTRbIQkZxnrDkrgh06HNTpc/6fxOqT6kgMcdt18/YwmRipYZ+vEPlaI3uAd1k/9LKG7E7MSGzlx
Ks0fJjq6JW7s/qaUFxsqCzvIkvaKqwT73PvegbSjiRxWgPIl3nY1tf8KNspQcwlsP+8sT9Uvrm54
YuxhMaJz+H1xiZZxMJz0kK9YvnbIwRPTQP48ckIqqfsOh91R+31J1CCTTzhk3/adQqaNN02TLAUO
8y4HaVRUy7kqDPSNy8nlOHPvrO9qHkWtLh/EOr6BDwLFYctlGe9MfaTzEcKwkPiCj6H3ex8q4/1A
JC8WHA3Jdyn7N9FaBG+xT8az1D4hNSYLuz/ZV+sLAYeG8AnJvZgvboRt2kwAFj/YHZkG1pwhDSfH
ncuGnqsvCyAdniGXkAxyGZGOPyRHvOAn0BtLhTEN1E4C8/xQqvVA1/n6Pi+RJ3VRQiTmPCPx3Srd
rhkEL6VmHXb2PJd2R8fdubHIlQQZS+NP4M3T5nyE7WK9RcoTrbA+ToT/Vix3SYgJ7FQYOkJZUfrK
sPtGHX5SFuar8po/VaJ7USfrqlgIEoMQbXrS/olRK8wsYkXcoM5lt4AOHcsYhNLhRHq+qgqcV1rB
tiLmhUGs/3agrUlJU0XlJwYVXo8eUY7KElkXEyCkrU/sND83qsWtHKHnc0H4gkIL0YNH09biwdU5
oRvNrRTxXeJuIHr5ufCUQd2LvhzQgPkM00xVtXiBbtnRbE1ESqzBHXdDAptCTwqXuiU/A5rrfcap
pfmneMWdklvOWnzCNK8lGUeA5YnETxJvaPR1gGQvH8B1drL3qYwr6C/j/05mtAyVCAtRGvsXqSD2
SL273Rc37VDbT1FQUE90V4dtmgMLNDPs35cpE4o3e5TpuVjQNpCKqtK/HcnwXhlPoE1CY6Pgc0rX
5ixD2yabk87Q+afyENNSkmnDAvIQakAIrh7V8t5jeHyMMw0BEar/uWkFtSzzhFzx2K68NuANXiMr
vV4aRr+vMO+zfeNRCBrGUzrr5Zwx2/y5f1SIjvNNE8nsF8wJpidg5d2t/oWatEsyY2YbrBe1rHes
Eqcf1uTrgn3s4XirJDAEcch07PViUTXdVzYPB0c4CiVYuou2JwdtXyJngoIsWe5r8vxJvXIcteJ9
oE4blwrEImRC2sueQNYUcRRZ1RSAtWapJl/SyRVawJfxvIH4Rf4Nr269ZI331syxX6y4xqJqvSXh
Fl8wHVn36Atd/3NYwIfBxYeIiGAqBU7EqkWcag27lZBFlSM2gWU+u7cd7+Muz6qdNLy4wHWVG/WN
v2JSzmJ9U66S48KUoJuxJnKiFpyTePyjbJ09lyzNh6OwdedB/Fd62WaM16djPqwIW8QyQ/5INznK
MUEyklJNV9oOFIIXwlUHwcTSHE0K+i2/NOnZjEaUY/tNawTSbA1Q++noPSnlMxKs38DlnBwCcrLy
Mo1I+SBFJkp+N7QOkqQctyU0HWuij4YmXagbKEIWnV5mB1LjpUHPUEVTyTE5SJUb+WH0l9eKOe5e
Zn58FXvaD/whqDr/OgQRZtd7Q6k3PKfjwSQulWbUmuiOYX4MF0LF5hX8QutSa7e0dORfiOqtpWww
4c3NeAQlT6GvRje9nODF31isfZKs+9Qc6qViubbErn1H3xk8orNhYj15FhJliWtiuAj7uzGSbxri
a/4H9uXszhDlVIjCyopT/olJe1y1czLXJEYNH8aQF1TF+Udtt6UlfKH3o2A4Dp0zFlR6sUs77XB/
zKbCpOBxowtzlzzlY6G3TG2q+gghPPMcfqQdKTy4PGPeOZV7cGKGPYfE5hEfsNjXcafYZ0mSxXqk
gThgxNqRICIMvEgSCL8pvEXVODBb+3ozvqwMJe3D8Q6BK0a6uf40/7e5It8xcqvWoOzmviHNwjI1
3leriLOcRuFhnr4keYJkeH6x656y5QNiZ+HAJhStuCfxzeadfi4nCuaxsgCSmucQk0BmBGgpopMr
nq6LwrQAr1gH90Xhbj/axFq2KfJIurr6hK3ngkiOZg5OMjTl2+ZiWME13IbKsA2MFb+eNe+jyr0z
HJF9H3RqjOL9pAK+QFTOMxjvYRQtm6tAXLLiRgkABbepIZcx3yBlaUYcZqszK6QyBSu4B3ZgxAQC
S9cdT4ekSwL47fPqvGlfYcyUWHQzAh1wGhsdAOTnK4og+7G03uzjeSwtW6Hbx9lcCKchIYUqWSkB
Eyv+RNSJJEWtqjnigJ3DDcrW2UGGoDgZKBimyXGA+GO3PqYdRv6vd93HBhm85C268tk3Tjvamev4
VKY0ncXvbZP9+uTyClAPPCtrnES4psjcXBSr/B9Msa0ndQ/PhpiHco4JRFhLOWn5sbrgoX0zdTZ7
8tL8eHqR9czkKhQEYunAgO8Gx3aiU5orxd9wyrToNH0gav59/OdT3GRChKEvKKNuqzngfaFWH8NX
u2zaCsstAUYMUXRmOsdnHlFxNQ8cjw1h8/s60EZ1fXJlTDGda3TP4OyUshpbj7np0RwvLysYbWLn
/TAF9glALwa0cIjpeQgXk2wRgp3FnajYtgKATuVoTdNqgsqDjfwD679w4aVc1Jk6SKHlzwmip3hg
SWflBK53lDuQ7umIx2Pi89QE0CyDGLoeTRxKtfv+wVZU1TE+1Dv5Rm+Sh6y23ZdDoC78B2zFe0Qp
pXwWx2Ki9HVkh7PUALH+/mC48cQZ2BmaFgzTVe89rq2Qm3qNYb4p2LTFYCMpVsN7D1CTlWnOxsPi
WtxoIsLf9q/mC+e0x1hQxOnfimYasNdtYlB6VZiv/OSIqC0EXFTFw6ePx+W0sHQO8FHiMftDky8A
JDy933qysHa1uz0y0/BWd0B8WtwST+/b2u+dfQLYcGKePcVNx4zJsalwaCfNOLHnJLdxCW60kA0T
mEty2wx6ldhZq2EmLSQ43DTnx3lecfihSORc1FqXF5rOWkBtfY+cNbfC3q3dBjJhl69qQi433bH/
1b3KWHe4dmbidonY06flp8UuveMVDhxjQgksYgfuGpf7IOXrpQyay8jz3Qcu6j/wmNOtdSyUq2Ho
n2fAaU/hYgFSYinzemTPoGx4g5guFsZCfMnk5CAA0dQDaudIkatsNTufWjpCmMBOK6WKvkGm9eK7
AOo1/ttXbXvmsDlEJx5k2znbV+rQ3dRkuyUST5POTvdkeV0LB785ch0k3p/uYAkQijvwJyYDXhQe
B1sZqxItCGmad5Jlufw5OgpkbgA063sUlW5MzlxKykzoHjMZcQBFZrNLrE62rfymN/zZOr1AAFfB
9XG74nXmkW3S41D7kCiaZRCKKvRFVpxxupaKpRnqv0NIC9s1BPIRdPZNRTzj2Y8cjSD/I5wf8Aci
sSWRRGhdQf/rSQIoyC2zOPv7tpnHVtrfwsDSU5VHVPD2kIncQO5cVPEtKBNfSNUe4SJHGB1MUKno
b6RdSdgdU/6EHuWXgkl+kEODPgUasdevbP1fcON/BtiyL/OCSJ3BqqA2JmbkbXPo0Fp3uTEO1wAe
KfzCGvKKNU/yoKV5cHI0ce4/b4W5ILxnVQDxwn1GO1XkKm0mwvOngDjsB+PtsZeacSEmqAMPNDcA
xDV590hQCIGee29P6GEzzn22w+c2hhERaazOo56ZkD//oX0o+N9O0k7kwlVgIpWfCY+C+yItVX8o
nNa/Nr/qv4pvQst9oByo7/iPeInYJ5dxQ5UdnSoY/R0p9oSFiNZ3Hrxuws3VreSJ6NSc4yKKPaHx
G8fZ3NZ9f7Iv91YulgkSZ6xkFI0ITAPYko4vxu2A+uJ/KU6C3PLRI5BkdRGnkdCKTH5amuKZL98Q
fbWFcL35kC1yxwSzlmQhQp6Kum07yk1sV6F/DgaTjqDlSswV0EUOY9U4w4E4E6ft2PrsiDKdaTmB
Og0B27TCMgkEa/y18Q8nviGQHvYE9dsESY0fTzACSnXiV5epzMNntrXvGxmncPd05KqNB7nIy9AG
9gUJd5bcIGOe5pnVCW2/o/qnyPUcQWTd0f5gOpxbbly9oKu5A+1x6nNWWoVjtvU1rG6wEeSVkQlW
8KA+6XEJsnUMBIfL2NuMG4qCEnaKSBDM0nx+IaeiwH4nOyUXg6ARYmN+eVHyc18nC5dCtd+4sGcc
eJebnD+kyHbpyjToDsrpyePJEm8+EkYJB2or2j2124bTbIOdYSuNqt0Ire0kn0Zb4lTA6EHT4kiG
73h5VJbteuF4dKqrfxovbjA/UFT2apQbNelK/9lBqyNKTm6Yetoil0JnenFTo9scecw7XCziWTpP
CyT3sDyGgVhUTtHgi2on+NXMSO7Amkv8bT8yCvNwLlfNpnWp92ffQwqxwOW2uoWKgp9isnGR3n+5
WOcE7PVeFGhWxSNt6xMxfQhIbuog0Qr4zGO2FH6WS30TMvpkTkwn/6duAoCV19CPqVxavKgcAWxf
8a/kjk4ZqZbHEv+8daPvfHjVaGvZiTWG5XCseDwpSv6zyf/wIWyrBI2jRwif2ck+ufi1tAAmQiaA
Zd9xubj9V9f3y5L64SuZ+7I4bzYN4bYxDuhB6xOj7YP14UBntgyBkBBvH8115t9myiFrjfO+/yqp
UAq5BazAkLvGMtVFdXPCHWMiy0Ie0A8GWGMZ9bgN8LUZcCrLa1T6iZwrlYPuI/0sNwb8aLeIzbf5
/NCNWjstDWjeri+y8VqAqcBWOKNvGe9QgZYQA/av10xVfoQOqVJ60GaqfY8oYOyDOuZOOTB8If5F
PsQDTrwyjoGuFYkLF6BtHNQdyo3t3AooEQYbIesqwLBMPzWVupANZh1m4wDAMnwuK6Egj2lDn41c
Eu8gZfz7faSCkp8UcXTwDpzV6ObMG71YR2Yw9ZtQLw6qXj5ISZuYxv+iVze/fOzVJIrnwIMZIiP+
JZWHUQIMLzjqHWdEpcKWi6B2QvU8L2+/JPzZXtDBChvW1midJMw4LKRPT+cBVR9dEbwECT0JEriw
OR8syN6psiAvTVRE+ZgGQEnddKbEIEUYdUUjLPfTqDdZCBLwZmnRG6rE0gMRT2gxn6GKl/sj05nN
4wa3OcIPW9bj/xZFqjV/mhY7/PT7v3665TM9E7zduESgCXoWrKSTvu9d9MipJBVT0fGbKjAOs2FK
zKh7pSf/fLpDIJ/qJD+2M6QCVOKS1Qd7XfjTuTXivP4R+odXmwHWsHDSXOmo6FSPVxtSVNxFXvye
bBbqsyfvLcPMkI4R2TsPzKERInTeH03JbLItHsrnCRvq4vWO/Sa6qF+8g5pnSxStu1BjG1nNeEy9
A+1BWYhBOiTuKN637M4Hf/CubGry9glF3RF4pxxOBbTDa1VG9MSPmgi23JD92Vvj8nH2RXcNEXcQ
hqWSfXxPqVSH2Tu8M7hd66ubqmFdXpusi7woqkqRlPaO6qN4evG3/8l3Snw9W0DOSGWinpYvnr4g
o/2xMDoeFAFVBQEK11koD+iFbk0OYfkDIYBu4H8C5zAZBEZijojEaU2hK9OOFUP3RCrij0+9YNKI
rfFGA7iQgTJOc3LA78hjo4TZXDbVuyTk6zRBDDyINNKktT/p5hUrEUP7ZGlW+kJYzlCq3LPlb2AL
7FmCWpha2BFcqi1CHSeyQJTZbqTu+EZnIMgbEtEuXQBbCwK1qUvE0mMrpptvDzoJeTn+9c2TZTG+
P9b50fwpCkDvzIVnzBZ9WHbLvitWfqIS4MKSiBEZHZCqP81jR34ibkGdvymlHGSVD62KpVfbW9y3
402ofx4gJb8Vo7FmWwq0Ivap9J4b5sDmnJFDTQpHJl16gtRab0R/mvTPdLKOJzQJnuddiPI00kf2
AJy67WXCiThMtZiu0fN98drfs+cFN4hJ/U8ZO/FRPBwCw9HuVYAmtbNVwAPR5bj75SVbpj/iJGhS
B6NYkBra5gca2NaNoZcApryKWm/OSlOLiBX7d/K5TPv9dlZ+5WTHb9S3BLy3YH9TvaI/GZb/Js62
6a+EDqn0dCbSlXL8vHQLaUoPb1+C1qJw8DyK9SKutklOtZq4YKjw1TosBwEzjQTuhZsvKklBvotF
Y+6EZmgPoUMnGKHhY3UNVOBcnU59gbxdaOKCYo3IafRLM+CCHEWVJBDSOTQNnUCJbpm9jqc1coFl
K2XL2zEs0thrqaU0P4hWpqRKtgGiNMH7X/C+utk7oPthTQ+9qX3irknA0h7N0199Mq7NeYMlT34v
gbjWvO9izLv3NTnByGQ584A6easoFAFC3lSFCZYI+7AQCzgg2XLAb+ltab0JAipEj0tkrYnfrnX/
+evi4s+Ppoo+4+P4JlEwUhThdW8JuVhAtPq9MJN11j4ay3jS/lWLmc9AR3CvdNVucjf/JvSsOF3+
4/mf72rfU4nVVfyWWSW202C6r9gqOr6MpGoOVpzKZrrPnNgfu+I3G219BtnRbsbud0zKPumkOP+o
g1SA2BuvXRIQ9jpm9F89wM98OJ5UwYjidAuZkKUw2Dv55ugUUumOblS2uZucalOf9LgXBeqgsuV7
j5dKUhTzcmXWD81eK6EgmS2fxsPwU6Y94OLSYwG8LipLzJbO9pyfh7t0rEgeQZbOlHYkZYciwHw5
4CNQbsBhqHiVegaoqylNo9W2IqcNazqt2ZyUfXUgvmybLKLZgbgW40s1tp7L5r8Aer2xkkKoVp+q
QpweT/jZwCJkbJe0Oac7aGcJKKkCrooBDli218X/J3Dhd0DDb3JHZ/MyLbiDpf6we8DeaY8Xi7c+
RQTgpSjyCpCs+06NCHtpp3eUty3LCqi+PEElZTAAP/hFARZYQETAzkcn1kTTERWRLFOeoAdKJHvo
uh+rXHCknKzf4wD+NUI4m/9l9dAwwG7G4bWw0RtnAt5FGp8K3t+TJbYxUdMkmYlWqBuZOan5+uZQ
fteqwLff8M+jVib28Jl1sPrMDAeqlKUAHSGTv3ZSu7K4NNuNA74WNWXdzeON8dPdHo5/Q+B/3HUY
HETHPq1byGJAq62L5YA/CTCmZgeeaHe/y5TqbOozviMJn1OqTYt16KXaoS5lkK9sw7GilWT9K5mc
9AAieoI2oGh6GimilhabOQ/Jn+LoFgK0L3t3p5B9Yql4cnhOQouY861ucieqv2Pa3gxUiXwM4YHq
//koH+Rmsfai3FW7+7eAuQQcJTb0w8/cDIPnk31bKDuhKGkwnHo4TRX29zZ0sa9SHX7M71MERm03
2c5SCQjsh9hVk6HsaNYnM2dA6vRKUMc47vWWXoQvtskSDiLvmScQtwM11vRr5rNt7zN/8RU5xM5G
i6iLxM9snmwXXl8/ksUdGeSN0/vSGPqRMqe4RhWCOBH0YvqW/YGHjublXr2l5AUs7cxxHbQmr8ZK
LIWoOzfKO688GiDWJ3AjeCe1mvuwDG3VssNDZHR2I3dXZzoyT72Zf8vYXQlxWiPmNAzq1c6Gr4yg
Y6KlSqiZtnPbk2++zw3kUqYKdhZe3QYZ8I6yVyqiy7SiWAwSOvbyIXEVXHGewn/0JYTaslSRbHyN
tA6h4Gg9LGFbdv7Ka1dAjn7tLFkJf3ifWJi2KiYYNNQM6n59LOLIaRsc6DgrYXEQrsZ5NbXpTqt/
Ho/DVpcuzOMKe2ygtKeQxdjapVx4sr7H4XmO8bmSCJX7XcE3tbRGCsEj9/In5D6qy/GrTJEqh2eb
MvnqC0pHi2g5l9aSzHTI5hEI0OhpTwhQnnKy7S97lBwfAOQhF+0vFKPa9rO/9ErmkMAVwZrR1ZGq
WsGpbnpzAT/Q/9giWHamwOGephTw2dTCRW5QsQDX0LUtMqFJMbKhdhaR8WeN1RiLncvxZMTLmpBT
4d2aZEkOjP0csJAuD4PjZzay9SdW6sdeaqF7ZCG/q6JsmpGscHanItituOzWqDVoOHQ25U6GAfRf
hVa+ZBMIdEvhqp1WmlT0AEU5vbecyayaw4ig5tD/BLiBP4HoS/CgV502IcySp9kPzkbCqR16sn1M
dvbKHwM4FsiMB7ywRiR8Q8TOMqD5hIdNohh7yJuEm9ick6XlIZm2m+iB0ArSBjtxnwrxTihj62qc
ndlyolyphSea77uwZeDBV1/w2rkbwo/8p/14ECtZeIMIrZMIOJhk8WC4VOTTNF19Brl67ZKW8+S9
mfjfUibcESb+6PxMmxM79k1T37mxJPcO1aION28jPVeEbYjqyKnd9Pg20o6jJIITdUUrlrNbgGxU
lpXw/kHKIUn6eC3th3ZaL6nhE+JtEMbXWhUU/0WpwzQLlpVSjEpH1oh+DJqji1bzncBvOTHH7fO6
FDZNxaDgYrtLxZ/+5WyEwEN/88606iRewNYeffpwY1jIIeFxiHkQiowlaKVjWbeRGq3c2cBX2qH1
Co34CC8Gt02v8Q5zQPnvv/ZPJXA++Azzm7o2NnJpoGy8gARKbyAJ2YM/IAYv5Ftw4UsP7ivGpely
KxuP+PRgUIHoOjE3OndWdjE0VRuyK5OW5qkp8TxF+Q967ww8ytt6kIJte1CDk+mL3FVO2Msm/glu
C0dbQT7PE5KdvrNd/V29ikD7+P1T7L1VoojQZFNPLclGWOLK/X9l+8PR8f/mnVt9KciwiwrEHDip
H+xye9OQJ3CnFPbeBgCePY9Y7+lX0pzLtkL9iD3We2U/5wcPCqee9/vJtTFw8Vx55zuaxNFp454J
BC06epmKhM13ICCsnBJoMeaj9VuNMs3elbKLdKRWCesXdrXmtI7ig78srKVw/TcSsLKc/HWeKAfQ
sqj920ujLItT4F9dPN+4043t5biNIT9jbh38JbG67DfyuxnuOjWiALeRGBAQVkALq8Whj6hfUdTA
mXaesJITMKvHbhkJ1pWBCzjaNm1mVYkEjDc74W56qD2KtB1V9qspY3J/sozTpigR84qXdN0LqIHo
qbEMj6gedQ1hFOsImY/CLrMmrY1R7vEZsQ8IQUaPDXVXB2c4pCAs3DL55WlgcPFvNAPOf9GQBrmy
mnsS1m6T7DCpZPx5rRbcJPH5H5ppAfMvOJrJCHaRa2vs3B/AMIcLykjxHTNKaWJJp3PnmGVh9Ab0
LqO4kFTbbEZYaJpwLbcLpzuJnPXszVM7gYnMkdLRjr96mVz6eTnE5WgaLzu7kCZy08DgEqfssIyI
bacmxURZo4T7tXLrJgsGw2ZRfCgFVoF9k6BQUEDH9YJM0LxL7ZTNAc9FO4uYkud3yc985poe11y6
oKOHXibA95Zr9FgisZNmyPD2gTigcf1tISLK+HfManhITegu7AGOsud36qPyfE+aVxeaQTcMIf9Z
jDNxdXjBVW7fX6FJB9c7qm/4tJqbHODn1mEhoJ6zvSpTafM7lOhmPkkYRet/03vArI/ZHVxRNeQl
MBaHTgQ6vrjH8gvnZU3IkIZfpHoHIgj2NOPABVTSkWYMoNhAweeXIzwNHiK7lZpsvi02qnzZlNDx
HFkjWTP4WtL68aQHodjByNKw16RjuioNlt/hRh3QCqzyAB6yaao8JDqqcaD+8GNEavOuNp64sjv/
MvQ/7ow24SgvwDQfuU82lxmZYUtKgwoXBYJXdGZ55H2nECHZKeDJN4e6HIaFMGFwPDU5TrWRi2jM
jCLhdjIpQIM/nHcKiXsg7G2ey1h0pvaHiy3QPSCoD8N1XHcG+ngIll8083Ju+J4Iq2Sj85gvfc1m
BT5/S3zdMCB7qzi3Z6PN/TLj0MHFOPV5tKo9z0Mh/Z2t37d/TdQTw742B+IkzTqXlU6Y5z2yZTi9
s0rmmj+cQ1xOCJz4JlhhK4uAHMKAquJOTDE7DO84IC0pUSrknClEpGOmLQdwSjQFlx7WzjlzLB41
aPQ6RKSafqBkSbjX1/k6q2fTXpAssrXBXPHlgXbylp0DcH3tpLzoIKiy5L6WwO0op2HlUN1R7X6v
vOtESlGMFaa3N8Cj1E2Fz50hlbFJLY/hCNuS4TmHaRZ2cIc01gFTK0d5HDJkMZHRky1CyE+XSB7G
CPP64ErBhQlRtnXecab2gNSu2bOYbXguLAm5WT3avClrpWRVpSTK2Sp2+8yEjobUUzFb6eKrl+Pw
01IeeX2DzlKYvvd86g2mT8m3GSiJ8ScwZitKoz7GlZQEPKxT8F9Prd6rIMYZSbyqkNSBFYhM8ZUK
GJN7vWjVAn8gvdA2hJTcOBJ0hrapmrriUEBATSD7AuJIHLSv8kR5RXH1wnUh8VXIxvHAMZq+sT1A
i6jcJFAAKrT/rEE3P/fi6KGZ3EFhCCaNWscFUIKLA4z/WEh168kHglwU6nasJvtFra9elq+dtdKN
aiG+KORHAPJetMl/1er39tUPSnrlfQ4HY54NGCj3Wd0ESALTpb6BB9zZza2pcgi1Xfe9oLwroR2Y
BPXd4GT905MkWcPOAzevahHpokIiQ5pAvC13Xhhw+fRAvt2PB7Gc7P7MlY4jSQfL7Fvqj5s26dqH
38KiqUKhOscnzOoaGIAfuZ5HJhgb9h1PGSWJzosJx0cJogLDLhjB0fMiNO5n5cKlP76LX5CI/iFt
9GAm4a3cYY6T0DQK1BibHm42apHkNt3iPGZePKjcDo0bD0tWVGnJ63yRfUwglniOzPaCbg19RqjZ
sPz9PV/vHELsNa1CNyVHwXCgguwFyO5UtJt8D9i24ehYRn2QRTiEzZgUDePe+y9uUVPU1lrYiNhI
bCgUPu5OfrvrZ2ma+TFendHGE83EfwK6o/2tMP43jBguaVhQqWTSur7wDwGsPwG1oRqOS0PssbVl
StFvDpDbBodzuEdcBLvBJBlccB5+eDFVIfXDLjXkBWCXEdJO+BlbXwU7YKgPP9cR1mVC/il09RaF
A1pDasuq5TqsH1RTSNa5ZHu6tOnxLw07V0JoOh/5ZRgaCT7VT9TKzDE/8sYmdALtNHmPts1Pt4A6
8owgTmbTRM3LaOrQ/USLOcFnmRc8jstoy3xAQQzdnv1NzYkZbjVwmaQnMtD9DiXnPr2+BuSYfS/C
QmplYzi4Vp0ab3Zn18dOwTx7A2QrxfMPPRe6RK//5FOn64QXS81CX5v/bt/i6Stkhi335u46gCRh
7IZuCcYbLlpFLeBhuCqrKt6O3aXPA0KR+ZkaqxSxLuo5oRkV021ThTDPUIXlW0t3l1AjQKvJQA5U
JJ4jMuJn+1PmF5d5ULDlm3Xvz7dH3hnZniTkYtTPAfoTYSFIWU5aGn0EV0cSFob8OtvY+yOX3p2j
GINiQ7KYyGkcCYuaexNTDGtXJjI7qTp24jPDw4i9siamLsA8nSvc9n9k0V0Yh6ivS0pb9TAXFjbW
Qs+TefFatus8cSV/EYkLgR0gGLQPPpS4XiKsmwUpb9cxytadl99KW5kV7HvnWQHb76bLepwT+Ixb
uGy8uVpZupsn4wibOcyvT9UOhJTCSugIpkCNG7R/FpphdjtQnUesrTXTRLq5VRDCObOuhqjOu7Ld
cdBPF9vvkGB2VTZyWa3OIX9jpu0eAa9nw8TcHV+04/4GiG1UzfQxvHoWnsQFHp1StZeAKGWRL3aG
niJxLeslbIukQba7sP4C3YxFIkwDsAvJ+qCr8aC9Snf9K48cr6YahuXciCPRivWAPbVSa1FOGRsU
pX77EDq3Y80LIQPcCBYcQmUbgBdpDaBrT18EVoKivgBz4Q9mgAEoZOG/wsnzXSrukDtZYzW7cLAT
Ofvn5Bjh5SczCISeG8Whkt7ixVYB9nm4O8AT/XwYnN1QUUfSnmXQrZLSNBfvGjVU60spsyPYeeVD
/GgCH5wW3sZEFEaXLWqV0gLMmqYqUP/drlIjwHq8Auj4OFkaqSgZYW3HKCMtUkFbdWXuUUQuW/e9
vPfTMzT0hgK/SCxQK4BFuhv4gDcq3JFV9AY1T0LXL9UYv86jvqsV3b2+t+m2i3voB7ceghsZCEfh
1d5Hl3O/xZ+qe/Ux6v+StrdOS44QxfGCtlBzf7Mm4ccwe6f7yKAktxMXDo+F+U2LynUmcx3EfQ0t
MQWL70/l7yRaJLtATTGWadv75oJHqVkVB6W3QGFIl038zWG58848wPiPjkfBlRmb+1e259wCJWcM
AnsH0l8N6GiWWxIhTaiGgb7xYHFCUDEZYju8pKV/1U+CDfiKt85tHLZF0jXo1KeKclkIv2adqs0M
QkFu0jL2nL+v47aRsPI+DTbyYkwneEGr92/pJU653IxB55592Bm6ZJLNrvx7D4MSrQwW2D9t3KHA
X6aklh91bd2BTYRQ9TZVUi4dxLw9wnE7xTwySfM5ZmC30DzJdvr7Bmy40oidSNylb7o6gJe/CNOg
O8NXRqDtyDOQzgCWOzJjfKMmDk/Gw3CjUcyVi4XJRIeRELhCDULnICvRCIG9Akb07C5T0jcmiLau
esDzVo169W3dYZ/qFGkQDwPAhahET6JOXRnL/+aC6jpilMf+K8uxfnb/0wmriWFkP12vAcBqpdX9
mkppkVgvnOzvisPPbHzasvHzDwfGa3WA5kPQGLFAcrFrdLUz2bndKNXQwuSlfGzD6yICoS8pNjHK
0OCj3JWbe4HYuSklGXxMYFnpfNUfjHOPEIdqBenkNaCJ82O/kQVHjYQJ7GN7jX4UolsgPjVL9VWc
ccO9s6pz8XsOYP/mgtnM/qMTqaKcD1UBSuoJmh/UHp1gZpwUEE/7kk1FVaA0zdwXQLTEyOxvjRY4
9guFDsC4Ccj22Nr+HeuDgUlO/J3sTbxBf/wMCbl8TXSL72ui0cE5UypPTeferd4EPGf9j7E74i3a
iyCYqf5+svald+wOsBkHDhCuVTa6R3WlLk1JYWwUimf9Z6vTGTzw+AGkK7+1prfzPWA5pgafaTVZ
c7/GNrn0AleOKY5IE5h1K2XiMr+zxrvskWDULzLAPGUjfMcB+UWnxNuV+prKzccNSTgI/7nlr3RQ
LJf6h5DQDLHx5YkgusHl1c2YsozZHshLgtuXY+B/XjwFylroz6CVMmgnBly1mddo8RY2Bv886hvv
6nGZ4ihaEIdWwZbDcxzKVV3xIPNYEbIXmUDHhNoNhDYDfd/IyIWEejsdunIX4Y6Qv1DNAH/LTsh9
P0NBAHbyrd8DI1suoUVKGsjc5j6bAGD53/1rbHYO8trnnJDS3+CuVGchY97Ke/ZbOfxOYJSKEjhV
WV8hDgiGScUI9cU3wtbp78YUqvWDUeiZcJJiY3uAkArWuY5C8PZSFO/jHZEe5isWSsLmEaJk9f/P
6odwEt8/B6FyOFYvxL7gI27hHQkStt6lN9SSeFIkbICCBXZkYWLLa0cvcx1+nb18FSACVdpwiFEz
iu/ZdjJbOqKbN1W10LiPW1NNuUKSMp1Jk+U4rvNvG0kEVCnKQ44Joi9fgFwQJ2upQexxrisLeJ9Z
/CXfWKj1FIt2VBVfoQQsHEzMCHy2cWPH3nzOHplEX5BF/05ebuUg+IlAfZ58vMGVvVAxQMjKPwng
HXteaMqO+du9m0+6QroOJ1p1Lol3evCJTLpWEdPhXf1nY32xVsWvT+rfhye4uvESE/VcSNsswVCg
kWSiaL5D6zM2zmfl7KLa/IT4ssbxVZyU8+d5BQMV3S5UwjK/KjWmac/jKitCX7QJn22/Wcjl89jc
r0PmREYzFPnrybjNOCiNWJIV5Y+KkzWSJy7D9x0ts0aphApHdC7bI4Zlz5Dq3tbzp31JZcfwzwAB
GWLalJXQQwhic58NrIeqMK5MNdaEpAeeOtV8X4oVaX3KXnWvy661nKHWjuAkum+R2o/a89C1QXqv
szK3vj2zfOixuq2CbS6YOLipEcYaSenkUsc4HfKdBLH0Zbs0eM8NlcTYIz4M4YoAxoizhNcAVhTU
WLAvz+rZ4puUsA2hogFgoE4RbSVK+U6hpn8J7xVnx5Em4VTfwKCE4g4gOnHwdfNg3NfQv9F/v2gq
Ld/dGmanvilPdJrLGtgBOTVKxTHGjscRrvmzFscMFqlak5ChJ1HMEpzn8zZdNB9FsYgv8N/w89li
2g8WCCc85PTRdr8NvfTe2zN5kWiZDPJATzmwtivmb74sB5+kbstxGBJoWebhGXkThqWxnDsWDDks
E1hxnlUQ/1/i44H8rirr13LOwOvZnrkK+kM9IkQSeRsLB7qyYdY32OWUy3cDzY6mFtd8GYcrphV6
Nc9WSKscAcl7UV+AAitaCUg2ehurvS1Z/MDOWca3Dw1vIagfikBJn9+nvQYGGnk2z4HzmRHUv+2m
og5pZQDxkTI5Z3NaVe2sKfzh31b88P6a6vYYPbWfAK3xsYIHpodwD9zBNJYMAKIBMwTQcwR/reO1
Ppt/LIDzwX+XgUSXlrnuaFKW8WK4vK8UXaa9gsosJUHkVZ+atom5s2CWbGJY7HEkkD92usOkQHlv
FV7atRGI8PvxfsHt8uh8FPrpfGXH+3Ox0ODqkAh1S9F0MqgqrtxJELf/q295wIesj25fkEt9pyYx
MlHeO9TM4C+zZCRCRFdUD7GeXtaIrxlKjSbTMK9q1unaEPSRz3xbvlzQEfKCQSQRSGQmisWwgGoF
wWpyFtSf6acuMcDEEPrrgVOiDDxehfXq2RtF93dr4qXj0Ug7C1gD/D7CAfN/GKANvOahWdXjY5J0
F3crz6uTqev44Lm1yRMfJ94XhMvK5lv3te7+FckpdZxA94KIOlHZNoGFTrSp/cmWXD/v68e9Et5u
X2bYftQRPRJe5bNsp5NYZyGshm9Pj/jjeY73x31HAGu4o8ebUubE9aGP3te/j4tIloDYnx95Q8Bc
G3wkhA9Y6hUoGOU/9BZeI1h+UYMYP4BfLIHTyLR5huFmZugvtvU57U6+KO6+aGUNO2DL0PrpO/n2
wuHiFPbC30ov/mM+xXQDmTWYInNX4zdFL7FNMgsBRO9a0l+7Cm1YCwBYVvSVZDlTuSBOwZ+WBE26
is72l8f0NEPeuWQWtjYeoFOsGLJicfoGRPOzoTRwXKK/FQ+SgBlEtE6qg1RnfqksLmoKw9oueyrq
qGSADRmn2HdTzLtkFcGKJlbyMcxZPDQGWj0qck5XszJSCytWTXU9U4JoOZcUfEK20Zt88HucV0Uz
t5Lsio9kBP5lKsNxMOxvf0s/kGpIq4Xn+Dx3SDuPfLOCIPKuGFrGuXC8WcibUpq3aJoPPKb/HKzq
wFVNgxDwgTQzgYdPYy9EAF7ZswQ4L6AGwMInN9DbJjwCG2Z7bGndnDiPpGsIduCJ6PKHi31oJ2dF
G2bhv1nHNwbVD/TEPBWxaLolG4QGxjWek3WoiYuxGVH8CLkDS6IbLwG9+CWUdVs8JuIK76AG1cZe
S5XS/ESCoWLqYRW1nGl2ljdqhQNidNh5ATQHLEtMfBvz6NMZZJDTd5fvpPtymeF/+ciLPGZ5rARK
6Jx/jbh/5QfTTezfCRtYFviLArmvOmoNdxl3Hrf5NzABki2q9tZo4sC4gsS6aEfRqA0m4FAUO08Z
wY4/Pq7Fg3bclD07WfRxPdzLIwKndA7ZMYUV4/vcM2+f1GGU936JiZsFwOlVlmgZONi7R0StLEt8
yRh2yVdyF2JVg3sW5rmRtZjvXFiZ2JSUAYinxR+sCx5ZrCDB496yz1GVa9ELSo1CGH9vdH4EPCCw
On9ECKWxqa9VGLM5Dn54DwNEA4g/FWpg3+ip/rga7aXvIC9zM/UWJSTtCsx6YbS7gwr6gb+i/l66
SyBAntyTo1LdTq565co+eDsxrpdBImzCQ1s7jIUVgdgWVc+T+j6KHU9NemO5uekb8qHTWp05ogAN
HrHREzcqvcmo6KAIMw1HrUQ1QUR1c0ChLPC5t8vAPOKxOIvCasEmm7q4gzSpX5UtIZxjOEdB+CQU
pcNECJFkCoLc2a3flPgMlo4JhNny5dQHUnOOuqyaWR2Xys2IOZ4cZq35iyzITB5T7HTp4+IgMaXn
lCHjVRmpK9fNaHP9I5HK+cnChnd07Z8nO14ZOrdZg0Zkz+zvvsHh/QmyUnXO90PA3Xnb+WHpUhKb
hrAS57DSwN7PitWfNt2dSsGNSHV9J+GEOgTWHG6DYgi7PnxSFyopE4SJgAO+Ee8K3crZuEwU0Skm
NsNETnMGIW4uOi3p/PrLi+hmBYGOrZGGSUsIEW+w5bMQAtjPceE6RVKuNCgfBylHRGrxNWsjkNgL
uPOY/gA+pwYNlc2xDPMGfzdCp/dievJoJRFrtCld44NvULZ+IMsjGYp6cHYfQZCcUyCrZ4irLy32
O9y4N9HJBdGmLMkJkeIR665Ti5j0cL4m60PFJ0CQ/TWsEznUWdOia+1ig0UZa+q7jH+gA9bkJLkh
oPmtxlpRl9f/WVdo6BCLAF+J7miEii7EYYi7du4riq0flMpEHpTjruxMG4LT+HhCr/pEfvWeTpZV
c5VhMQnD2CuJu9r9m7geDBamN/h5OPgfCf/lRvaEsaSwqRHhmt9RpGx/DNJKRNcnx1F3jYHr3Dzr
Ou95SBBzso4cYrYhKXrfolJe5eLMJDtJoSFEeAxW2rlhVsACXaQnjcpBq9UlvztOyWD4NazPIQSi
zZe5fXF+EIMe5L++yBgrATHXLyclV0NvdQlW9rgYY4/QD8UXX7lBcHpcJZr7R0oOnMvLjJ+9aKcs
vrNxx1ZQt2HB26k8tQY6RO1BZP6SoDR8/Yty4A88glCq7Tbn8W4aHkkNTw/K1bSnk+jsWC/fX6P5
OQiwbjRkG7ITA7HwQF1h6GbAWzyWhzg26cIUDzt7W7uxtrvqwoBvmY5NsfZlgzPevuaoRNwP/WyI
4PHGov5Y7teYWt9/B/Lm3Od8YYMftNk/1aNtnkq5pu7DgGziQtxLEZLcjJOS6U5bPCmFnFA0vjJ8
otgB91borqg6QCHzy4LFhnGTRb95qU82Egg9ArT/cBSmWv4XvUtF7bpWlEK/0RJxyKLFyNohSGMN
rLMnW9+BAtg/3g8q43eMIiv8ixinx/NE55Pt5KstbwtXLCkOEc87e9retUwr4+Bfkaay6c0j1XDx
zs2nmmSoQ7ipHRwHPJBCD9xKSwpii3J27rE6TA33VwId36iMkR9LbohbYZ1LeNXyFOWTTI5aWbFE
vKI++6Ol6DVW7xF6Iuuwmo9+DdL4ZNp4KXmHVHft+E2v/GQ1FHdKB2mjVM3jd+3u7gv1rSZZewux
zTk0RzC/8MolFv8KDryxZdBHdXMXcRpaXSDt5+/E74p8pTHqY5J4w3d7LKuwzfT55v+lhYnrgRak
FQT9fWptwiRHmGjcDKz7dUqatqhS4iEH1zmcr21k9JrmvtJ/+EcNrUje01ylTIWD8Lu7j/vzVgvy
/0ymbQAU90LRK0M1zFkrokMb5VjtYeFryW5y/NaMl8iwFSzW7kv6WUWcjH+BKHh4NFPDyW5dKgvk
9XbuADL11TExeOb6KKwOUWB64dNr4d3XFQJtsVpgEM8sSrAhvPaOrepNJBuOPUZki2HC5TkWRjOI
gJCpT/c9Skl/VCMVx2SNjxksgUofozek1E8kQZ9iYWPQTurCnsb5qfe9ttF0gnfKGx/ot9I5x4Pg
IHOvRhsCHfoRcoXb0Ox4cqqCuBgGAy2Odavz0tJ2SGIWyI2w+OH63Idx5BWhbTy0TEK251o0xJ9D
Fk/DM55iq1bdC5XWp1geyhxlr2LaJNLAc/SkDMrY5SdF5/IzqSHbKK5QQDTDD73kZjhgQyezB91c
vJa48O1bT/H4iSlOTamxF+pXvoLwn4BC1zucH4E9FRzX9sS5RjjZiobs0NToVNUhv8DL4BfkrlcY
gBPU/lv0vXgPdlBu5GHXiMJqPkLWJ7qRAx7OUzDsdUcMQY1z/Rm1nU8fJBoUu4rWMoB6ejnAbuZJ
vgZl86VCc7sHaKX05jTwXGe2e4UObVjyeFAFIxwzJ9gRyqJtTFcdNs/dhzdzTRUm34ER6SK+keuE
W5BziLNZoSWuonQ63F11mUG8RGR1Gmaqxno4zjWKPIAgnKK8QSd1plKentInZumgiGYnYCfMEAZd
ouyLZNgMci+TcUEa+1p1V8sBKDZ2GWIhTwhuU4ydnryB3MhRaQGUH1WO1ce5TWITiOFK015Z3tcu
W41IaLYjUGpt3xJ3SJ2rghyPVTCz00JIzINvBvQWD8JLuruUmx/UVE+nJAMRyZG4QezSvW6xfXz3
gnctoG+TS29R0Mw8OhCqIaD07rP1lIn/TyT2T3OEQCQqDGHMtxqwiHQeWFCUqBI2yy6291luz6Lj
0HNoV8LCqEX0JIKzwDMib75ymaT3k31Ki2u9WL0sPveGPr6+IcvkzlcjAxXB7HLTc9wlVlrQ2diU
9X75PYJPV2LVVy29Dn0qiR885hMB/XUa8Y/MgEnTFtDebXHrkMZobWF8dkp0LXZlH0nhEEjqk3hR
8JAWaosZ4KP++lLUgdZUmIrq3i4LwYmplZVOuFTvcoIn8KA+Mw3BcjGUTRrjQaA2wdWbNoZ0/s4Q
4UcZcSbgc9eYOjQUx63Z0umfoanL97FC59rpdsSlyWK75isOD0/b7xYqBJIEt1Izpn/+1/UAWJh3
na6NSl9tpdwDxjOc6cAYYE48lbFGy5oQyUgMMbafimVR2n1SF4GszkfArFVpYYG3n6CT1ak+Surv
9WR2xZVq8cYm9u+q4AfhAC0Tcq4fq0t1iEa3rX+dCk/kEl9+FF6alY6tFAdfUcOsM5CGwk2buHBK
EvXbguBafjSUDG01MgxtwNIBgHcMUt7NLqAWuSQ31LIEcxlK8G4C1uE/n4hAniVDwHNenAaM46yp
3Vm+9GUI+MERDQzBNZQAK+JMnMnumNt+IaZV/aZigXhwnKRlZvSPnjpuzNLfNjDsMs7VLIwsoRfC
NQoO4jxVKd/as3buphgiY4sV/g3bNIVL+9geS6PTprJ2YKyxW6K67XEYpQNdeC03XCjc3rsJT2NQ
+7HkKsisx3YpoRrXj8iRD4x2JEnq1EkIIu8bRJiiPqV0MggR6hoA3Wrc3BA+dADOnVEOULtpQE3X
+hTywYl1X1x6XJzMHaJsrQzXwxZx0SXGka3tqDOzCCgIZJh34mM7IxuhAU1ICGAlKsPtJh7NWtL/
So/eM/G6OMuxm05QEd54zKGftK/nHLNx0v/QV422r6WiBWMZakhMMsetzfSad6moMr8H+4vYCOEf
vsuY28ME500ht8y4zl9H6Ll4DhFBAq7yC69mquCNLBFISlV9HPvu7PR2I7W+oycTO9NxF1Lbu71H
UCSFn2XTFWAMeAhc2fNkOPXZEJfjGrYuEFiRZcFkPUzARLwE3xnjeCJL0lqZUIT0iEQejb5B3VXr
hzHcXmOIJuicic6JSgy9+SiKWAiTazD5qFUAGcoIMtpZc6MAgaDnDShRM4xmvCUyDeTfB6otq7jJ
DaJPzj/FV+X82o6FJBxaSMOGilmnYnjgYAkc2n5fqNvGsqlYzeowGOUGmY6oK895tEQ0jyXezPZR
sd9bbejTEb69bciQp6qiAp8L9rNGjG9uOX/mwWeSbopzwPXHzTjjl4gM2Fi5/HrXBJ8ZUxpSSWNU
T0Kzp79fX67/gb1DynEciMpbl2FeO+raRiFk8m0PkuI5s4Ay8vsDg2GfCs56GaZQkVq7M6co0F85
s7m82V2/sD/MKyKMKwxaHSFpdW7GOUjIdwIEBbhfJ1ibl/T72GKl9bMWyNJxiK41meVqE4BLPFeV
KPJECaKKPhxyk+2IhL+FgIL6SVFVSy1z3rM+dxJih+E7jElLpAm8P7xfcKmb/MN2cJny2zZqKszA
AOvpIv8cDO78uECCUfd6UjdBMScfmUSFp/VpUB81E78MYc/hg9/WqjdLJZSLthZUyB73lC49s3ap
q3QCL60aNi0D44bvlgGLQYFz5zyyU9bEsV67Eq6EIwyA+PoZg6qvpXnOBtZQDnjqB4DnDAs2uHHo
LIDq0lUbO6NT6pp5oIXCB7EbmZ2qaoxVzV6AffzCNskK2WphdDfX0tY+P9m2yvDveiBBKj5Y6Ecu
tcXXwZqYzXVQsCfjgvoLEilkmH36dYNJfQef774bu3rTSbWiNX7dxYCX4Y3UioY+1N4LFelrBGBH
Slsh2MScoqK81+qPUCOqX0VFMFunUTDdK/TbiYLeYlhv5Gfto4rxm5K17+eL7+JzK8l7LJTwBOcX
mevf9jilo6J08X/ANoXZyt6eJqua9IjxmcAG+aAORi/jLRc9+rdV9VfsGlg5KReXrCVoWRMXTuFl
KhWkBQB4TC/qZJuTE/pMsuRNPwQW+UoUw0J+B9ebExd4bqr/mIMPot38aqntgANwsR4Ulre8rkgx
sFKaqdum5LeBUiBwznTX9W60Mxhf5i99cJLE0YXJzgI1pFjneeYcgtd6EgVsV75SmHJA7tH0WMwB
j+bW32ncu6lOAs2OnG0cL1sO6IvUxFdVyXFGi7m0NPvJjxdlTRjhgJCYyPw43WABsIyOHg7Qdqdb
2LUa57lgrXGoy8nkTomPxiDNZ+KXHPg2xzYfUOk8jPBQYPmYle/UOLz1HT0QPR4sftzwWRtaM6so
pqiG2l/6XsjyPhH+lkarFNLyRs3vwIJWjhuXEUZThz8u3OeKh2JHmfBCuAMCK1GJ+KJAeJiTwiqM
mDDveNoJjN2LbPWex1jM4IURpoSyWA5snGSd+zfZE2d2gC7HG8+aXUtyno+jZkmrIkI18TAu8JFd
sGSGfl9Kcnkz1qKstra8IoV3HWUVhAdHolBIWOC+qzVPNWAzCuen6fDfpdG7nG7iF9LU/jes6oRL
ExasE8LwiQDxV9xqmQrs5Q3jbD4I2b4evBW+GH7HKSAkiL52S1MdFRl0yG1U3fvIYiBKwbNKk/NF
RV8QoWGUwhf3c99p9Or6kv/h+9F3QW+qmGYu5JFLj6iWk7/QT2ex4lU/Nr7NPsgaNh8teaQEZKOk
VeGijDGRaN3xh9CJoBZ2POp76Exc7Jy0olID9ZGLP5zw1PH4om1W/12iPhc3xdohAxreHq8tut6D
XTyem0Wu0V9fTRFsyii8FPxbLBonNWBDHbBlGQLyAtw+yV+Pz7WUeW3MawNg0ItoBy24OeKle7vs
eBOTpLCL/GfHcLWRXIk3+JfD5aMXoFISmnyqtx+PJeLCnx8X+DnHk36ZpeLBKpjWXjbsn+DI8LNV
AISHZbFwBvEzUxxuz43cjRd9xwqVOeJk22g8GpoiFYzbyxh3s+GpL6a/AuWfSvxeaAmrKIO+zEZf
EtfrVwmRCu3ZlbAV+H97f+abCvHBUaDtYPUVO1FvwcMvB9A8XCWfOTB666q7SsPUUPwVnMHk454Z
nISJ2ovAZsRWeX2JHUysaOqFszfRzssyI35e/8x4Jan1H7Rjc7Y9Pu+tRR3LFKt2bWKALRsslYE1
khG7nR9JANzUAk/Bpc/8fEQDKRcTC+EJC3EN6Pw3AU79WqiXgGjblmRu1XtQWzwJTlJT3jYgWR4f
stc6qn4i/YxbKHk6MxImoCNLDiOMVZ/Y50IfXuXhcsENYWko7OYuiMJ6M43wnfgRg6r5gjdMLgS9
Vgkecrbe67DWF4URAFHv+1KRvQ0XYORLfv26hhPYv2qCsnpe64hzFmsrQzVT+b4sYxVw7ORG67t9
UEVmdl/LUoshlPG3hOsonBGTHW8JjzYxc4fau7uiuhptE1ud9sJYIlM8VqJY1lUA/OhSi6fVL14d
8CiLZMWKpXodNTr7ayEiJcbb3Mj364CuLUGT0vV9ljqR3aoygTYsUatqLNbnE5iUwu2lMNZaTOre
Q++hdDInyKxJXqq7VlboEDBYLPtbsm589avL+vgeL98gCB31qVUKRmboQ5ChI7ZyLjS3gp5NgJph
YmXFp9S9hIAFrC6IsSLQfinona7t9N5y5wl3PjpfiS4Tu19qemyt9jsSYWBqWRGVasrrizZJXwhs
dEV4n/K8z5xY9RqmQgYbenvSVbprptF7bDkXK9OIlhTRVgV1P6JtP/+K4+sbT+jWeSWGKyWvFozB
oZ3pVuvT5sURDBMRwpj2/WoknXNdzY1SOpMGMj8zvbZ/HdEf6Pdo1SF44BF28qN+Xrt9+1hICFJ0
QxQwj6urm0f19uQAhVc7+h0dQW1kxblI7HuCk+Wixt+Ybg0K37YVuMWyxy2I/A8zXrGswiDk1fCq
uu5zVOeqKgDqXeG50hKpM4wQvD6pdqOuW5X+IqRwtsbhSqrpx43DbGOiimQIvyzsctbiQPHAns2s
oz4Af+F5FkJtKbqG/IodDqtfTo98H6jz/I/KTnS30lCYxk6r0jVZka+l2LpUVDdkdUeTmDbVmZ7j
BnFjbLHKmax5U1+yCEhtefCToA84XEpdYpdXWZyIbiO+gDLw3xM2JFrOlnqrd/lXPbwIZwS3RZp5
C2oCvTQWgTzDqIsx4Gpnxcox3WDIRVVGjcXIfCDBCLU/IkzCYDBoGkI9riAH3FJma5BrhsIAgqhb
jsbjg0sVI11jd2NoU4Lgay5PAyy2vIyOhJrXAqXTjzHqT3u4tx+VGz3U1q2jGz2RfPiW51ktED93
+PmJgN1SUo/Ou4aqA+lux9KEnCa2yYZ77z54+jvMMsp+hasINfhmAjdpUEqhrRDcoruh+7b7gwrb
j5687t95G1jWaMHsNA/2F2xdPC2QVEkgtZ08d4xnp4qR1ZwSbzTj5L1RuRvW7uWXhJr98XwBPM5V
+Fc8HF5kcU8Kg9uC+oDHWFoTRepnQbGaQGmDfdMSwxH2NbTQFc1rCvJbIrdvFgJKr/nFYlgsYkZc
NlZY0omUA7gMKFNogUlwMAcgx9Y/T4z91mmL4jkRukIHpP/zEuKosciX3vCOx3xwYI22dFAajXGS
U1IabGap/xOOWQyN0VEm1UTsbNwPS5FIKZBQkiDy4bmvSuk429Xl+sqlpCBB0z4wESahGgd45jXp
qu6LVuQx8qT+Gb3/O7dALE7GSQCFW6ocxm+qDc/1kS/vqxHU8qfV4TKzemXrrWWrHPXgVgrdQe/7
qp3JeCZB3Ypn2znYdaSdpx7Zu/7tP040/uq4jrRysr6gD+9tr5B3MNSBKyn9+YXn1DFj38yF63px
VqeLnEz9lqIMwkUbF0II8ztdApzO823jjpFP7gcAS521lrkflbvuod81CYBeg0Y2T/1zDbCKzLQy
EHaNR69lA+hbxFp0K+uowpxVDgeCvb5JDuoHSK9Wdvi20NFCn1XijrnvraLtRtU+AYyU4QMiDuMP
MsdUU8MgAViubNPsX9SLr5xZVTiOiHBa52PNBokEP2mXUmSp0WTuEJRMZc97VwgLOYsjdcfagjE7
GDZZZoAsgCJotoA7Z4oIx51ICFHUPbsU29GtZU7g7oNnungueA9/AQFX6kWYeNqE7j6suPYGSN7l
/JObxNa4Bp7i8xYfGISRn4VYmFD0/8musa9mEFpQ7ENSVkBLx9wD7WzvmGvo6laP/9VL+BwerpoQ
XitybvXTbEZXcjsIjhrh1DLRaYv7XBCF+K0i0QRyhR6ECHNP9ZwbmDOT+jNzZPOW+VuCg07jVAUm
6BJvxbKS2R93SgEZN3wiGNZe96KtvUvWPmGV7CKEeiUIy0f3G835ea58QwoVZ/NEuJYUJ5cIbxJw
miG2GU+nooRE+tORUO7BdmOt1+6CiVFc+ksAQ2M/RwIJPVbvfk7AT6B1ACFotmRprdb3eDp7stMY
D3R0PAh0n0wAdNkCuv7ROrs9i+UhD/N41/N5kgymSjInjr10c+75iwb83xcqJVpweHn51uZ9i5D0
lmJueUxLtqzYTi9W91gFzxz/M69YHFNMdnXChw1lN+4gmVUg46n4PPBaxs3pGKtz/GmcIpy9GyqL
CXJoacraFBwPxjhqLNW6IRzngZU6ymZTGD76iwfkLrszgvHhnLVUBdsGnHrWto4YEQFXDMjqD+QU
pRGUkrJ26WGb0Px2G6l1JtixjdBztOqziL9NeSJL3BZKq0cEy9K3Vn1pwEaqcKgUeAk24GlqWbYM
EFkVK/P/C3IDtHRUTobYN3bxID0YE8g08y/OH8NRlkS/+3CKf6MMVwAVEziPmIhzkEG+7LEUHG/V
cxHJYsminlk8ZGlJpoEG6imbJR4285RTuBJK7tCX9JtN4/E0rFH8/adcz7it+ATeNvyGNmHRJj20
fV+xQPHqOVawzl6k0UPfVEDqfOIA4WY0iwVZGthTv/NM6NJ7MeFaYEntQsJ68FJ61USAfRh77Fsv
fQ0a/RkNrA8XLL6junwmDjEdXFlfpVVzV7+iyxjBLLT8wFk3Rr1MNJ9EkibP0spfjTVpOIL/N19K
8Nm46unfXK44JpkrQQ+RXCIPE1Hh8z9gXIQ/FEdKfcQKCvHGLX/+3eixkY0bx9b3RC+MJPiwIB+x
HiKZ083U968VI8o9uw9hphl2KENALA5cUWFLNlvF/moor33X1ab+Uf7inwL1wpFYDo38CQhd74C/
5ntz8sTC3uz4eKP+AS/BjNtuA5O9DKqfMAIiM42MIMT4FTnB1IwOoI+3p4FZkcgslucxmpfSPuuH
+4kNFSeTLpr7+fFMWhyzON4Z98jtKlJbVTAIMjCJ1EBRfBbDqdsbBwUDmE6bmwB1u9K3KliSigxz
9Fwp7851+kx+yTl5LsYop0M2Me5ATSa7Fh4iRDzymHL7yA21VcUSieCnjGOIroOIFwYAKo5r0izg
UKaoBwCVG7geONPQfVzBJjLMXrOZQGaf6rvziFQzTGYNYLmFQp1lpP9G6fV4xMJ/pOjhTZMaQbRG
B7IJUYZTCbPWuHJa8/0fvVwJp0khaODdgXRIHDJVxxNPXZrAK5IuR07I+D7FXG9Q/o/c86+JL7C7
/HNzmW3BU+4BJlGWNqaHDKMJKaq2IJaRPajacVfP99/FmYehgemlD5j8Mbiedq3t9cY1KE1Lwfbq
8d2AIFK56JVtc/QCF7Z2I58LuD8G8iyZqu+jhS97wbvDQOyDpTTAqPtaeP+VcZ2VtU9kORDBjBcE
Pw0iXYE1QUyBaZfdZSqJBNAI9lzJObvvOzMijXD2XkRaJ9ETvNsQz5E0xvdlZPy0wuo0fStM8ClK
Ip4fHzqW1RXc1D9qobRRiqVfOzDgwjq7n2mdHaUlDh3t3WMYl5lRhYset65KEwf1fZXXn/NP/h8S
ZJRG9WuKXTX+BGMQLTSz7PytcYd9YWJpjq3UlHvvSIwwucvUIWGsOMowNLRNIbQhUuVSx6I8SWBN
qMR07wDtOXktVON2f7syGIedDZsYvXWSNVVolBQ8xEJaOO8vFb3yr8YUoDIeithcpbV3A7BGkSsn
d/lpE0km8u0c2m4rkVWAN7cHIquaY69UO0NOiKLnuARPmQu224YvxzJNxurHMvl9W+1oBJnBNvo1
gNadNUNkrepdg/Q3DdXdmd5iScuJMhMC8yWlqMhgF6NeFBEcx7zkaRTjY06TVLDghZ+ebuJMwEyX
cBgFngbVLq3DENXGHioIvcr074wKkjF1gYaYFERQmaCLZeFd1xC+ZoEvX4p0wk+d+FVTJsH4LgPY
hQ13jPjcGWputxP/9YApy9eVT0nx486Ld0QrBi+9qv/hrfpynUbOzuAbuwIhRLTeVS6KIKyN2NFW
NQac6Z1RwhhkkSoNKtMMhlHXvieP6n2p2vznsrQDUAxRBnJWxvzd5WLVZGto5VP9lT1QdS1vh7wG
67tXT8QUAJNMeQBiYNW0KYKPDemqvo1ShjPMRcVhrJ0bzpmYsIoncHnqWqb8/6zHnMQrdtp5dtsp
rhUZ/5Vt4gx0ZJfmaTE5zBGKPdyx4kOaxmKzFdBb21rq+Ypdaec+SDsDpiy4G7zdkRJQc961+Lbc
GGKEMU6cSYRj/R75yk1gMbZnm9kOru/kfPiDdDL2fQG8LMbYLZezcKrECY9nd7/tgfScHfBZoSx6
nSJLDPWTAPBvOuAY15cwSEPyBNfoNrDHmRhwvGWLOMlG40h5MSw8uto4MzQrNiS9zA+kHYHLEz7m
PbLKW+8jQtcJxN4fZX78AlCCmFBX8FQDDsFR27siVHEiQS3upPxfzVb2nzjcAjBVIaO9xDSlE4jQ
fjiYfB9jMsZJXkDStIr83rZgVLvj4Ubwc2o2pXdBX2wtj/1kmS9OKhOU8pkmXYM8BuDiYh2winxx
dT6sPr2ORP6SZbwK4Q2UeecXXqWfNJocm1r3v6ISFObT5SrGD1UVKjC4Wx8PNY4EjgDcjWlTIECF
zEwsL5Bgy5TxdoApgDiFWAq4xLU9H78yijX8IhhjuzpWMA2zxoLBo6NOSkFOePmdqz3GO8lIeV0x
xIriy+PbkYY1cMs+9oi1LyPsWlY8e1lkDn9gqVIaMaBpdXUSKOjk5cp1rivSRI8XpKAo/ocRqb5W
swk7y7cihSCr8L9m9ciCnwoUTyopZAb4uF7sUy1KzcEKNgUjFztjzPC7cpYmQ2P7Mjhj+VHz/VKy
nl2jZdcEUVq5ksXDyAqkINis8aGcArPr0TTE9FIIJA+IJYiv6A+ir3vda7slpFbEJId066LZ815/
e99zTy9c8oyXcrDhjgHCyswc/iziRlskXqPxxzgiI03Mc676B6iHyMjwGgXak2gHHR23dwzQcTMM
Pu+DbP0GSE71/twugssNSbxRR0Y8xPh9lV9j4IQL1TCjtSxoUiopOBz3nkWjtu0IM+dTz9TBFP7g
tF3ObQvxAUfRODrI7Ch9gsuS3jgzFPLtSfjKJ3Tli67l7d2MaOhcIwhn3P0odfuoWnvJQXhBpTUd
bsE1HMssanYrFA4p85bPHenKwbOz/pDv7ADdn98A6sRy3nZVYhA9z+xaU1wN2YA60cp9h0yIodCA
Ks6pofIFfi6nHflTfpMYAjbQ+faGIO/bDCDqx00hb/7S+3fVWTo2fVwrreXTGuHqbsdyieODc8Js
OSIaSoaG3KpXL8D90jxcksjK8bguM+8Nsho/kGOrv/8FuygNWbTMjR1lcJetpWtjAy/34x+Y22so
kzJnSMfuDETrR5PyUETZ3V3XzuQWbQG4DvsQHMK+ArgumEl+RpaGUVr1+Uf1MzTK4XD0qpTPPx2c
xmVgFHqUXdLEXpYaSsnui1jQy206+tWxjBCnU9QeuzjYrxImfgSa808XnkAB3Gr3BCYG1dGD2VVl
VtF0i7A/DAPYRHiApxxLmS3Rm9DcGhTmKUpty6vGaaNtKE8PPR89OO8ISh33v0tB6gDI73AKOodA
m8Mh24PwM3oCBUKxUmoeArpNgmfmjIp0fhlnhRUxvxaN1M87v5Bu/tzzxQpQI0pfF3+JfmX8QSao
8rvrFthgbWBZ4CZrH4GroXc2/PUi7Jd7bYDN5Hrw6C7LWyLtsHXcByT02rP9uE8oUXtSAue+XI4k
mPNMp2KEQbRhpUeOtGOniCirZ25y6IFiYjh+sPy0xUnAaCUrM2rddNIylb3VSiBYJH6futKGU51Z
VSjkqzaCvORp3gu46dFWd0DCUe40iM2lVlp8VcSnOrr+l599gWKDbnhK46NS8nRaroIBPCA7mot1
C/pSHemBs8vNAInz6R4PCHuPMqjEvyyBTCbwlqnE/fjZF5VZiPlSdgCIzF0mjM3VHiGUfAiLhnS0
a9WajXgadjENF7B9y6pbMeXO5VAJKr/P/f7vCVbRkOhxXIskJkkVWYIfyJRlcW+KtMdOjRValaTH
TsUvJgwwj++ECKvjerf3G0pDbmqxwgbx2+VEKdF6gqk6miQfcjK59H8oPbPqby5fIoQ2YQAUcMgX
R69p+euzn6Ejo+q3HAtK8o7IFCFYZzZjUqz+VzA68cKhI3obMW76KNjVEQu8AImAgdMOy42govOb
2ZAFMgeKJfK/VnbUb8lnE8fWV1ST0Y/tSeurl5w7kPUDmcL5mFVB+O9FU2js0vxvlOLpPpWo4LHY
VG4ujOkY/LikGwhauHp8Jx5IJjrB86jEBYXi89eyLkoIr7hN/0ip/1yIEKdiB7Iubd8WTzgiEC6h
YrMqgc6nyKeIJ85a66lGqPxk8yQ8QMFZnjslLdk4FDicgjO6+mf04ypGldV9+XozH3dRDBVzfrko
PyGmgE1tDGKA1ukLEbWkGXSKYTE1Q8mIaKRZrTP+Tyk53X8E/9ctiVYrYLsircC9Z2pqy8TH0el8
UrwQIQhT9jHVGDczaIIyqQrwZkrfr6PIiv/HRb6OwzpSbohsLhOhtl54E+YiR0i+EcY7y1w+/iNr
7peeqDHYxMt8fxSb3dgu79P8qGcMyhHWM0koYy0tWAj6zqYNrRMDhyIynD7YMrSVCTkPKjCNgH6L
AabFg8dEW7KA1r3GtxUI4Bt23DfAVE8sSjn65opAGNZFr/yKQq4OOnAtWK1PKQgk09xhiywEYNmR
4PVzfXbgngDWWlCl28j/U3ykzlwHEa1omkpfr0aKpllWRUtLFxQAwl8heKAW4a/2KpTaEdl87sJN
RuQ+hx2+2euvP0H+ASJKWZpSMHU9ivEIHmrF75HtcjSekovlZ/JbRF0ReGtpvKmvYWkmPqz++FJv
25wCrltlDkMqd2B2x1Zwrus2GkNJfFQ1AMCDmI5BggA0nGy5GeJqyXEAPBiJv+avVwoBfZ7mFIMy
G5S4n9kVsS4Bsy/8vkj8wo3sWMzVYtEEtClhZECZYpX5Hhpw+cCweRjqauZkyfxeoA2lxCQ73CJv
eNW8S4qx2TqppVfCQio/Y6MV6D2QGOUH6dxYOWsdbFRy//HOoxOhFkCUJscLTrnD50q0OwIpnSfE
6dcX6IKKcZrTyM4Y4rZV22yJIKmDzUnKerEg4PJTutfuyw4kM4rjOaqLzPh1JuYtFBwT/zSLuafp
cPv+a67LaruMs0Top75duVTDDEznqHfRGTOQLoyGg05iEF8ljGa+4tDI4QfV9QFkwmwBmFzdDcpf
GaFgLfIBLhNlp2BYIv0h4AwBBG+vwME/vjFc9IOzQ5inGv2fRdjfZkDGoPryZjNHhF4AiUXG7Kyd
jzvfd1mRC+MjABrakuHnn8Cmp4jwFxiRdwl3bLUMbryH2iVK8i7ZxB+fSa+ccJKF34OtvVqg7pAW
DZgoF0rWv3qx6rVkCrP5nPBEBfVkhBtwRPkWgn4l06i5lDZwXVw6mXDYTaPIqlEE0PZKKaWGoY/o
gk+On3/iuJzlO+GGx2WSoqZu7I4P31aFwU/rVrxF/6UIifLQb/Cx0WCSQgaJULxgVlloUyuQTJsI
57AI2cm4xSX1XTwuwgE0QXw2N6OsX7c4tN7kh1dteduJHSUGR1dsXgih/kdtgQrsgb6WmwCiJRsx
tLK9E+ALtWJmZyTQPEpuS/XZ16Jn3gLh07gE3Sb4xJ1UweUrleMM2gArLsk7kZxAGyZyOtBmJs0Y
IcJFIwdCAdjehzjvr8cfZ7yguAJYJ9toEIvSbgm0PqDvz56LKCE5Fu5+/kVKDVzX/DdIT8X3a+da
Tm1acCx26P5bTXedJpew5R6PQuBqp2Pl+vK83bil+s6DFqiJ3NJ5NmbxuKjgGsT/e1Q/b2dFYtRt
lW9uc5lWVf0oH/NFPHOkjVa+9Oiv9xkt5GJywN3llg4phE6psW92EKokHeNkTkRK7AgweDGpq5uI
oUov0peywQhDnO3SKSRnqp8a3hkbPn2RjMIyk7uzIJeZ8uTqpgAZUSJD99iJLaVxCHq5ujTK13EY
+Y+QmWTR8Gnjd5DomH9eDg6oVtMsy3GkGilRCSZiceGXNjwDe6Stvnnxp9SuOZz8aojzcl0HuAk6
Gx3tOYR+c8c6WCEKBL26WZLeJ+DlOdrcOmL96xRPBJjzrajh+xASqS3/ERzqA+ufRHO6KEHnYkKk
T5fsT6OInhSj0KrqjO7XuBkv8nifUc5jjGYIoqKQ/sf1jpOXX7ot24re+Uvwe+uAPMqPROi7ZWGV
xme4hxJtwEQolsjn4npCPvTuWx3gOnABjJrOKorYSn21TmZkk8IzLOxfuY4NokjeF3rp/z4CuwNs
ND8HvXTZJlELpL6NHQ89GdGIWwgmm2bXFKJUJPncuW1d+wJ3aRtd3FhUZtSQ8MuVSem5O4p3b2/j
dRl7d6q/yboVjFp13PUlPt0CfHBT10LzuwOlChXSVVTWiizxpXsQdHlNBszZ7mLpGWMcEvpRf1ov
5lGKRQN2+xmSkasBfvUcAsHupQ48gjEfJJ8VK3x/CJVh9BwRJSf9Vt3NWuaharIJ68KMACoi75T+
J8Mkfl3l38uJzbFocCRMcbMtmUXNkQ38GtiH+XXe8CRyqfhAE+78OhJJ4zKPuoMBRF43diZ9AMd5
oG9Ja1LNQ9+BWUY/GeNo66hKs5aXKZho0IpIunCIBCUSFfAp7ehvSloKfptwAsFW/gNz3xQBxAuS
ZcYQ2S9w1PB3+H9TDBWnPKjgcQDa0PuLm9kYbtzdhCs30GEX05gG7GJLSrsYIsewzhCEwPuxHQGE
OfdN4nribZD3CZOKoT5SuuqNonA7ajW433jDDW+7jkdjDrjFHUX5TYAjbdqdjpLT+nBppV5aKIKk
pUa6ZyVHzoYmpcEkc/R/QkzfZ48jj5AzjAXcWVbXd8zfixwHsCKmLv/g7/X5nbxHTyEAB4QcpVWo
Ug4JKX8GxH/D08d4OZqBG9zZGTIlpIC6nLhb+hEe2vMipD54X3ccdkUoniXFVT1zgyzBHhPa7Niv
wGVLSyWOJs1B4GbMVioG5feq7nDfxH0moGROVl5wvRlDe9/dNg6gbOHvxzVz+C3ThLF23p+l7sGx
dJHE9OdTeh3AysNKU4iycTHsWtJ3DrGuZNdKNBEL6ug33EIhsWnMbvTU1EhVjNGcKbm92KQU1gIg
/sVMoNedC44Bso3OJKo0OcQ+pP8azdwgT4gUzFSnooWYacs7vly9pOFyn5V5XgIEHLC2/x5e1+wk
qW0GqEDf8ULvFf/pHrUg9JtQRTvI0oFhoVXWEXAGCap1b2/uXCvfuzsNLV9XL1uuc/kWb4MLo2hb
YD/1WmcyVBpL0uJcopI4p6/FHUO0KIdVzNKpmG+DfiFpxokMlPc7dIzKRYssWDgzycuEDxUlWqAM
HnG4gzgIAJE3WwSsvzU6b2WizVbHrE3qz9BpctHy7Sl9JsUsPW4vGDCowEECisjZK37VTUk1Gs2X
I5e4QNwiaIrsrk+GXgmUCpl6MvMEw2blLPbYoE0bKBV2JrOYNnrGe4rbyKhCVJDdlhiPAc2pwdR7
N67spLYUzKPu/w1RbslnU0mVqHpAR8W4wkshmQK2XN+oGv/02ie6wLav1VDG1jgU3yRnl0tGRtTK
bL8n9szObBxteAy7f5Xvh4hyewQzCvME3VR3z0dzEpEaKEfw9F9u/HRgQ4VVMx0uzWyeTg94WF+I
nOWHnjxffNipc9N8lDPMRCBghfHzExkXuqhnRto3eC1yw29SFMN254rpV9dJJ6PTq9MFF0xQ1TJ5
zKy/PgSGvZnTDEcXl3HYu20G3aCNhAwBcmJo55BIwfOVdHv6qYuismboNlSrTumHiTaAfo6KGt7U
s5ZTvpn4BAVWCOZB/nkHQlZUNXYNEWz07gC6MaEM9QOg6CemI3GiY8lqH3A6ocFVTPDUJgQGA4ft
Pllc2b8cluFfTyLb3F+pd/ta9CXHPNX42iaISU8cC7LUff38RpHPmsCNzsAN5tUqgGP2VK4CBhNm
iB5mEECiUbP3cN7d4Ylybb+5MxwjZ3+m2mz3PSaXixBv4Oy7MUV/DfEHr6EeWNpkr5cEUZDaZS5L
6Qv256BrTbjT8pxElYKjc5sF3DyJCdGYWWtm9ukFKoEJMIAnJdzaRWzHgNWdaQERoJKtcoaG4EZs
X7PwEprGtMdiW9c7XJ638mxqbP8VOEdVkcR16vdiV/O3x2zcUSr3oucA+yX09XXl84DwAYkQWf9W
ku5OXOzZKnS0fnXnLjFHkPANmraNSVGP9E08+SuLDyotEnHs7K42mODFb6sXGQdd/tF0M0l6+Jqh
gGqT6uEKuA2XJLq0omxHf0n35UKCQ0MIKhzoEQ6gEhVneK2tqygtk+qGwVBz3DYsaHI8sw1jM9Xm
b+BVHeQIsGwY3bhZcUbgkI4w74faMVP8SxTux9pynsogA2peF7s6ixuYKpPtslwG9h56k9hwlKRY
7wQYlu6c8+aZYBKtjHx9iLHlPWxTH6sEgL/y0QE8/8ZrFsdJZbiWhmrU9Me7IdTjG+MIa+ClGn1o
tyoLEZV97cwws/weboqHs33MdXoKCg7PbRJYqG7xf9YiVFeugDkxb53Vy6uNHtMOw80xUMwLlfJx
ZhIuB3Q6PE0YHK/poWWQljWfyM1nIMBAaMiKSCE7XXAeuy+/DXy6rJpB1/bPhwhfLez9+GFbBN0X
sKNsmLHd2PXbRXeSdyBxSoq401BHFDNgCqWB8y9rkKjjAJriX4ThBtXarPV6GHlzjKHftv7NdtT0
iG12EHeIhiEXlvN5w+8nzNCl6yylYh/Aph1Rhvd78lHXNS+X+7Dj8dLTkKQSEBBjrssAAo9WwC0e
Ehl3vdo8yWM692KvvoAep1EC7RsNlqDCdKjwksg5dOeaYW62Xc1uK5FaRjgRX8yBW+MwUNZ/hMDr
MxZT1o86oZYNQDw4gxYab7qVcRp1y7Ff/CkcH5HwD1CzB/vJQUJPFsNhudR3F5h2iZYZ0jW25BQ3
IG8iCwl14C8JRSPgbhHR0cnhycuG/Q9b+MIaAcxQv3hhjEzvQUWo1j5EJsTlBAU6C5zbqCvb9OY0
JEtizJRsX1AF5fmfI99forpnchiSWu1Y1EdNI8/BaAvdgCOJot5eLphNgySk+GI2EqRl73LwZJqH
tNbk3XjfmzaLk961nqL2AQATuuvwchBnUjPJkBOBE6m52ojP9x+jkcAjxjKJ3me9qTJASdUYPRMH
8wokL3iD+MFGkXfkZvk36X45Nq9Nqq0qG3WJcNSYP7oV6e5X07LKVloHa4e8CWp8vLlpePljl6KV
7jSNe1Rn5+hnD/7jcK2E0fPBYfiLpOD8MDMlKt0WbIZVCTepf6vXFTDHXtmCk4M0xjRmGQuhCH+Y
kXyoLtZxictVG19KnBP3WuN2K0CC0BWr3jKr3pm2G+5lC+v64HZHSpyZ9S2PJX4olcEPcqT5dhX/
TxmKJgZhwAj7Z8My+C/Uxh/VOlsrmpq8JDKEcWzGQ8zkUttxCwY8cvni/lXZ6w0y3SoqrKZUSwdd
bIndoSjH5VkFO+CrWa9DFHTLDUyFiBx5zYgxMR5D6Tthx5a1Fe7SAE+diUu8rnSYpA146jxqnmXA
/NO/DZdgoJO7Obb7hb1aoi8vlao+o0xPayW2MAC9ZEwTW8hBIhD6xDTymMPtV4nnD47aFEUK4vZS
TlcPg8rs9WCYMlZxAGuDmtk0y7bObjo9dI1/Yx53MUgVh3c6je2kKCa+Hm2xQqzZE8ZQuaL6JgUP
FCL7JfG5e9SevUU/LopEUBvXpdGBCjQja4X5Ieyg0lIjM7Kd7CBN4rNpj2y4feosLhqRVof+R9K5
cIrrKxh1+kehIZn5tio2GXq+5im2AQQFKZVcjJC8iu/1C3R+ghS/CWVx2yilvS7cEw0yqv3LQKIr
WTNyx/2oRneeP5x98STbFCk4OYO8si7KXNeQs/YFRho8TtJkIRBkxaJpcqxGum/QYGKlBIcx217F
GUFDJ3fDOA/DvQa0CSiRaC2jCPMXNntLxxJhZvGJP5540t/yZaPXndLe//LbSxODClQB/5jH4Tnw
H1T3bW7/nhHJhy4EetBoIuJGHF3UVsTVPGn4Wra6CVEYwQwopF/2CTkPlkAf8p0i5IkxN9RiXX66
A0D2CAuxHyLDLppfnzXvlwQUgHpzVy3Y+Y3GXLaKfLPzvCiJWaQ4uwlKuU/Epwgx0aRR1pXgnocD
7qFV8xhAojFCyV9h2suYbJqLOY57h5gN3B6sMGbScA8xjB7nBc0qlyZSzW2suqZ0SzBPToub6En0
9zwO2IHs56JmNu0WPm/YdPTxMBskAEw1nHmNGYQbXvAgTbUvVy1hQ0jwyrlibPf+lFDhRoeR0BhU
XZqSLv0MK1f9935YeQ12HOxtXHwx0ahS3KwEJcmBr8gr2+3gNoq9NyzjETJYVnOygUablDkzjKNC
xMyshWHCHxAaXZJr1Lmm9DUTxAZs9LAUMgWByTEJfmFwWOyKrjA5Jab4EPZ+ZjagBR8GbqWzkMXf
ZOjD8ebvv3y0/AGu9i9NZZbg8hAtB7mBTihlcKwbC6DSuz/MZFJwvjo3YCXUG4GPtBf2Vr7c4V0f
SNWd4bI+QSUYfVBdqngxZZ2oZ3qcQcpBI2Sllw7fRpFocQmLKR0j2MAld0gwbQrsJm5qpcbdAnP7
DTTBDphX8pzJeLMJhESNSgYeMqB/jtZxkTeLitGSv/m+8GQ1q8WvHy1cgxk35FAvEjnzjJ4gX5FH
E3aCU+bxT1IXkS3A85f0h29/k7+lLD4ISkFgvHTT7cTp+r/Iym8tA2vxyZK/kJu2c9+LRe7TiiCd
AuRS0I/m+F2yRsyBfJyO8cJE5r5X21NeADh5ubjaacPBvWUxA7HU78J0iKdIfce6FFxXRwPaycIh
8XjOsGGQkF3mj0Y92CXutVYaC5zFEBtUofVob0QiXZ+ohei8jeo6ng1Qf7R8xUZ8FyAynJSt6jCT
KIGfulqEEKkwtyvW+J+pdNUoXjvpKObMi+wdF0FLD3AxiNa/Q5XyK9esr7DtCnbs86DO0EjdMpw1
Aq4VGWH5ZLWSu2YayMP2ppda12OU2gZlCL3dRcVY4f65Ne4QF9jQcWleDmP1xP1FzpMBNldJmzy9
4BPesnxMtEQjYgzqnEsFW9nrck7rEZGs3u7j0qPb8k2MMNuViJJFOYQ83lnvB+cNOOe8M9FkR2NP
ri6apv4I1H9C+3q16ZMbUICqD3HWAIzckKUmW0ooGlgZvvzrtOqy7b7lG1VKw8WZNvyc1dtUomgQ
M3RKgZq48+NE3qnl660cBPQGO+EC4N0n6ElBOw4wujDnYGMhhkt3XINbaDBSRtjPWaw2jiPyQAfm
RVPB3ruUuVCs78J8kaeflTLVtAGxe6ZkHFT0RHZF6Cbwsdgb/GqZ65E32K8kjUW6QcvaurRz1cQp
9Aa05kJsjFgP17Tu0WT1a9awMsECurSdjSzD8tUtWyWO8RDaqoI+3UQNEf8V1fGyLFtcPzQkNulZ
2tysE4BNfGMFUCae/dEvKDpy33JJ0kPO0sdmQd+vKrXnFgiqVXnp9SiXfiR1yHIW5ZZrQgsPbDNV
N/zOmPDEOY8mFqZ73BbFIYjF9xJa2qFLXlUxZwWvUmSXdOQFOKuucFa0JumAUvQyk4r74Y1QESln
TE5/+jpeJyFwRS2xR4CjdI3FvMX/h3QvkzuAE7x5yQoHMB34JdnYt56NbZ2Bv23j0bWc2Clex9NT
bsu/8OK6mzlpmeksVGc/mUXiOaiUHovoN+qnqjoqzWP4QVPHO1kPnGVzbmF6aCX86Zx8trZr8NzT
KC8c/6S5GNrWzWNVmhOLNvCoXV1N31FvDCE7YM42Zvz/3qKVEY1AOw29nmOvnOC2xWTqGjklESqH
rvdUAXp/j6KqhI4yXJUEqAzP9EfsMNz8InzNEZCIpp1Jr3WXCGcWDLGkqAqUdQuwVlR5B64rgOXM
422okBAWkCjQiWNSg2GgtRnMtD74sNbndQDMar6uXcn0rREp9H7iblc9scxU+jTsdcrBIqV1e13m
Bg4sNz5dD6B56DanxG6OwCPgUjt6OhzGQSK9IMmxkLucdy7XbKZncPqU2dyk+EehXQ/RbC5PD98w
UJfQhNUYnLZsffb3cuRSfAYov25hm3m4XhgT6CA+2y+AdudfDAYwGSgdn3E9p/RPS96Zj73hSTtY
ezkdLXbZkGtP5E1cZROsWBEw1YmmoicfyXeg/Qlk5w7zdsYLuwrB+1ipvTl8c5b410vwZyFMS5uc
IItD7Eyfb3bO0EYbLWxKXWCUkNVpuhXKz/dv0qDSXLGI4dacEyyeYyxq8TchkFrMD7PbDDRe7UKv
Oiek/CBuiNlflNbUm67NapzCnVxDI6DeGODKq2zg8W/X9NwXFiT0DLDt0pipyTcAm7LN0oJ7+za4
SQC2brjl+ppyyXer9O9H/ROfgHAX8s9hPhNM0UrHEzcfte7JixPzhiPyEqxOt5WJ1WzZPJpbixFV
nQ8TvYKa7UZ5/amBFlkMrUlG/ift7OfLULGTr4pXToFEiQjlSfdvwxmwB7dVlYRxAMj8YrHuMDdR
Q1tU27jND4mkWyHrYSZe/pQY19nKDNMszPW2SHn6Z8XRnBtAcngNtYjxBNdt7OJK3qiP0hnyeahN
ktiN+VcK/xYDTSwpnTHPBXTVLmI98dgD05ie0szgisRix91lyEyIE2pxuUNlwkXTk5O5TFUp4A16
D0WhJS/HEP4gNZuwMB59b7zFOolIsVCA0WInbw/ci5ZTXtDGRwSz3Yrtyq0CgQM+DXVfDIh2sa1L
0dIdrnQ1P2MlqN6QVAbijMdN2Wt1kot8Ly2HAj2tZAAamcxsFMDwauje3fv3/unPjgw8r/Buky7L
+9iLpK7wE+4K4YU2LbsXlXDUUno/iDp8J+NZo7e8OVgWuI3DjZLloT0B23cGL3giGMiHjpLZaHF9
28CKFJF7M1lQEVEyAMd6v35Qnx8M4EEQIxVl0k7bQ7b+fJoklR3s8AMrwEMxJbA3X/fvuPdmzuK5
bsnWuz/30c1Fot8MypqVd9+fCgv/MuVwKXf2ww8dfK+lIShHD9W+j91GY8LsLOrnksFlHlqOHywd
dM0czpcplZuWDplGlZkWyOc3rtHlTyQHktjkRuGI9YcXs3DsMQPcjtR8M1sVbGXpOwyrNSSBHTip
Wyv3Erg+ZbrE/FposRFOnzK5A6MRgasIPlrl1e4i6glgmH2SHmLW4A90RFoSJP+g0R7zdYwt9ejK
bC5llpPs0YR+o4KoJLT19f4rY/aywHZ2Uf/1M/Q4WEASHV2SoJVAHeccjUJe7I34jH4gAvXY5C1L
i0N30DFZoClaj9mIZR/Hpjtr6e2sSd4GwghXy091P0CTpkGoRU9qFGa4gP1HAF3TBF3AkY3k4aNj
vqJ2nb/IdiL+PkT2TnwrCI7POl1v0o/XEf7WozvAmuS5luYmXDbBYOcfip1mgqz7+Yjt42gWjFjt
oXzK8GIrtAGp1ySJ0949XKdP0Mx+yZhiMYYlofjNxOV/UjKSfhmwn70z0T2VrEHGPGtDm+My9Y6x
ZJApvKBzcTmx2r3McH2/P/QYXbOgFTXGS7spe0ythwtWQxk4ezXhwDi9IWGOQxwuxTOnyVbWgbIY
jEol0TccJLTjHbEmHAGqcItFNLpHDqGE5gM23VZqv90KdRz03THUkE49BMEWdImtz72APqpxtH6g
gpeWroTfyPNocRCHA/adqLYuNMMV4s4wSBj4zTlPAVHYXAnFzEaTajraAZZaKtMx1Y1qQDcFBhN0
FSsf6g3Ef3+ddIXw8x2uNkX2saRUlsDIoWkgiGMcm3vpAwpCHvmyJcwiKj3lADAQfo0dz8I0kEsx
XtqaPTxVQpzfeclUje5/gbZTj8kpbQluS/nFAIrViUV1SmqRADnlK0e3yZEigsKdVrKrscGDaXWQ
DDyYrSj6kRVmpiwR4ADuneFC2gLp3bfZsGQs0lyh5HkXA0dYilP/+VUJL7XDMpVuBoh8mCX/PbKC
GXSAns2/Syc+zx4nc3Z5DJM4MLIv/xx+MB0lqh+qum8tiQSz/HsCNPe5EW5PARx3s5Hj95S8GaQD
BitZY6CqIzDHtBfoG6RAooxOjY7HQvEGdC1j4Po7TusnAEhJwRwz4hs3kpojMP4LJePEhmJePPXG
wp1FCOMNfnenIT8Jshp26H8om8hcJ2TjtK8QQVumarZX64nebIci73PyfdMouCWlpxGuIkd5V3SS
jsIQIjrxVscHFl5IKPQ9cEUx6zMA+9+D17iX9kKpsc9AV81g1uxq/iirU6KLdTyT54EzDaXva67w
/izCYRGtWmGvtzo1qwiLJAdV0naR+LBsMTQiBKLuFC9XUXKTgcHq5z7m+/YluL4yBzGkFaKsW0g6
LtQl3Kwk8ezsEan6vYt551PGczANjIeXOeL6BWKqL+xy5inge2Vo9kWUXXmzdCrXiMVE8LGGp1dp
j40j9NADigShNEvJ9ozONEt6EWaoVFf1HZb1GC/S8vDdD1t4pV/NfeTHnYFRUXLpRtRk7YllbC2Q
er520ryZFdzIB6Oe9txQCMuquOw3fRitRoEogWb1ilnsOIuksmzAfOb5BwXUP4fQZwnpYgmYI5uX
RuhFv4F3uDpNruiE54k5sz+AHXMuUEwJ+w2Ofl5CHLaLfK4Xt5aKpHk1jgkS0kKOlpcDYOuoGKgQ
s+s8n4eYYC2oL6wKyxZHGdMaDbtKdHLfO/VX/nZ0CTN4vJsvsP9aat93R7K17gakQEvzZLFy6nAw
UpVRPfIqDqGSDDB+6hpVpLU7RPq7B8Gzw6MQHzun2YXiVp5fn+29a0ivxW9hErWt3Zw8eFmbvhxn
Zcrqrzfz//u1gLFb8TAxxGmsg0PAdC7f+qeYn/C3n/ZFurnmaEKCV1TReB2HgjDG3U1KwOk2l3kD
qHAjbJc6x6RVaivPbDlw804b+RS3zVnurioAtOZNjU5mOTabbBs7eXGcM0d1ILeGBr2hc3DXa2bT
lFlPSka4tV5usXLRKjQKu6tGhiqXwcz4cB4375gbIEkM0rl7VwEw0zSRhJjaRUm0FTbPXOpIdvTb
Xc3bcT1v3O8yzh7x9rX84m208hxCHfEd0y+YzegnsZXkrFMk/G5POejy6J+ui6NefmVfA2JS+9KE
RNUjy/5nrgpbK94vxVd7Tzh2+LtlOHgqqNxbes0+cSWNUKlcybTPm248zPZAK5GdaBQNjQ7AYV6H
VtOW5VGRvRH1YQeDRbUAYV7jwDm8gdRNirUHaJ687tEjw2P5DzHNrZ6WA0u7/kyoULS37y8kduNi
DYonAnglmQCMTSToKXnx8X4PRrBO3X2xS8koQsGYLW0fAR7DdBMGYkfn8MNFLyYTE2Yess7ssIe5
3FqDvC90npXvv2dSuD4Oe9ocukR8O16s7cxOyPCe7oXiWARXmZ/N8KPy0c4JRiJLAaZ3tKoPndnt
zQx1arck2T/EGc/64r81GPCIYiDRw3NaRitCf/MR6fMFxSzUYlKShZmyG/g8i7nwf9uQxZWPjYxO
ZTN9HVhve0hXxv2+E7M6+XijYSVkgRmZ8PwrT2Zr6ygcWbXt2xAmVGlZ6rrRWQiCL5N/++4TAPC7
X6OippKc8sVRS8NuvxL7igmZwl4EfOC0Fw6oI043IMEwTWrVlbQTADMezVKB9LZ4KfZ0JfHUzR10
IozN3N14RRRusSGUOjMPCRYRR5AyVKU34IMbO/1r6xOw8KdD75dT7HWdWQn83Ajwr5p1Drm3cxst
ZqmhH2BJkPfDZdLGia+sEBjWChuqrh07Uu0d8wGsNl+oUI21IrtVixjG4x+9MgMLPEuAT6wPM9Ll
qizfRAvvXBbgUg+rEw+yvZIxR9haKvnNYgLKadD/HWqPt2G3//A4fahMhrpABh3pSdEAFHGPen9a
EjaHmArq027hEcytobuJ0iSLplGXeMqtBS6yxvcN4lWqpKQuVpn5AeixTl6QAQk216SDJRjSNzgd
p83NaEtlKbhsjZZowhFIrbSMNNIMVoZsR7WimJwB9s10Xa9u2Eait9qaY1ERIHbdR6Bg2J0zVEC9
/g44SIQ8lfslSf9qzm9SdPLOHjVKU7Ega1L2hYViVt46tS+Eqo8qiYIWaiDlNTPKQSYhAf+QRnhf
7fR5WNuStXQKuWgzNb9U++fyfiH3g3W33zRUttrzBj1b/7duTZWmJKKwjqcpHFDVYl/H0TSB0XZj
5+tvwaL09gb6B1bHjM2bCcVVBakeMnnFespTeeOTDpM8dXpx5AH8plYI5MYdR4MH8D2+YwH3D0N2
d6FLfdigUQTz34hV2FsWm+GLjsjWTbj18NeeFfCpgHl7btoJBBIer2mAqrkJKhTUsvyG+UrtPRGp
AAPpfu/LSD0nEk5P5/8Nt1fhxvxAY7G3Q92l5DXs3PEtyNVyq2N8gZSP6nshfjZWjynUNZTGP4Il
drYGHv2udcTlLCsdZnUJkqb+ON5Yn01UC+cje43Fzddc4tyYZN6OcJDljcmilrQu6rZUZwN14so3
IgsSr5GDlWCKmChr3wnwZcfdq1Wys+dd0+22CC2Zq47IVUT92uU5u4BJryYpmnRjwOKr3ortE+Md
28ZaPGcRnXw5gFfnQ7nKr3DibugFGyey3H59Nt1QEHJGj7H1pemy8z1zrYKw/MHPtV8jl3E2T1Cv
bynGIaCPCcncbAVEhBBzK1hMAR8gjZ5ShMENEqk1dwfgsCQD2lOLK56WXOLTf8Ykr9CIpnM4PZiK
/OxRbJTwIiUsDSq/5QWcry4JDdVzMEGCOZu3ognA66aRiMhdyRu+H5vdMJ6FUcMq/lIpTzu31r4T
O7q9shvS+2HqfCgY41ANlxcUzG6t9R6sZumkHdteNpjx6G7bcI8LIlpPSyrhSTV61AB5v369mAaW
JJgENW0Efl+x3bDqT7OzEsBQu/yPQicboEMdqsdD4lBt5Z73VlQOTWO19g8/wizpJNBCy4yQVZVP
zongOSvGC0uWoXcbRqZreGMGpdWSZNiZ3eTXEVZwufJwgH+zF4uJQ1swogTQ2iDBgftkrTPDsNad
1tnkK4PeV1+Ptf3CPMo6+blPC1FXWHnS+u+sPrsqUIBZBSukYf/kKGj90LcgkZo6xxZ8Inoc3wP8
wlmd+OyJOhmlsLrQMVWnUIdaiRoQRvDPmrqNn1gOeAvjxlWDc2IxRnwXQhv/Km0msYjCLnxrvZnA
iKGhVEJlucMzeB11Bgll4G2NTnCbVP6S0FOp6jx/6Npfc+2aBXMjetkrweK2aH3JFUtLUIGAQBDW
WG1jvys6oeDLjaIfGHhq1142tYnKPAcrMcjrdTI3dG/6javklSzyMaAFvryyWJNDFvS1A3zzwR8H
Vf/pqI3xneqqjsrtSo41vYgApYTKhOFYLTGaU5GwIuaYRm7uikEKHtmfhiJrB0pYcmHs0EzHXAd7
dKEl4xaWlzw/s+azdYmsTa96DqvwZFwHgkB/NmqlwoDOLjwN0ECVqnK53pBQ0QP+d5nRxoJ///tY
+zW903qgNHaK1g/QkyI4B2C91dUYq+c6BkR3jDHfgegPlHjHnpceCkHERLWD11F6B8sJpUAE9owH
QxrDpBzRYCKvkltHvGbxJXdo4F1G4LjT0OVM18AiAvaCCjvWTQ2h5VXskBhjmRXHYkvSYBznJw7q
kRZC1b5q9t1sEZpUOr1QnJCTQopfkhE/lZVgYTWSsubn+aICYJJ09aUNPiTaoDeyiTX/sX9YmtH3
4NzowXvikduEXC7RiWd1FEe2aCETppZKaRGu7r6zGSU1eZmME88bZbmqR41Uf7f0fBUBncOeZosJ
pqMT41UGNmMmXK0plLYOHlvsYcFmU6C16v6D/k8bTfVuweXy2pIiXPiO/D9hAT252RQUh1wAPQsU
AQrVwBtEkeMl3LEVRniEwg1APooTvr6XdpeFwvR1ycYpC2OnfArrH97WIkTQj5kDoaC9/HhWEemT
PsT/k1nR/Ras4fAngsbebiKy6ZeexCmiuPcu37CzomVCIUL5jK0egTz8ouCGWxyw0r8u8FMT49C+
RiIsobyJzx+QCkXjxcH1mT70KaYO3itiEA0dbV1e98S/R+VEUBlv6XhIvL4DZRrCjb8zSU/feyGx
iQOqQn6nXkPtaMz7KV6cybwtmN59sUoK4iuw9hRHtXD0FPJizS+H5LB8yCz5MKoEEydS1k+gkt/g
ZNvah+KpkwH27Ry5BznQKRwzrsnfPv1zXt7VsVyp605fO4jBJawi1ZNmPfu/0V5ZNJWfCvYXKfvQ
5d5+2zGhnCn7ENlrt5OHHZ71Kh9U7nGf9+kLWdEiyAhYcPLxMLBce4J7gzqsJ/34x7ZFLU5+RFTn
NKNz7snMq3CbC0CUwJ+xx6/7g6Y85NFAkfn//9kr0BE8Wpe5XKUce7zShRwfzkAARDtROZRuyIbf
SfOPFPL6SRleRmoIlAim7K9OS9L22ewczb0nq18U1oxMnKPktHSdpPTQQjC9y5SX4G79DNaV3eZN
1bjQK29NPueR3FhYum8R0AC+TxREXLDWbrVjwJ9jZvQ3Z+6rLuZhmshiAjcxf/0X0bTUwo5TGrwD
xhBh0VbVq3tEAOLEKC44ccv8nSuph1gj29q/w+LCBVsyIu1BEpwHjvhUhg2Bc0ztPuVzdBFv2PSX
vKMjf5qVA45hXzkzBO4nb9PLBgH3+HRozdUyoQaMbAaxLTxnsAfeN1/9LL4bfP+C0i8t1qUdf6kC
gm4wT0cZbVuY2Jm4QkN8eFW3nJTla5YQCqZMY88cv7fD80rAMcJBJrY3iSoN2B8khpFsDrLZvTGx
H67BElsi853xeuWRHsJBNfFZuOCNn5aUunORf1dd1yHdjLgGmAS3kG0p6sjxfs5MdFsTlIiLJWC6
h0OB/GqDSEU/Ikjk6Wr4tEkvM/WKc94WuAPyq54R7ZLRYdaqoS89tvX43ITxuLwQjfOfxS5LFrZw
/vBydke5NWm67UcBl7Ox1T0WNV1lHryOQ5mLO+mVtjMEiP/+NK9cW+ROsggkKqoCE1TVtyHdaPRK
PoknduiqCKo8u3Joa5wJQ9DuoWGcsiAIR/0ShqhPt7rpCJoWkY87NevuDxqGINYhsst/XXnXxUpa
hJzeGuAHpnw3+J4kKtzM40alnLFfxAp4PZONxa1PR6qTOhc2wUgSXIPoQ2fwXWxikKQuhGomnJh2
Mm/pdPG0dVMDFRfl6NQ8ePMyU9YlpcXLgKxLbt4oFc5RT4yQun4yN8lEZtdrIr7t+8C8febTzbnn
uICdoqiMgRj62hsinSWTb6Dj6dorTK62oKPWo0wuPUx6sWkFQ6yE+ClamH3y/wbW6fDVx/8T5+gR
Ws2c9wuWsf4P1ux/SeX1CDweVpuKILZgtDVTR3+PB8sYF4eljyMHvVg21GVkDFJVoSeBu7W+t0RQ
It0m2sZiQjN7vZj9XwOfTKHY6/iJNn0O6xobUw8ObsxJA/NKFyAuwclivW75i6dt6yAbT9I0kQTQ
XtXnwn3bfj8/J8QiVPCey09lELOy9YOaqK/HaL0QDdx00+fCGLUXgTWSDcAc+ExymEoNYC4JvsHV
uBzsQkKpq3uJKsgGvK2t5FFTJ92ACJsWYZ0ZGMz4PibXASZhPLBQKcX5J2bP7hN2jEjzeNG9872x
JdmLBU5KFO7pQ5SogoiA19iKSs/1CShOR99NguYRJ2kfCOHmun+XWF31Ew4qjAaIG+8aAdFGubhH
RROiAzZoIHVv/JbmPOcenXf3mmF2ltkKKRwUjKWg4vJXq1fgsNWQNliQL/aHLcCHiAg26NkikI7T
tGxaCa3yNMLB3CDy8aWckOdmfmIZ6RaVKS1brxiqvJc/PGZT/BnCbBdI6+1o4fRZeiXgDaZoKoAt
2dnn5JnQl/5mWO+YIuN6Bo6mTQbBkyC1JPiaVtiTbSU3KGR/sZMZW4lgBRkT4VBvESdW6+zPiz8R
h3dSvbmfNqmK3R5Twj0/JTIXCr9/lT++ZDiN6sgdacsJ0eoxQaj1cYUdyh/FeBTuiP+99g0hpi5W
tmD8O39mn1nvzdArUtbGGrZM9pENn/QRYF7dABcOO+FS/XeZdCaRPvMzEO+J1T2Cu1bB8hmldyJR
Kr1ZmlXudejoNaWHZCbWMe5tz6ZOHVAthigUU4ABrhNqBoQrUlx2/fSYGya8Zb8qrr9YZn9U2Rw/
Zx9pPpO2fOAEnUN6Ql6b4rjTFoZad5U/Yh3COix3RHg2QTMNb3XjRr/OdCUpD3M4OMHM6dlCB9ij
QBwM0sxtjAKJhhjGYEKYQXz2ugCfQOij9BzVTdRb4oSFvT+b8v5WRN1476MCpTv6jHdrCyGQpWqr
ktgz+T+pwG7bgMcx2Sdno5wXgLq2/Zj5aqKweYAjm5wxurpU3w5MuR9vkpLmaH/y9y0DTM7GFgux
5JKpodbXyeAUDcuRo9gr4C/XdXD2Dqs6+2qECCt9sJvH7ko6nK/cQWe8HmlmlXArfXThPOSMVvUE
Ih0VmNQ2caUYsakubLnuSfyviC7sO/w5zh4Sb2FJZp+tkBPJzSBVxNGWjU7PWI+6WCpdofhP3bG+
BWrMXj022K3ldaLmXscNQV2z5yvHfHeB8n2jIKZWbx3WRtmfpTqzWEhEKBcjw34HtLtTcsunFBsv
NGbYIX+xB3W370+AgKHngIKnaWaeMzRRDY3xl8OB680HCyIrJAnA8eA5/Lfh0QOhm56kegj0Wd8o
p61YUn3lXFCv04cFJc1Zb/wGAiJqb6rEw6q6PX9+zq9/+TQUdJTODPUUEEhBXLDFNpHuiosW+VSI
qFunO3GEWd3BnOTiQPxdpzY6r0JAUwVTYIbpeMp6RVWr5NvF6eaWsjrl9IyQ/MRya88DBe1TkwyG
jsAA29bw17AHBdOTF/VCSr5aO6ECefzUJvK8+UnLMBPQk/ZPTI7UMyXH5uw/jICXsO3dXD47NFd1
IrCInQkecTk8PdwHpw2/qvlWxeI/WsqpRuz6TiEoNMMN3BCZaC2l+Bbt55ZuWOJeKUTCDSQI+DaS
LCXBbWsYQFZajICP1OOen42iVKokul+WnpdQdzivj90CRsPO/AcI7o29FWIdW6ZlfvK+wivXTqP6
O1h/qThe43jaP0RkOze56HLGDa3Hu/otGyz+97XYDX2i7mBMtgSD/garTCbWZjburMcsyhHFL/VO
G/ui5q0VcizW6WSSreEQQLlsTmXDgVN0o71K8COdcuFK0TolFKefOoBqZGC1sJhns8Rz6jeyMa+C
zLXdoqOr1OQdS4LT8Mv9tGp1G5Ir5Rh5a/gLcCxQy2orG+9mRMeQxtZIK0mujBkY8v098lVbe6Dp
pNPfO6gl02iHaQob1LPfqdv9tdWm6thW54cFS/x34G++4Sb5MYid4i/dbGLNCXOr8sNhoDXU0uAu
ZFTkDuHAxjY7+2FFme8Jb/lbrtmcXZzHp8iSFgMJShfDK3uLtcL2PnzuhVjUGUhqeLi3mZmn905s
zWRLEy3khJwEK7vFkJ7cy0a77IRCymt9I3hZb2Psh2MGswKCYAiBtvy4dFFrmzT0b1u61Q6jBJUe
BAFyAmfUM4EwPwT2LUQ6KoAeDqq5pGRBGCzR9ocUfxVTzFtgavuuzkrkSk4X0oWBPoPWkZM4oo5+
gBtcx9e+enCHFKycw+Y3OJYqrtc1piZYaWoyKZbsXhIdeqWmxT0aKTIfE3U/H3nG18SH7T2i4wK2
bMBS9nOWAWQqW/UPgGHBWRjoJz7TRiwbYKgJcC0tiyjxPY2qRAXCEbgD6v8p504hxiUOCOo/ILP/
3csIv328KkAhNyQnwGKM3emRLCe9gIL/KpbLBqeQE7zETTvx0SnOIhes821GiVFkyokBipNphAEP
RPIp7iuuAAgEgtt0Po+ur58jllUTnIEPXgRH+ZH1k87Inu7v0maKZsp0o1VAI4Mbouq2eptzqgdH
mop09jxF9OTTEAhyz3bDJmGOhQyUQQK44ZK/P/4+mP4wpfS3gEaU61C/T5Mvgg+xeKSXmhm2LOg6
I5XygxjgmW9adkqDwjS7xweM5Q32rDMza0IPzJMmvYWbVswHeVadfotKOcOPpEe+BNJKb9TX0IHy
f17ZiXnfNgwXD2ALb0nbJwuZ53ioznR9uuU9uvorMUeDzLtnr/F1iOh2eHmZNSa6Xb0SorR/j3wx
LNaJBzG1SK08XPSGuq/+3zOS7HNR74OR1vHMt1DUoodrRUJaIzGvFOVm9eqI9gcXHY1Oc6+eEGfx
sv/VKL6FoJMFVLLgX71xVntEi3CvjggVDUhWjZSic8oNEJJeJAj23KKGUm+lcPWUlcowhL4/aPFx
JSpCif2gcVs02MTLW8xvE21KM+KgAlqjsuOpl8fCGHY0wumqE6wYJOpca4Z2xr37GcMKG/tGXGM2
JTjldxr4whAlw5k+r89wHcjActf3d/8PPfcQrEZ7RLE+2ZisemZ0XixIEICBik3hJW7PvAxYSiit
FVtCqoUz8alr766WDjn14oMbpcEnpLOMBD48EoGVosaCvfewbZ0NqD2JjhS1/uqKLJZ2to1NLNmh
EADDIhCAM5B+LHHXNBWyHMh5fgd+gvfDuBCGA36G+X+hlgTjX2JvEr6gYFoq+YadT6p35q9TfCb7
2M+IZ+UPGr7AlbAJpmhcncE9J2Mi+W1Jby/5II7KMaqSnAWuob8sZwfkv13ixLtDMKtS6dCSskcy
/OOpN/Ta89OkKiHWa7uSllJK8nefNqNq3F5V0N2FPFdMvtFScJPDr4BYszZaQgpvpxYnS6329CA4
V948LI1gKQ4yofms5ZWyha+KisbKxr+z9S0zaXC/KEq2rJ+nb3ONOMF22GEzfyx5k4M7IgS7EiMp
DSsGu2OBiNeaBfx9QcX7h+x8rmRVR+cYsiEkkCd+taDF03ZtvgRbr+ORgur4TyiJWdoDtZ7xNqQ+
T17Ht26x6SKeihp+LIboh/YMtVyw8ZXOwmg9CqTKTzMlbyDqu+WreT8Frvj2Qxj3+r9x95JassOR
6FKEQDFoBOKwR7MYAgWtkfPWEByCDPbV0gUyoHI/Ow+moDkGV9HgPHAerjKRQ/NJw367EkplbY5W
+8HW1vpoagHxYS33X4ILbIi+xNIGnMwxkK01Qz7EImQT1n0tiELLAwO5DBuo3weIkoQP5FpokDzs
LikaF88UWGA58/+2lYsFtCEk1stSiVXy3NAqv47r8RrloZIunkUs7jhCCptgKq0B5q4uNhYTDNm+
2Xb3cryE7fd38OSOsoNsaz97KHE2qnzfFCz3ytKpQMyAAld6FrjBlR3Q+mXlU5aYLCCk0xnbGYaj
4Dyp9DhxziclXfkPrHMgyUW3NOVUO/K2uOMd7VbRYZJ7VkjljChAPC66ORUEBv1E58imkNFXcRpc
Vs557TOfF6NVmXtzXGB07zmqADvFRw98fOjokKVRZaPPjTDjzidNUShEYRe55xlhRh3GERFWLL3V
Z0GtCiIg/artcK/isg5NVqbqH2FSCiQQxSpxrs8A2JnokDfD+FVzA2Wt/RAUAmA2a3xDkRYnJvpa
/b73tHwPI/v3WJq2lsmcfEYNT6wBxiDopn+mRm3RXKqNCQVPZr8roLHp1sO4JmRtdkFRgtv3azfq
btcc4ySIuQjKvi8gc3WtoVmAAvxbWMViZTzuqws8H/bN2LgVIkeyGVnNUmnXjELzoqMC6fPgiijt
CocURcf7TPx3MNxRW9q6iKCgsrwZKfPC4NkWbmw5fcVzP6QZ2IJb3DRbsUevPgu++I5ntA6yHsG1
25AEZUKOkewM+7lRXTo8dZQzNh9NjMlIkw9keUdlG+WVY1l9PyopxGUDF7HaViEaKT6DphFVayP4
8Ou+HomyyvGn4U0ORAkPyr3G2IoKVnrDVlqDkNvnFsskiFDATs04tQnD1nHo87sQmXOL6EgUQVQl
CjkZIbRj40+F8MLQ634aQrZnnLUv87o9ix3xrcs8AZKHxR4MaiG52FRsQV7IlOFQcruO1QqZWJY0
mIA41XL9gt0PsK4sm8wgvVIjFd9198x67dEonaWeUAAcJes+1+PttjLnZbXPIak7nPLsq57S2cgB
uf5r2KMyaDYqgxx8WPpDcedc1pB9HhhCPOoxTlbe15Pt0YAM3zAFfOYTH84zpRIvoAaN10jgTt2P
v4xsHJv7xc+ipn7KY2x/kYvntR5yW5/dTHdyh4hpHTcwKrjG1aq6lAOFzAanv3Tk63hQMa5rsv4L
sj64cmvDf9n3VDUCaO0B4VIV7jKy54r4cfh3Xm6k6LGi/CDfMZXuhR4P4ACTEvg3rdg3/XzJwQNY
BJM6h7dlA+w4PiMCYHIUuNzbC18W5U2OmATk26z+LhGoSSMy9WMsq+2hJqRs+aiJr0xd4mhsOlkz
1TvSruFCXX+pXZvWqDywe2He7z9qPOMslmHWRBFLHMKehY0qZm7XgY9WMYJKJyC6deHOLCl3op0V
pIszYZSU5ugH9xCn3CVDcPywamYWRlG1I3NC9LYGqF8nwEi5GQexYqfAkE9cZgThTHLm9ayLYjVt
9qla+qpuoOJatKyS6DdzPrKXEZ0BPo8P+Z8b0XgI3ldGUA6Op+U4LOgYH/iyxwGzpR+1rVza76qb
HTO/PsTfxwwSDAsnglYBk3AiN/REXf7Rpm1FJpEIvdRGPSIT49FJURFj9NgQK9uMDnXArQVKgI9z
BY1USMRWRhJxc/rfm5N58AeHPa8vIdPYH5PYJ+rufdugeRDP2AII1q7i4ii1yHEIi+rDrE0P2SbX
7cBMHYBwwel9/12/p50mep9488CRQKkDMUasJFAf5iVrJPyHJGtNkIfO2kSrGtD3jQsoRhnD3LI0
qc9P5/w6NJC+SVglJH7GJ8HzQGjnTRx0RyKec75EVq3WYS1kk0AtXKaNSe5RvSh1nNWnye68gGFC
n5K+Vq1DFNZzt7DZttPSUWaa2iKV4f1dOVTFbMUwiPw1jKVs3ciK8ikdWlLN2yzFdZHwSZY9Lpn3
9KtJsp+wWWA7N+ZZE3Ko9hKFw/Obw+JmEAFs0BDyuZyQ+wXnidpwUJiRvOGlxEDPCxFyBBL2Z5uR
e9s/+5xgE/sbbdZDWfuehvsOaJa79Wp/DP2Yb9Ca1MtvwUvs+epjLJfcE1RDmJqsoITux7GUf51K
eVoEHoh7Bf5KWaXNVclDgWFG/yb7SywKwbKehG957hDFQZ5vMNtmTY8MbzUqToHIMwjQxKAH4qW2
Rsk9jwJ9WZ78WLbyFGmrANrzEB/2mJ9vjowWtLzItv8uGdwybAJRiyurZL6tfDMVxEok7/bGDC0B
pbnVrNYjXFlXNRC2GUKpTKANowIofvc9yNCeJel4VquPoYY4uEdEglX34kqJuffu/2UEu6mh831J
U093Feir6vV/AObMmBhipv+2L4ndGkfvYw8MVW2DOYcN8rM66Kt1hMUAaHyItSgIFy87de6p2+YI
HU1x4RZNEfxUGak47Ke/Lw9pu8D/xwQhk2fIvvDvoARUWAUEcjvgP7ZbqPuAcUyUloo2JKl59/UE
A04pFtSjJtbarwN282fqJqJDHWwSjDqakXSkgiyjB5inQlXFk9zC+w8rOplwHP4WL/8N12H56PmF
6bNMTB8cgSJXTKXayqvEeJDCrMOHcQtXeSOL8X62VWLM5VEnKEa3NF3axSm39uxluzY7Fo+McMS9
BqPYW+Y0/xAUtfjirCFAP4Y1gI86aXauStiWXoQHBYfc76CVB3Kz9GFZAwy7OlPcx9I0LnoVTKGh
MqVYdtBpXnNRyq57GPDOHcFSJZN4YjtegBGuEFxhP3WzIke9TVTpVcySKUh5D2agfxNbbBExU+xQ
DsFjAAbS2E+s983gfsYXLIr6w8VcyThuf7e7KK4AH6OLZ0MTbT8ZnarHy3jQJHDBVzinEpXeg3tz
NQZAzrE6uREJZYiPMLilxvXQGptxJtLeWVPHiDDSfMRUuzCJ0VuebznIyGWeNAfoSnGNZ7l3Cw3V
ccJA2Zw69idVJLHH7niHz23n2oIaM93L82ALbv35kT4xZ995yoHk0XfUtn2WnpZdzef0F71M/Ih2
Dm4WPJuuiMj6l6LNNy0+tMmXnXCgiwj6NHzGlbO5pJvTCF3lW/GA4sLWeQKJnEyqicdpUWuTIoc+
+7WhdDhGAHoI6FUkUMy2m4ZJp0x51r10Moxv7zvqTlp5Gl+PcFJybD8UaME8SstHBJVi/082UAhl
7CplvMWCUiQb59CMcMT9R7KWNUELScdqbes4kSpZsQcqF05yhR3xdW0D3odNEDV3xvDWC2lwLK4V
iXs9BgfVo3/z58JtIL6QgEV9PTWbXvG5LPuatdKRzuNIna/AMKksHIhCu98L0es3/cFOly/X0Kbm
QQWajJDLG+v1vrEJF40cEpqAahF/bhaCDl9tDgIDhcO2oNL3a8/mW4XLYL1oNDWcT5NADotq2jux
7UxO1Reyv19YlGh31zrQlq+tMvMUROsl/NOvgeU9GJEMQF9b7WLTk8U7fOt58+JvcTankY4ekN6L
hNmY8ZDan1A+mBzu7BWty336ilm9HzqMF7w4VuGR8bHUN/tOCKAcW9kP4m3vw+pHs24lfKesMTz/
y3eefaAnRqmjaOhotrKOlJ9smoFFdJP37uvXJpaN4awr9BrKyIGMrz2vy4zuPfIVjophtY7lVdCj
ggm8sOfvrz6l8TymSpn2ytzh8QMtoM8X10fDso69kngGBf9xo7oXKgZRGJyggMCXulHAaQ+a5q+B
iZToqwxtmzQhm5Zd97aRtB8hqA7AgKgIyawU8k+Z4QGHf5KZZafmlpQH2r9+rxXoL4Lgz4gEEsEp
Cp00AuuxmRLUEU0ahUkJrrtnkSAssrQT0c0q23CAgkqmSg5pml9xzv4AUtHLRKTw9ewuZC9Z5PS9
IIbW0PLViRjLz9HKwc+iBWUnZa71Jm/Ha5ha/dO0pwNmDBW4V7iUGihLkd8mT/7dbOV7BKrl6qdD
saF9q5ws25ZruSKIge5yFzEw4bXH5kEQUVilvo/uHeySxW1IzC+JongwxW2PAu4a6AyVuTBI/Tpe
dj0ATPr9k36wRXt00SGPLlNBqo1mIGAcD8p44xM/7kVWGQNE8rPUdxQzijHVsNEtfNbRh8osY+fD
98hSIRq3/GAziN/19ZAud06jiFfkRdR+2Wjev+nk/0Mlz7y+zA/0RU8R0Svc6AkQawhD/jG4ykRM
sDexonemV/ZbePbpHTqYb3Kt9RbLHSboIK4jddm9weH8iSa2hhVerIUajUqWWaOsRG65Ss2OfLql
Ctyp0J0KhTCWEfJnIZYi5VDlM06+5YLnzYcrxAmFpP2BGKNwUM0JCpUpO2nDdvx0u/h4tez3qfdm
vzYChd/96oMJK/dZuWNh/xVVzC+KFCQg7pl/nBo5o1vaWm35hvcOvHLjHZX+RmmHTmWqqCQ9ng0m
j+7llAB+0VIoaRLR1KTmX/3dNP1PDspn7yk5bkI4LNW13qwlLVnW4gS7+bqrf2Ndpa5py5HUKMb1
X2hrhX294APIPHyB4gjQIcG+MyCwEr6ZTYfkHWxi0S2LSP7a7ZuAAtdAAXxjHa6BO6tQMslqgto1
u9lhrPekARCoeuLBpbMcTwSMxTLdfbxQsIfkzDBwyvLqqVzeqObPRLKNWNT7z1R/JE3JslyDeC5w
Qsv8xJLN+jUOcVY9SjFRPl1SxvNlKD+j6GBSw7RdB4vAU+SVljSqxk2BUxz+CUVWqM3usJo94qvq
myjNnAwGwbLDhsJLEfnLjpRrbEuCROmcmRCdzyyGCfFeCKtOa+glcOaiNO7EVzv08VsQXM4iwSPP
MO8kF/dBZCky3faZ2qQWPxXdyzNDy9/Bp/f9dE1LAmENELaMqEJhvp2RedZieX9HzAL2fc4FJ0+d
2G1YUf1hz0Yg1sBtkEDNYXseYRIBIQV8ftgM5K/oE+FvHhXQ/5UgjM5DX0XVSf1L5LzJ4DjLPCNx
j6eeBP3qkGNh+FXb0hiEoWGTipU+0nakUeOeIwzfgNCXoUvXqLVKPADLEehLmucoR02UtPBFI4Qh
3frlTuTsn+CHFarEgE7p/PNmDXfK2fGtmvJYYbfXeLG9xC5GPMnU1jl2lNRuADyjtfyqraOGh1Xl
wvx5hKuteHICpj0LrjZ+nucHyMhVS3QhXZc9h0LS8tlaJh/YNbMoTDgWE4N3JS9IpvCPv/v8WC/V
caHrCiiymugLxHIzkTyW7l5BYK2AgYV4UvSdfAZwXgLsN5meJW/AXkWq6yXehc1cRDESAAuo/9uf
XDi7ClhkcASqqSIrQnLnUSxAd8m7MUvoqzQ9dfey/m1IudJ8SrGaLF9I4OU9FgYRveF/kKJTP1yk
e9DwJBsY+rDt6d0s/R9xo1vJQRQX7zZAxKQtXNfYqHU1ZXwpa7LX7jn0POKRxb9MH6m88XW0adA6
+PeNwpeXPYU2Bq0QEzXUYJ4qqP6l+POecEbSVrYg4IxWItey2vwUQaJwEFv5k3R2OVYjsQ2IOOM3
6nXRu3PpA18zcb+VG34DawZ5K+GK9GS9YfDCwHGfFU/G4pD77mP1Yvv8UiB173rhOxwEpV8jt/lQ
aRhJ0MFCxFDw36GIvpL2m4QlDxjF1AWOdKpw5NXeKQTRXTSYApOzrPE8jUm4CkFMEaD9CKldHMzH
oG5Nh2FocU3/JFdNf+68DiuYiib4MlEQbo4JNIMx3KO3aPplP1giLjOtuXNY3JNGfjW5nre6J6FR
atfwwShxzQoRdP8c+jUS/9awASgdjK1paq6K0aoswqmWd/REBtatlphRntrvv4WVZDRMEGrI8EYL
lxxS7AEGyExecWCBcWylU01vJksF/NaoCsJ2tkXMThEXGBBba/yVFf+hH00DbwmWYUe1so4g95ip
rAlr0DuELEKHFvRVDvd8lJ0RISNjRtH5q1up2ioGZDag7tkGAtDXk5V0EhsGpI49TFrHgoyOOlEy
Kv7TJKrnT+3eUW53anxEYZPb4OxIMb8gVzL+pQpJjVzqs+yyBTMF0w8BVNF/LSYyLTdWWmzOiPm+
kQaED8sxc0s/bklsCzCJe6TXzy2dJtQEhLTD+c0rHG/AVHQt4MjOmodK9tr2T9PfwGhdxsWSBWOR
VytIMS/mc4gtavPM4cz+hkBDDgmvJWVr+oG5hkUPVaKiwBvoeEGLHb1xUqbcNv+Cu1PzM2eG0iWN
X7DV2b9ayGB54jbY1w76i/ovcC2R7gm4FZ8z993XFcmGlMNCpUDU4v2+Fye1aOLR2iAX36MTItKm
EcSFOglOxjnWGY6nKz9Ad4zb5fIUY+iS2CeSzWxQODnHPYfHpcySbfRYAC0FO08v7hDgPr/fUQP4
VXIbgF8XD5K6LHlHTO/HEVckTBTtJyDbC9M9HraUiJ8vW10yq1U8w7kx0fbjet9PQ14Pp1nND7nT
JHC4wsVc4I+1gUxHuCEicfxgMT5XTCQtwsyhddVzKGnIr6LyreXNp0xOiuVJI8A/MB9TMoG26CUV
JwLPSjQaPBz+dkRn/hiq4NP1rvknXpRPUcbpjJalOU90XyMVjJPf43Qdhqy8ntRHT5aLZbaWzL1u
RB2SKCBCD1xppcExY2bZprEeU5Wk/viB+jKNFeVx3cCCWH+T8aIgiVFQTau5V4ZwqTfZ8mOwXqFm
5sF7WtXlzdItmcEUPJFXOs4IPoIfFFlKheKm6JrfzOTRr11TtObuJB5BKmIkgE5DucYqFePuCEKd
Az4qMGBNLDpW7IAsTCMCdFfMls1XnJ0FCQTvrKT/noz+91AoyPNpPe1RfnHR97Vu9+6vbbYd+RL7
Cjlt0DK43LPKoBs/dmooSeRhASeBsMHhB3LHM4LglGAPNU8WAyIhb+kXN7z97Xc9CWhcRLqVbiDD
8wQA1NSIVqSjK/RZ5iGvYnCVMf3vP5ZMuSc7HH5bnuSTaF9XzGlkgE2uoYg+Vy1xZp+0i2IoJZXP
X6f1jNa8xq/3hvkhSe9xmoKMSiSgqfQhONA2PCaJ19oTHXW3Xd9FJMSEF9OMW5ehZWl5E2g4SSvO
ra1fL7NipYXXoOuD5+98peFe76G8oipPdnxmPnwb5STWw+SkvohHU47L6O+9sAMU2MUj3F51bBk/
pEglMGFban3Lu3WDzBl3+bcTCKIsQkXKbg/F+FmMnktLv/22UMdXQZglJpd8jnupOozulD7/T9by
WZT8POlOqP4u8SwioIo+MkSo+geVKbLE8eViz251fTe4nyi4MTJWgzZkh56+FB04yCyp209sZJHK
2la/6BKXbgIZbJI/C+WlyJZ5031owdIl48LTnYguwMQZAyp19uSG2bqISdSoSdUT2/SuVMRNMnxv
neQ+hFnrN4R0sAspE69Po161lJRx4nJAfQGyZcyqAUlMPm7myuL9iGE09OHCKPkrMKQ5DoWXbh33
i7QHX6eChUSy7yLjUvLJECSOlMb6ZsCpt1VsJ5+bgbu+Na1PvQG1cEl6lL/dIfR5fdcPjQxGEdPS
xKvnx619mKqsKPIMvi1UD8o5GmS+c1OGJ8d1qLT/cYxgRAgmoeso6GFm7argtSixdLxV8LL5mSj0
TXLFKlGbxcVXRBSjXjbhq76dInxlOw8PHeW/ohetARnzxrBq+WQCxolMn+YQCk3tvze5wu565a8t
WRDbkCW9VRF5FxRdpqiYqI4A6GiBnXV22dHTPjU93G3t+neWT+4Gsr7dGrRy8lyvf+CTMoUeeBZD
wh/8ZiMjJV4QHqObw8BRrjClf2c8EUVlgpba71yomA8KLuWlJPxUY1MbRRcp1AVHD0Mwq/SvTplT
9XXihYnd69ywEaUH36Z2bazdYotloXMW9DoYiCrRSlMoD4hIyLksCgZFqhjyNDwjsccN90D38Rsu
mISe4KbZKJC9JtKIp8KfHa/cfDwhH7CM9kGj5hidiZMI00HggljxzEJjqtAWDQYgxrCmi+8wlThA
tmyyYMmbAvVfAP5cLVcjQdMx2839voY3rPFJNrPbPdt03OlyZ7IP9LSHUt7nkQf//VITSXwjK9QH
g8DrJZ8yxQwk/ZoU4mOmt2xBpyLxG3V2of5ORpiLRUtNbW8MNuIzjvQxfmU4T4eQV9benjg7ZWVR
H/NeKCrmDDYEtgA7DYJG3NZsuiWXpEzOos79V08VWeLwAPh6t/ykEaEvQFupqOeKUKlWWT3IQfFp
dLbm8L4UFWHoP5/tr1S8ojJdjrrJXGJOJie1sp0K89oEDT7XyHl6qXD/IY1Ma1Fc46F4at12XwkQ
xTfKu6DREBS7mFw/2RY21MghzXSSz0eJck9l26Gof76RRAXt4bQGHXQuzst8pmRUi1h63hm7JE6x
zLNRsa605r/bpsplFl+b4CQA9r4aZmhsw8Psmn1cIyZ4I3Cx/gtwP6rpC1faP2GC84ejDSdhRZTm
D+XLklCxtoHZIdqohN/Eue5v3G8+rWqarOuCW+Jf+q9U+OIvRNvuCnYqy3hSWRjGFJNpg4aAZqQN
TjzW8Bk5TkaxxdlZBQtpc8/D/RX90Lzd6Xp7ipxdl9u4MLPqck4xTpM5r+5+SP/L6peMHC0N7pIk
XyVdVgUirRT0EpvhIy4kJlYm5dBTfqLRww00vtrsH13pgQCyM+7hBcv8Qf7oY4H2qXzZDDD3HXXs
ZkmRBa3czvJzy0+VDS7WV54GVCUzuE5ilztox9nw3QQWw/yVRigbPU5P2rx2aNhfWlCdAEW5Jjek
DjQyNnk44RgFiiYUPHi2/8SYG1ly+uVN3gUmD4bbcuaG2GfbIrg8/fmHyuyRZWRoNFl5E0WPk1lI
hortxXFgVVDHXa03fyik6II6vhI2A9lW4ZwNWqeBIUpK1CfOgFbnbDL8majxXxu3UkBFA6b3pn6d
g2E8GPf3hYbRyHRbCK6ZFXFK5jP9CKBT+0F32pyrRekUrX3LsI9fAdQifJ+H1kdMxw8cOzR197vr
IEFr3hAp04pTX3+h/AgRXWqA8tpNWxbk8mKQji7m7HdA6k262ZjGBnjOdcc4Ti1+tGsJotWjYU2p
3KLHEyvhi9g+l+jgysX3lkE4Ak0AWO68pfXFgKq/BcM8+phJIr6PSKYlyLswQb+hrqRS1aUFJsOL
x7oiH4B+gRE/3QsfHDVOcDjLHfRouDy+16e454igZgzUwogXfG0KW7mDZ9ov+UxdcnRDVpnxW4T1
COJE+2uWN/LthJ+ziilf/GhltIXV1wqSpLb/pm8laHOEl8vK1GsIiFE1sEP82dpuqOZZYIJBKlNM
RzdRPXncIVxhPXhh7684UPecYl2idk54uIDDN8drQegonpnSQ/lddhoR4PPvz9kW1nB8ehrjm2D/
7CtYg7GXBUhhnvwGrSyK8dXBHicDuA5tAP/dRIEPGij0WlOK+9JTnNs+1UJkNIpDcnLkwOzco45D
UhoMGDIcrj9EXZJ51RgZNHNR2q/bWRBSSDRtsy8H2th2F0uj5v0Iv7h9N2pBIUrlhu2SrS0I8DX4
REO7zbsLnwrs+AmRof1EeX1RPyxlhQg4zrfLO27Jcn0c1Ey0VX4cKax3K/HmnXqRXeATkGgYjlNj
6zuDeWuUByIcK0FgqugOk7Xw8Bwd15VRvONSmkzToAC/efyygJ96IEu/UZp/0Py4WO3sX2d6es5N
ixNczg55WLQHMOuoDXGPW0ydj7LlxDMSaI0qc/ELlEt/oLHMjZc+336h/2GSu7xobBxJqZnH2Pxr
Vmimyz+n2UvOitd5Oa9kxlw7h0+ulqSH6zl6amiERAbSSi4tqvdT86dFNCwRGNl65nZez2mY7orj
5bOFUmvwLNp+jAEMjK8JsErcVwOrNXO4+oMZRSMX3CPxq40qWGXcnoeUkIZ/4R0Yd62trcSIQu8E
25/g1q+99k2RD+G0GvnlMtB/DHpUqfWGcTvl3FYmVYuWNOV0GNOZa9cWF6hcnfMAhKQT7l/xs+Dr
vOPDX5z9/ffQYiRHEGGPNrWcqNjQi6Ax9VsAqjxXjngbzPS9+HUy5KBIkXKhZTp3X7AZVbQB1vtW
TfcZz9TXtQQ6WLo170DnOIe6aoCInu623MW7xnRWh+gW9sdfPGoSXCHnpehWqn8KpcQoLgJKUS6U
IuTslaf0sYnbNMlJNdbrq4MG4+KZhmphP4EptIr05MLCPbI894nqMQSb8cCBuh3AUJN/2yMzxZUK
Odm8ZK2aU/xgJQWg7gkbE7YT4IprgPAyo2bQA60OsIgZZsB0d0zDVZnr/OORXYnVRewRNzddfLAP
0GC0+zhdSsvGBaqnxlXM1xRpMalacnvIS5iJQIkja56PTBf/UrQgkm2ScWXQCRO/UnXMCNSQCH+k
v5oAjcQr1SPdNjJscnpGNbZIht9dpieZFZHX2xIpmhdvzur2kU1vAxJx+gNBtA5hlBKun8j6N/yK
h8LFsfyw6Q8sf5bqztRZJKYQpbUCR3/Q5fzxC8I+D4AMmof0mcvMiyFVUe95hNNeYK2Ic7nLPLVx
RkRigz7xwIMZgPZlhzGsrm3rJiB3n11VKiXmsj45aPp1Ld5QfVrt9TWXKBmli8ZvT8qWiMyXU5U5
kJ+tdWbCtcW08ySnLc5nNep94nLmBGvKSJ60iinLAZlqaCMD/KaWdt6sovSJx2s5ZONBOgRgDlZJ
WG+tp1+iSYrIxfy1HjntC/NvzsQ+kq6wrfvAdt3B5YsRpaDd2YAGEBLXdi9pvhAwaXDCllJTxr8m
wSdUNO1Pu94c3wS/Tr2qCrbgs736v0vvmxm/PxqrjKMJnFa1u/5FHYVEPBaYa2fpgwIEpNZTqfBY
+Z9f5IXD5UeFlDISQdcr0HPJAAAYRoK2IOS6wtqtvS7UuKid45oLUA67VdPg/+W2SXkey4Ggtkz7
i16aC/Er3Ph+59WcjofGic4xzP2MxK9TtyUC8pQpp3caZSUUDoh3JCS93W7IAbRH+kfgG7VYE8UW
aqrWFXAmlYZqlT2xPt7Vi2TwuVkWhlpb/O03rWyiBnArrqGXMkzrt+SPNgfYdG8UimfS7D8CGIy5
P2gR4BZYM1h8x3jF4UFwRHtAUw4Kc7dOTDGH1ri74xSSw+BZqY39nSruc4wSI2DUS0wxFwHsXAbC
mdc4aAKZGD0bMMw+f1eohSlnw5Sr6X3fgNshwNEyVXX4cmFTnv/+Oet1xioBQXSmgVXs6znRWbnd
KSPPD028Noy14EBmOqOrObacqGTIAAvqXwM8fWzPfNRtyiMzXILIh0Fe0+wNImaBRcblxKJ4Vzy6
/1IE6aZXx4v3xibRi7PnNjt9x+pK6rNccAIkCwp4JCG6gn9qCHAYpCHW3mFIccsY10jV6YTbrmjj
LYtimOvYSRw8wzhNVSr8JpvwSUhRAid2U0+4QykRVzrioWwmaJyFZb/sIAEXA/twNGK6wlK/pPfo
2IeG2ROdsEoPXk7PUf9cMkkhpHCWXG+/lbvqmU1YWXVUhSxNYvMSksbUQv0BI6nNadCBEMoOMDrp
2vOLGiahvtBXKfAEGBtnKxiUDX26Xld22Dnfng07SWowQ7h8TzwbCwDm7UmpUcJf/vSnmYtRxL5T
dKWGFHhGV5OWIF6jOZLqrRR01+JzV/KOlwXd7tXrmMGpjHjQ8oBlTWYqE2zAoAn5IbPQaTOB1x6s
zcVEiIP3tkfbl8PO8LZPPLzKDIX/Jdp8Je3uh8emAkqmk8uR3EGIRZfxLl90QmLfcVZN/NKtB5tx
bGHJq5Y+QRMobh4TrgCDsUwO+WOBMhKlJ4XFivPbXC8HhNtYBL7sWKTZN8J6ALTZMiRbxY/Y26zr
bHguB314wdOdeJHkZZPpjYOSpR33VmPjzyWU88FGZcrBzpdgktXMaiHll0J7Kfq6Pjjkd9dSHzVY
vyIuhJaQbbV2UzKfEOc9EYrSpKmLxR98S/k5TELGNQrn2snGHZugIuBIn3XvzTjkoINZx0OAu5Lv
gg5Oz8owQBYaNqQhhGbfCvb9in4Wtkyro9GodBOFnO8npT7RdpJXMs50KK5vnmiMnBiHBv2J3cP7
V6j/OoFoP+Hl5J9bzIyA+Sbum5LrmqV548nPRJExqtPu6cZAqVH2ESc+7UiD87YWgepC4YmiwVnI
Szj6AUcz2iukJE0ccfDIySC0iqKqObzi/+YMO5LhM8YL7AEx7lrJYZaSyr3K/lrpCxbgfLB+rFY8
Xug7xMZQdOamzzGTT+i+SUOUcpoXlTBEqYp071xQ+gtfWaPAMfw2sQgkjVf7T0Hjj5pS7sS4KJJA
/DpLlCLFpuO2EX3oOvJ8K7eq9g9he1t9WRDl/JAWZiAAFmyNATusHafbXgZGRU8fYqERJSLDeD17
JI7VHbf42lKrX1puzjEAOp44oSGYa8A3YoSclsnXpwEVmnJ5HcQ/kWr+WrxQ7IyMDevMdcnA1a2B
j8Rv6hxcnjM9PXIAs+RExCQI8GjC05GDypd93Cm5l6rUfPEiBZ9O+Kp5uZrrZRfwbPSpBBQn+YQz
rXYCf5jNSToMVgEV6K237W5c0+66zYF40K4hqKWzHm6GuKdm8y8MUEGPBz0VPTX1faqwWEsIi9A2
qpWU3x0OjB5/eX42DfZEEY6vifsevrENEnrRtpm8u6W0gkzh4QNVdLZeiwPZC+FF0MJV8Mdm+CTM
sXEfhIefpTv87kDNma4KZ4qyte6F5VX9RTGVYm6GwZTu4ldXMtrkV0pczSYu0XgaUSkE424WmKug
bpTnkDOxldzkpuLa5UFECg+lxiuCQmer0Fq40tD3+J6PikjZ0oRrRRMmrnZZiEYVyW9/Y0+Cr4ph
sL0onBN9FNw5Akqe521LJZb8MdR65O5qvzjnsm/kezrRxqSJkN4wGsRgMHmzUYbPDE+lOZFvhrfd
97nMfwC6w1+Owql2PJkKCz0HpzcTy1DXD6QTUtgyzvMCPXVITMWoW7agZUAF3pxItUz/RuWosNmC
sSL5OFnwJc7lXA0VJzXriXpdTvyBYUtljcOoAZjpC8j3fZebZUf+UPZ36lK1a7OHeivAkZqHxu5d
GHmTaKhJP+nQYtKjk90uuMwIC2hEUw5CTN5cdwarXM1PK4cRvc8PBDyYxvA/WbAhcgXSa8aldFwY
0RA8osnLKg8HmOf64x8W+j4Irq5YV192pne8Za27Z2/Qt268HKcB3x6V2M0nyyzTh5O4syfsUywh
kWxwtsUKQ5MxmD6Jea/4vffSrJktmo8Xf9p/VJ9inQ/QJtTysLsF+N+/e2PORO5y42fqxYUIpxfs
Uawj/NQpx014THj6EigoVsbUkGaknsBagYTrTW02c3qyUpH+k3dowav+XLVcUNgDmjOTL5Qn9rFL
7/ZwRujAsS/jGFtHb1xzCa5TxB66osfKZoLnR2X2ZzeI5rI0hOgP7AY3Q40dkRlMGNzfxCk09VUA
KU1wy+hWqqVZe8Zn/1DCbArq4BUChQa6PgFq25aHrYPY3KpCbMdqZDBCL3Bzv42U7bvb2oX88W9q
PjaVr/BLjGVh+qnTIi/7aCkQvk6bosb48jJmHYkywoofHPPK5WXMOlarnCwdRZN5M5k/Ewq1qjjz
YOX2P5vX62Dh5v5rI0gB4eAuLSf1pNdtz5V7RXJQlw0EwgVHovoTsKF2C7uc7WirOqnatEtrZXq3
5LM7TjJqU+rZsvaV/LLEP1ThiVUJ+NHwK1/KPf90By+EekxVK4/JW2X4Vuysyt1QX8O3Mc53qHtl
D9ZWNL6665W/WbHJwNgD8ux42bURBzIv/0WTBn9h5G0+1T4YklgOLZgcG6NtMtICV00fUgUSftQp
Ujsxs73D4QRS8jJzZ08IsohiTdpwBqpbxkzj4jP2LlX+D/Tsrr3AT++32rnJw7bYQEmRIC1kW9Gk
WxN/j81Zg5QoCZMkAiS0X7EarMZTk7MmabrdkpTrPm508JKI9bVGig8OprL6FgVgxPSFAsxz4pon
/pa2ZFdcgFD35Tv7S6S/zW9VZFTpUC+fVrD3dA0NmZa8YU1pw2mWFqm9qz7wdX86S+s8dq1ZH+zm
Lz0WYdfyIGUMt/vuSCdivBYlVWEN+7ZpLH8a5PaFlBRv4oLOWBD2r/goiQoCZ/QPNkkTBEEq4/I+
1jryc9qPYVGcNxllvqmem+6DnLApVdb5+TOWO3BRpjKY+kxVoQhbuP0scKc+qPWghJbve7WqoRbV
AXNz5CANFMwdYiA835wfyHe4+SicaYujWybssjWTNhkMa7KIsGoT4cri2g0skbxqRsuzXTJBrrZS
zXLt+3IThuXg6PRtcqu5LkbhFdhixgr8zjtIrJF2GXuLst8bov8WUv8aBhDGI4M3QpLU6so3xWSk
x2Y0S74hAT6oq8cgB4uwgiaKP8Yze8mdEudza4fzYEzGw8W9xQLFthTak7PfEbAdh9mfIlZE35ox
8LXaTo8Z4YSfEAqOi0Ng55oSF0+R/AZej70+3uxr4VEMwkRuVelaFikjaj1fqUKMz6+6KugBdtvs
WPoLF1yF3eKpabFOalw6njtPeBq2lonV0/+I1sZo1QPkWOuWOIT207yMfGIOHhXPwkqTjcw7WkFf
fWw0iQf1DspI3nE4IGHXparIZIEf879fBxWJSmCwTpGXNBdlTPp14MjLzokuGZhGsetZXRvcQlW0
05oOn5bX/wXpWBCoXDXUpEg7voMHXMDL2xa8+6pZM3Cj5wTF535g5P6aT8uBXRfz4wCQcShggmVr
ePgcSLVf/bg+jnps7+G4M3sjhyTIHhQL0YcBbEQkXjmzzv5kdv5+B5PEKSeNB1vxTOaSFKez0XKL
K1JzilnflrfX+GfDCYnJSo7maeBS+0lsxHAsY+cdnBzRm7RKVeCtMqSWvB6vtwOvhNqRMflmW5k9
fwUpMwKrhQv1s8OqeEGaojYUcoPvVKIzl8Dj1tzRjh0mTAOSfVkGOipktvjqcfeXgHZqXIhS7KxV
ik/NKV7KXHnfrA+yMRxT1udEzUFyx5sc6ZvI/urYPdhX9HIiCRSk+FXb3woqKnNA7WvKvcBZN0/j
qX+7QgH6pgFpxXtApXsodNM0dVBD2aUJeIzYP2XWPhKuEruitAXxChwklzvSOg9EVCp76ZUKNk+U
QpWolFGnIlyN8iWdZ/zwLBdpJ2I1VZkSD6BcptKvuFaKYCKCVjIjyw/tfx3LzrRu/nLGK5Uu39hg
IlL2NfXQOjhUa1BirY8dXrONnQyY9CQ44OVHLr4r5jhVt2XRvTFLJYnoHSFik0CP/noLpNZ2VnLr
nXQnLdxDnNDfQme4AFUVxXIygj2ErRzUqhzYNXtT6jKiYTDyhKFsyZNenbZZghF1lN9jeFyklSNM
c5l0YvTqSEC6wSl88lbr7V7D7T/Utn7fp+jp63g3b3PIK3NQ8zpmscvy3E+yZHEttd80BEyLHUAs
pQRIMhbRPP5DMUuJE6IGEsFS87D0z2j7zxc0TCiHn9aLcImCdRH+p65Hw4DlX4d9EXaVMu8KwC+c
usJL2Znj0UXlVmw2+jLs45xZnTvqHm6c7IKkLvjzaTwkb6hgyYoi6/51Y3fVsyrxOzEYQbf4dEAa
zvZdZPoQe5Nr924/IBmuUANDHlFaDnK0nNRxEqgS6Z6i4uDVyiP9EUp638sNV1giV8tjjTr2TVo8
5P/Ulk1quapLLrE29XIBvnveynfB6SQ3wAUR8tgDNiwTDqv6JfAJTGHiwpht62++YHIq6m/Rnrn1
ZoH9wNx1l0KBUrrpu1oofxBUCgTExRWQkShAOHZmHuwd+sQT+bGJqqNlyZebc4AMC0f+sgfdFXsK
AtliU1+N99sC+ObUCP6c94ceZkDfU9NlOc4WZI+uodwWWwqgGTDqADKRWfgD4jC8M4CZ77VyN5uY
0GbuBKIvHo4K5EgDirwMP+/EV2hyO+on20He6XoOSY49oaAhC294ghNwqbJwTdjNopAQ8g9nXmhf
zCRJEi261thYzrLiT0dQ9JAE+VtpGFQ8G9zACtVG08qFV3fN/GimWSPATb1iUux7I8O4zmbXZXqf
5SH6z62vIUjwYRTfuAaFs+x7kdI0nPMKcsdjIS2wz+cTp6sevHte4APshxw00Y0C+X0TNXrqpEBC
mKuPnYkcH357z4rOZxDNCAj+y2QpBKFfPT4/M/wxWszAxCgF1KlBszJMSTqkkcUY1LoE4gAcDoQt
OteUU8dGLGOqjvMpw2bLNG5SwFjmolUQbstL9lhEi8HAtUDRYqePQxprz9B7F/VdVK0Bht9BXzrR
41cZJ6kcun2ZuXUr34Ex91kmSO7pBT2gzoCkM+LbylSrL4B8daqx5L/YuPwMSj7b+AeXRxUcRugy
9EuUmMDOU3Z2e16/+3eqaEyBrHo9eqracpl033LL02NooKT7slFLaSoeN0QXEEHWtQ/RyQwKUcL1
O7n8oxf9dQcrpokTpSmRaJpDta2s+HgWwYsny9G9UBgor7gMoYkm2WTIuretk6NURZYozzaeZsex
2NqoyaExgQ6pejHV37p/M4w8ZcnOErhD49mcNB83Ahji5sZhJ3y8kti7DjFtpCpHBR3virR/yEf6
9KmL34RRNhs71BmRrp5y+rpT4nvkHg5yB0gMIdOxKYlZfs5ImWZXbsmAHp6gT6TKhPyMEWOHiz1S
6gD0jrJsp2waGI9XwuJcduiHNL8XBUHjwYN6ia+nRNAvhxM6BZjjf679t6PX0ZRPpadzKmG5gurJ
W1pT7i2N5P6HT52KYh/bccqMStQ/fS521Ox8jK77P3okMeYX2qvT81V6suTyntHqyDyKLUtKozEp
voenpQQTw/TgWvmGfYT/axYSHCDPi78u+ptrEbhPwEAzkzrlUx4/svSPsaslIcwcxy5teX9Abcaq
o4Ha5EAiNygMkOcNPuZt8xFoRjNNxG6S8hHS4GnMOZ65590QufD786cTE1GRyLj112Wh2hh5XvPc
uF3xUBTDzyyw7uPbzOnmQsqKiGT6QGVd7NcXt5hAsCFQkqdmLnnNShLZl5lvzgSiLrLhQncttF0g
kIRU55q+vbKxVVUDyIxgw0cs1YadXx5GiVfeY57RnI0fAl8S5zDbtzKSkWeGOIh+ZHeKek0D1nW2
FitGTaHbICxkRKjj8NR7gjs46eSPun6CENqwTrZSEogt/OyFxAPWLNJyjNCedKWgls2uzZYYPL9i
Jc+Wm7Oubwx31LaVI1zqCIPrcGM0ZljqA93M/Uy5yU33n1/VG04naFL+OyzDnyVFYcaADkshH2QK
fa/co/h0Ow5K7Nv9NZy9fpkpZEY6+xzKf9xqaKPMXHoFybACawJ24VeB+pPa/s7F2LdtHICjY5fq
h4F7yfhPD8wKW3qImHEey7BILb62VJPFnp5j3zw+An85M0IJmCIMVUvAPBKFdYuj2kSr2fxSSBgM
Fj+OEerz/5MeR/1+mYCw5Wc3Bjc7C30GVNDUtJ46aF2SH8nwnria/h14i1aIBVilwvd7eXZ3TfkL
OFX1NA0QJ91uMHy9WDS2XASxR+cSTa1tTcNMgTyQRZuzb1x15F8m4yH2OMtwFnl/r8V90MdgDuCX
AEzZj8Z9WI2sVf0GxxTUu4PlZgvfjBMpV+azXB3UQxhjwJ2UwS6ojO8qx4dZ0YSiVpv1EXttPe+R
BglhYuMQyJVDt2nPNk7ftfyKgJO4ETXZ8qTGwr9M5cDDXWhAHWqyYbifb6IW+6SxxuVjaf0qnNwk
+1hp2kzA20Bkqb8XjPqZo4yzLo4t0GmyNSHVdGV8JxHmyHBTYmc8aFLitzse1iREBfSTHCSkAspV
x8wDgGn6n9OsFD2ndsEjYELXGENQQB4PKgDtvjxzmvgKQX9026AYRxeDaT7+s9s9zVk/zh9a8kOi
u8x8CAUQn74JEfVk9F7hdGx6ax3oE7SZgR+fXNy4yCR6UNb/WJcXSJ0HUkRJyEoE7EDOYyyVZaaE
CHdjXhEUP/da2mzrVyBXaPAvZnUpq6GVMk+TYcs99JAsiGA/2eLUbHWGoItllpMNggtHqgMD8a8E
RbWfj0xpsMWbr35Mlh8vMHZuzhuQyCrPZPaKmmo82+g/c19yQ+Cr4e0fKZhHDVN2Ov4a7A5jKJDv
G73Vt0aAIJOurHvmMRZ0OuOoG/q2yUr4PeFxksZW0XJXzmyOXyiPvrJhwPlKYelKRL4LfKhNLd92
2wK8r7+UaxJjmMaGlz2PCBU241z0GrZfs8JNOPOqeK0WUU//bmI/Qb4zr0JC9ZvEg6qeXRNoq955
i3yDRCNtO5vuy8vhGvEEdQ0kObsP+5+ZE36IhFE3d36D0KGcwO+rHcXnR2KtxDGRpO4be3wUiyvq
Y11JiIVEBGZ1dRXMnPAshgPp7otivAVL0AZPdfkfL4OKlU2HgYkBzP8zKekCKOidykw6+E3Fvilb
RbLAjvdp4TdERIMZ/JAe5sfiEmKW96HYs6xc+b+iDjUmNN90WC5nR+B0VJPTll2uHbd+vIqQ0q4b
clNQEqkM3ZGysX7KjypG0pv4Br2NRxsEFIdJsF5GCrS+pTEF1UPGeNjPBivmjjMqRhe8fEWVBh2W
9biP+fI+2yYLt/IqA6TGqYJJjrAQ4eFxrbUy9W87om0JRybcIxpc8ZVS8nseKDXWqdLFIq7bc2By
Y27KmjjWtgh8E8ePE/sgcY+Yg/y98od6+jmJdfRmiWjagrlax+VxBXg8RLjcin+b5gLEXt0TjTKm
cIPIB5Ov8reIACVgnXHtXGxQejPvu69hLyWEba0OX1lYcXjAdMNAcTcpfpPoiLvkZGEdAUe/pXp9
ZC4Y1R2pNJL7I49Ly3rSal/d9pqo2GORwQMWW0ZU4yPxLiMiNVxG6io+Hd18XCDAVB86mTJm4/OE
wFe3ig77yRuAV8YUJxZINGFx4mcMGHbPlNYcIgvleesEtuuda1ous6XaafvuAWpymATLR7fMq45v
s/rQoj4XWFRJvF4FHFwchhmy200tl0o/ZUAnFh+Qp8oV67Ejvk6s4q5+IvQN3wPUkjx2shy3mjkg
bF0qQXMshRSFpqGcpy+MkuG4/7NmZZwiA/Phg5tMplf8RfKhGEEoq0d+/pxBhkN9nw3T0NQbGQUI
9pWfFqXqatBMdNEL4LibvzgAbI3pUYc4+WRwc7erP28f96+7epfeoUzuMC6twUEmxgxzrSpIC5El
9olM7Cw1ep56YBmGfBv3Mo4BahlLzjvJ7mBTpRCaL5SK/NCwS3i9faaO4bMzJdhcirxnPgFALPIc
z+ER/8+TFAyjBb70hNVBqGpCNPlTuph0YDrysrTNEsxN9dcScI4ugFSrwcySSd+9HthEMC0Hi5wb
zx+H6FfCW1fQS/PwpfF4aggbqqkwZ/7civBJ2tbH06nIiQ4HE+UKGKn0WCwtgK0btU/Dro203I1H
uh/zOIzE85lYL2TJvCviTY9Prb/T7VXmXs+mAYJv21GkK4SuaPUzXrWaKdfA7EQm9fJiTOymc+hi
kuaEarIUEygGUhWT/VkFi+l2he89z9GBLPGQ8jVRIllOuNGeNli6WQUJy97V+xujYGoXMYd+enGn
gO0hUJCIKKxaw1xRGEHGwYwSA8yF58GdF7vEpo7DSh0yV5ewnW2KqHqypwpV+TY5yVNUslET8r7V
OGSMXYvoPxG0R7TX49k1cxfO1muy89rKLxDkEq4R0VFlYr4P2aYbZ1ZPQrR/+J/MU0VtxG18Yjf8
MYs7pwsQ40ypN3OY4eJbYkf0s0ta+Quvaybs9gEJ0vQXgP6SV365j1sb01XmTVguZV9nNZKNfXJI
Gs+xaxleWtjVdm+KT9o9y//DOb4a8dsp9ANcJ9REJNA0h+FpyW06SAd/85NnIZExAgltzTPcCJNp
pbXgTtsoWC679+jSxpR5PlHFaTg5hxkndlmnXs7K6HYRoAQ6kHxrBUCSwO3ye28oW2F7RFZDQMfJ
eW8e47zxEpzSJRfQMKyDq/RJmkr0iYhQ1QYn1e9C+147wYIyu+R6DHvCHEn8IKGZqvb3lO3sho99
gQk4yTkQvCh3xQksAZ5O+iXHezRVt9BGn26zluYP6eMFSSj+QS7f3ZJhZxoYRpRZp3SEvF28dbLo
+QJcl/h5Q8+qnrXoq00waKOFeGVuYYZaM4CN/ftJ1McIfvhhWgQFSWkn36WVa9X7FzL0UkUgDWJC
oMRt0X0Yav7fKODVJqPwQ8iFKph8H3tum+PujmnWKAOCDnlXdMzaKpTprSDIAMj+TJMFsSDD+a9J
F3AIjUt1T07x1oWN3/PNnpKY4DMh5x4Qb2SDwr0CGYr7r32ssX37OV15cYNfsYxQ8vq6vNm1nkKy
6fWJ4fEo26/qgQVjD+KfpdXyUhh+DfF5po0L82F+0iEJTWNgV3o55f4eiyvsqkKPRM/MpCp+hTl8
R556nkLLdloa7tRtPkrQpvGfJujQ+74rtzlJ3cIIhWeMuXTV3HjH4Sgd9F1gEyyJCIXXJf0J2j14
rhy82hKVXbBMCCkr1jtJ6r+qUBuR1cDJY6obvwUdnagIz+eykhAHb9MCCdhUkIBoB/rQn9BKVW6H
2oO6Aekj/0K3KOZ5hp5AtxE3qIKEBljUiN2sv/eumb50hKRf8NQaRZ5Z9IIh1gSE1gjDpHpq/3X6
nMFvboi6R253+othxvX/rxZ2Md5DI2tOQTvFonGrOwXOEbeKwD2HGmspQtG49E51xzQi5mxM8SuB
whd6+a37lm1XrWt/pTEVAjxr80u2NkaO7YswxqVVvBHBM4Ykfv/h4ejoMAwiwGUXF2NczoR1Z4j7
kdXWU0OixgoY6rUPurJl7j4sL/4Td+JrVC6y2z0EUYc8uYAT1LFIEHrhw+f8Hrc1wqap6mV/lNJY
F+3OaAchDFnp/LittvRU4pM1sgCywUZZOg6oL8yw+fH9DYAVVZx7xkZ6wTW+joYhEOfKc2gJNFod
kz2xF+7OyrDXesAVQ52v0q2Q2O+q4Pg9e1IbsmBksq65rtQ70ShS1zqrZAggN3VbMKHcWhVMTeUY
693Cjj0l1Ci6yOVInjSUYki2NEuXcqPdbXF0l3YItSZJzbjX8DM9VPGJ5nIfONjilN3lAfxDG3OT
K/lwfnB3Mworjrbu2lmi7SInzm1KNcq9MlYJifqumWvmdhIjJRksNb3k56KJ3y/dbPWsPz0Yqz6C
3sbewPqty6i4IGmyaAPQl+cDoIRSuHLn9+/HUz5VUDFceoy1g09tcE/DfO2Z2WBrAAd8M0dVpXfb
YemuVRQjQf2KafILEqOUlJbFsywGrMKlf7EPIECe5HkSDXf6YrdD9L7WMqobn9f/6K6ObAqwiyyG
ixNXMwpiP9XFw2Wsr2dEe9Sv98vqEfnXQyIvPrO9Up+dEwhuZX2OlCaAbk0l9n1GSgGa6W76m2m9
V2zAWFVGnTGHddyX7WHf43C+1BpcZ3A0zEE31Fc4sczYobya4fiNWEFBpKt+x7yC5hcYBp5wlCgs
FyfKunElt0iXGq5+EXsAT5W/4IMeedU/X6tJ1khqP5V/zOMFazHm/Z7tkSr38rKsQdpeyLLc/J9Y
BegveZsZxePdXxdSuPigxKkAuUrED+dlzkcwnHrDEX5w8eMUUIuZyHFpXU4jcbRvQRQ89L8vmjeu
WBiZgLsg3LaRG3Q+kryMk+9kh+xtwOMOgtt1TDUOCD8mrO39IO6zmJIJwIPSJ/yk2XFFZEjkPcQ5
ivqTrWAEf5HrjfndLY48LNS8G+4b/XVAmHiNc+mcMZPSstXdJrzDWEJjTM50ELOOhx0L7VbXLGOw
2Z5lEJ/+syOyJ4oouMoc8eoH+nWDiCmNpr0nubBRBh+UwnecXHKGbcB7Aquz0Mfkb+Z7e2pbyIk/
O4ZhRksE6usSzzzggSMKhDp+RA4k6lfh6ynQe9iZ/LcZC9Swue3F+wt4xrEJDdncC1+Bnz26dnWx
8oTG0IgJ30Uqd9fo3sxSINNNzUR14ZLCKm1i93sNrFJBL8hzsGL/7Fs7BIWy6u0saL8I/7pS9iAO
fo+pbvac+UtjQZrIWlbTNxORzrAh7jkEdbHk4sgoaxgrg9905OCEyBEGxrZ54GI642/kEqlDlUwa
BvuUP4MjG5MOVk5x78r+QnangW7zbfIjVy/PeZ+zYsfvwIG83Xik136gffjVFuuvsfB+TjjcBTP0
xKGd1obPf8Q6Nml7qFWnLjwo6nz7geBce7OG4zzgXnSy3dVBAZDWtKzIuQ2ZOOicr4XF8kl1Ic9p
jVv59Y3TRCc1O4tB97pFCrZ6ItKLeojv9fDEJKX5vX++QAU1+x972tgJk4he7KP42243kp0Ayu3g
CvZxwf5CiODOipp7xHRcRq8nBhJ75U7lbjC9R7JLLlbAiTzjW2/QPujMtT7Y4757aybpFBm8Z+Ya
SfB5Z8Dk11arsBmabytjwUBAbSI2JxIa82ctakmzZSfpeEM5/DRcp5pP1Iz9LOJApGxf6hU2ZCSx
J3i6KKuT5w93TfSclu+vTpxPqMEAz6nRpm8L8t5yp0oDCIirMKY7F5yboinWGNjV90PW6D3lwL9p
hpj+imj1YBmhIFz50O39PDGQf9WrdHFySajqPVJoU+kOTDjhWH/qLldBf4AYeT4h6iKKXBDm8uzS
ViWlDxcZMfWq2ZywANuNAzk+45ZWh/3CMWCa0DNkjGTDPPVCbhCb1VT2rGtu/sHp9LGFjAPjFEWy
Wakdn1eleh13l7UEdPc+EawyLKHMJ6jePSK3+PX7chC4V+f0e+5/IGbBpyaJrpSp0uDmQOSs72pO
8YY247c7aX5rS2pskKHAz61jfx8uOaOh2NuqTjMjctkM3Z5Rsnt36p9BI/jbtHMHFoQvQyb9SyLc
OhtuOrUiYSBX7dakLpG3xkw/bfMScbd21AVmjaEHKMojko3vILZDxxNHFQ2JXfYEbO2eakgO2pFI
WElG/B3W2KVkLorlAQygRxGPBBlIgmdOJ5nyu2yI0bZiuRBqDd3Li+MV+BZ/dLmraHQLiTG1wag0
AwU/AVTlZWtM7GZ+pBYfUsYY087ynGCuMGjJKtO/vGPv9hxyf3iTdOd4hP6oNi9elAZl7MaVK5l2
q93S6/zEZ+7DF6oL+bUQYvgFdsccSLLm3Xe3Cqjcezw83dKMh/4RsWfZtbM2EZLqrDGx2DCuQvNs
TpOl8ODRo0h9lnvEq7tysWcLRm51uYdzlFyzjRjg4zJnP6b3PxRSeRvv+5G2Oe0rMizxRxdd7buf
51OAOK6I0/yU0PUpbICsKr+sthSOuJfncOvpK3Y0gSw70MUT4c6ZEP7GkruoTF9+2c3ZJUShx7Pr
M9wJnse6t+MyYwphkJlZ8gXSUiX1q4J8z4fGu5g90YEoiBZdgiR07iQSO/9LvcQ3GZJDGLH4AK23
6jZtQCRBLoCTmTA/frDz8HvD09CQTHbJgm+EaGYgcQgAR3dMf6JbMML+zojaUJ2vneuHnnUYnWGA
cC0feL6LMmrpg9mzFEkbnP27DAoQE1lrNay+gNFaPLQDEHn3mDS+auLodvWzDMa1MliRaQP+DVui
M31AfVszLYh3WPBPDFRFbXe9E7PVoN4qn9ip7FStEotSAlgT7r6RztzqpWFEw6RfCj8d9A6fcNXT
TQCVw+oA6aSlS/DfDh2fS0kJNYgNTmOqr9Fs8mDfyrCqQzU6Z0I+aatcmWc8GPr6Z5M+79fYtFco
qHtIsMbsv5E2dPIwD6ywNkNslqbatrjr2szaj+8kHCkSEQTFzPtVcfGCh2jz4KM/gssiGOgJZYYR
5kShH9ZJuujmmwmACTNnZdtOSIvAviVckskkKPB9vNFLO+jw8d8NCDgGDuaSLkrQySMtbiKTpCg/
A0Gay0bPkKQNsw7jk4qD+4Se5uD0u+kQmjtSeRwWdyju30AieuF5tyQt2hzscUvi9T09ZmbZYZdW
95KWYYtyH3Kl8bbEbNY08vpfCeHf9iViEKKwpJ4g211s13P9L+oXJPawHBCClijDUxHkovfDm0Z8
PcfatomxhQjdcYeob/XB4jhKHxhHQc6mEkPwZV9hLLpC7Ax/DbhidwH8y0pZ7gMKhiC3Qr9gZBoO
f8fRjh4+VE5kU1gpKi9lnwnJdzvJj1kI79AvdQ0Q1tlaJn+0NB/H2/cWIoQq9/tP+rX1Tl5sSYjA
h99erDlvmYKlnz0G+gl8tFr/bn4IENVUF7+QHGBjvezv0utEygUuOh2jsj+Bpvv4FwKTdOPw1piT
UyqvbhCNkEexDvxffAnw+t161jOvcy81vakOlricZleglHVfGZizxoRGnGQ9WQiG1xHVejupsdFm
iLJssQUtHar3ggH/fk0KGqTQmXgNRn2F59KxgJEphDGJoIARdtLAMaVOQqjMkZm5tCLnSQc6MsS9
E31iQ9uAWmu0KiZuwgq3UascyM9FJBZNZg0BN5rKmplsuyEIkpF7Np+VPr+bP8PF2h7aKwLvsjS5
jdJZOL2F1R7j06yBFCVuXmD9LJxzjzRuOmJeHIL4U5FtcsLQnbwuBVFE6uf4kkRSGOE9C2lS1a+I
4oohYRcsHgdTr3l35XkGiDUStGt+YczczUbTpPhKG0A7DsTwJR9KP9gCleabqpTs7TZJ8BJyiJ8N
74qlx37zt2PkNAeGb+5yHDuzS6qcjt4sl1IftIY5swo2Pzd2ExKj/7AfNkJeXuPr4C6WhZMFuEDe
at+rtC4ENWfUvTPta8XsGhywt9RprwtUBvN+TwTB6ZsH+Fqvaq8hn8FpUZvifts161pIMw2ZyS9S
mxUzpxEp6E2x/viaOjXkg079Wh6a9gWJioTXhh/h1bhAbA6KaBnljenj7JKb6DeuVfWJ7qTIbPnX
o677ea9aQpYb3gzypGN9PLbxVvheezv8f4KvsFSaXSuhNMj+lZ2iIGSWFcmBrvPDEYrsXLZFUeVQ
LrT6kBLjxFtYBRxVA5+MqcbGJaWnDaiX90GQRdusq4epkKMVyRgpp0/Mv2EiiB8pB621slo/DbLk
WNegT6PZc6hMQoNrtx4UIFbVYM4/ZSaq2+IWqde+LlnmqU+4SlbvbaQ9XiV7KBpIayDzSYpD2krI
omN3DMFfmGYuDq3c3u58ORKhpBztCmLFRQAU41pdYabwG0nQ0gl8Y2JrptXRXMLhGyH5kD6eJPOL
SzZcPtOv00M2gitBnqMK4YZaoCavRdig9cVZO71amGbqqOav7r9PwCgEtjfTCQJpDL9JOQ8fNtUp
tRsl8smFKEG21yKLkd4ncHYuY4rXE0P/S1OKtEqKnHkzOQvuZLwvmv5KE7Qg+YWEv7lHT6S5KCWO
H9/N13clp+S4zCIB8GZx65vRFHt8jpKIkpJxK26acrG8N/D6JgikzVrIAmOgeo9YIG7rZh5lo+Bo
Vuqd7G9L7tm9NKeA3CQ54ypUWx5YviBo+k3Bch63DiOehx4wcm0DtAbvjSXwOSMOU5vHTMxxU69I
ntkTioIyzQJG2fcl278igUBzJwHBfO/iQNuJW8X1zJzqbcXBRgiTZTxq4tZc/PPFcpjuej54oJE0
hZG9FrARpe4i+ok/SgUkyONVg6LOlGggGtP6P38r1+HWBsvyvL4TiZDqF6QXz1F5CFofBAWHRTn+
G88he9qRISsz3I54th6ACsoTYE6hWm28ZT6ACsi1S9hg7mnkkz2kXu0oaywwKp7wiIB8VGD33sq8
9t9ZTZgCslyrbCITeAyhUUkNb2xltog0j/4AcDEC4ap7g5L4y5WZUfzdHoAMyto+0dX+DrpcsTV+
RZp6yGNLxAgKFDqMUe5uMl2lST93jj7vHtAmECmDC3xi314uT7w/in9jbF7kP+uYSbO3/WR9hjQV
2rqdaA/18bELykUW6CEp8qfuAuMfmD8lhNYbV33aUgh9DWLssBPTTOIy/Z0Yeg0zS7lebXGrxWL4
jeDEoaRzdUrTccWVVOqkTE032swuPRmVNpBXb2MGl2l/u56mZp8wl7RZ1Nlj/Jz79jVMP3zrRtSu
j+GlIrTTLFYNJ2HiMFHvbBP6dwtCnO9Yn6F/ld0EYeTL3vzRO/qb8U8UO4kdDOD6IEBIwxza/GpS
RbZBM0k0g+RknKEuqg9zW3QZfZCrmp7TFAVLp6dQ75WQ8ZOUDXZJca2VusSZXOXAVJajmgLflnoZ
q5EDLQBeqf0gJZ+TjiMMfJABUmTQSTS9CvsaduMCUrUA8Gszw4/4mV5De3UNIxWV8O+Q6NL4rXHY
4wh85dM722J8Z4d4wnXGhMK1Cjk9g2HUFY7Zn3R/yL503Np9dnE8ddepWtOhfD6uwY3g+64Hjsan
RTD+6E7SPcEYxpDROxEyuRywsTaQd2xinHeB8WyYfAlbd//zmajyqXs+F6pbg+dqnodpvp4wdV6J
Z1B7BGC5VngfQtmLId8ksv5SDA7ZBLjLFVug7aen9tjSR2gjEWMi7PeU0/0xKfCTfvAXc34BLvIu
ixqM7ErM8mvN8Y169qpopZcr86arPieOsH5VxmZ5AaQnU9POWs/Adar7HPF/9LkOgzL1ODtlYD3g
FQiSj6x5fDYZtoXrmHOsERR1iM9Hlf3LwcBDza655uiGtoiIqHsVwUEFbWzAjrNwENvA5gxy5e64
rVfU/kgrkSdpQyVTVzogEjDxhRJDh2q4Cb3FMBuuD9hVUNwaD4VqcqhPs1zZ59JCxEBQ9fnMjgYZ
+fBWrBa6jYwJXKGO+n2xcAfEAWRWV2SjFntTT1WlPlxdP6xCZ5FEE6BAyBpd6Uxbhsp5QbRJG9MM
2qJ/rlAAIRr8KHK8BpmM56pJQQaZ+XqluRbDtKlcRYYjxHkqNmcJ38ofNqoiedKWfFt7n6rO2iaa
qfJ27vpoI2BknRpcfQi19nIL/2n5/8LC4kkltcoaSb57Yw9o7RFfDdtMHBpb879KvH1QtrWMMrmq
Q3WqW1THxNPMwZagV28zOVVG0ncjOjoA952fNBa52xCwe0xPua64oeDdpO3SH+Te3LP4hBhcHxWt
LhmMsJiVQAQDlJp2k7aSwOT4E2vYtGDxwefesLpeg4IZluzWIbj74+fztfg/vpcblw5xSqkWhpEX
zV0wXhLzfwCEqptQBVkOUjwtxy6ZnXu2TMhEsSlY+Z6J0SipPh/yoKQ5wwOEdqdLoh02/jMW5psN
S0dyqhxPRftBHeCZaO2IGrhP3HD87oQs7wzSET8ZSmdCONzZvN/KPePCUgYReKe7Q+eHBImHwsu3
dGEfvc4qptg8ZhvVx/zK9oFTh08T26lfYXx0C+vv0PM5gsEayrEfDsLpTJIRT9veS+g5UoQPvHfH
Cxa+Q/FsCPmtTdgC+84yPpwl+KXRCQnjAgf/3PMQkO2Eer8+/I0hmiLCHxPcpYwiWhb2vlf+mBdO
YCW+lwWtWto2rOfYCIngPiDarsI41rdmtkf7H3frLucR8gj7tprH+OgwETupSPiIaF1VP/s1xtly
mQE7K6CF1HpQ+7wSl1ohCSpOuckjhOPwfwEf7pp6NEuD7nh5eJ1Q1l2OWVq3PYZNEVNnRRFPRVOQ
KyDVS30r7c57KVxs8yp7+cY6tGN0wDOuuub3dKwbW09E73nnpBWoKlRexXxJFp1BW2JacCWw1hEB
DSlWXLhaREhNAM6ZyvFdg5S4P5zT+b8amXG/s4llBdE3NCWEA/UPp0wCO0AT/VrkuiyZUCilCxV1
znpqciGcTTkiUe9RTFFgbOePXREKgtOUSQzinoSbgsy4ra70s7MATKgSyF29yKgYgQikoRAVczWF
B58awMsv7HXR6FRUkedU2smzFWKMxVZ1SGQRoWWr1FC7KAPlYT0OIxY043YQrshwstC6r0vKN6C3
qjvb5GKhTPnr8LpD0/DI66pPBaAtLbH1gvaPTPexn56IP+7D/POYhtrsDd+3/NlOLjdGI9P6+19a
wihKcBnILT6iNeklm/OUxdoyHRa2Vhmkp/hKIOJgajgXhihLMkNFq1+OigFwVKrEbSNZuJ4CANcc
AD4hFekPaeysDck2XK6ntWg2T4jwugw6tXL3mCWfrgAQ7C1xQwBvi5X7aYsnhDicEzBe5L4UsrFC
9XlAMYw/89h8Fo/cl+kwaUNzzxBfjD+KkVsyh2VXuFL81guW9obirHEriVkPLRMjIlyN7buNh/7b
c/8Eogg4gslWYdsdKWaRd0U6MCK3aIqjcuJzQaxNojgyZMUePs74GkCEoFdAJLq/nv0PKJ72Xu14
KsS0f21BeSXRIjpa6LcfEOTQDpU/etD3Z5hevbFNePcbkHza7MGxbncmIuVcTo7UUdsghricsYgc
90jttyvqJ/UAZT6BI05rSHEehQ3yw3YFIFw73WH4hfmthjDaJWp8VxPLeIrEYLLQAfERmTuM/1g7
TKPbyOaHyeMj8GWyUpf5sSBN4iZ6xV0QQiP7OkSfrNM4RoxlNZSsJmFXb4Ke6nzVmRJeUP8H0ybP
wIhYs/9cLCt00HxVZOzZXjx2A2s2St6+FnI5mogztr+KWtmflAZD9Zx5Lk8IoDISwnxPKagsCKv1
RMKOuaPJuNUr7RL2kI/OiH+jx0coe8wecyi79KD0qah7ZBtK7S0pZCQTSOelofmGFsk60yOvhQ3L
SeHvy0vHHYnp7zJDD/l4gi4MKAXOZ4RgWfVlhY0XpZ8g1fhJjp0rfnAlpjHT81Iksz8DnKS5YzUi
krlrSphJyRxe/4dZviFVjs05nF0BlYWaZ+6LOlbhUF+rWzGYJl60Vdey5B6JaahlpZGIOoA5UBvZ
C+ZFo5lgKXIhzCrT1JIE6ZSMeXKS0Oi04nJJhT7OKsvZeRKReYXHGUjG9KWflfjKFIGHjRyXjsFg
Yy69p9nBZ1w4PMr9sgnmgRguKBfypAWEzGOvxk+CPo1IAprIyt5x7xG2yEXDw6LyWofS2j38MHNs
Xn2vlgLJXeMqDMmX2YRV8j+TLEHNNW7AI8aBSZTUAak3EfqBa9SUUd0esQqOq7atSDVpngwBwIE7
ZuU0J6VX91LK/x1HWIfm7NHeoAAYFbT3NYmf111toepGY+RKHirKxRw7TAu9Ttldma2hSSsJBhLq
3nxXRNhYA7TLydMaJcekqk3EVtmUrGz0kNIIYl4w4sh6sT4zafVtAqP1J4eL98tuSJ7LavfNoGsB
Cw8sGzkUANKCcJoT2bppE5NOkQpAAXhJOUsDZAayshhx5OqpZc8NM64rp56oyPOR0A1fNoedazm5
8kwXPI3Qukxdg1dRm7xwZ/xjGydZY6XUFW3dP8HfMYZVY1SIDpJUcLOY8TYiOPM9CjImU4+V+VTq
aGqRjeNQMYeVlGvbsPXR2xE4v5/U15cQ8wEzubEoOWev8LAth2y8MtEkEgOZP7rjvPMhadRJcyu+
DGs/siB2TvVIn2Qw2lm+vGc4WWlJNKllS0WLyb6mLqC+8TfwYQ5eR9V4Axm9ufNbbqQiFXYjvBWk
ZttmNF0DQvEdosStPEgBFjiOWueOlTMiR69nxa45hiZMaX5dJPx7r5OF63Xm0DsBxDxsCaHI+b3n
Wy8Hg5EVimHyS6K7XafI9YNSV6R4The8ILdpcEcVMN1YURKpXuLehxDDMX7D47GEweZSQTvn2hlZ
AhF5FE20oCmiP1lQpNmDmUSk+VfWik7aHEelXnk8byY1oY2xg89BjbcJHTGnYTttfBRDpf6ot8Uw
h8+g5xEvB15TbhMRGrJvkmV/32FIt2FXtL4hSDxViG+iA4IPOx1XJ9f3EjnBWLqeojqwgkq+lOQY
1Wky79cb5ZSm+T67bDHZApwqiMllQTz4voreHe2l2pRWitl7V1oE/EJ741FcsHsqlAwSCduXzHuf
y5K3GCGs/z/S2FnbEvn7T1wA30CfYk0xSiO6wC5CZVGpE/H2ZlqST3cn2zdqZ2iAXKk9ilD/uljU
sch4uTToewf1XOWRhJ4I3xynUj+BntPkmsliQJ/hKmWtakvip0Swqv02FzMcpbD1S2b0nykChaY3
mRiI4CcX0Noq8vLDOtAzSyVXtExEnd6L/7r9AXs87UZNMJt3Jnl2/OpAkXEj1iPQ0MCtwtqR+9id
pBcPPmYwgVy1o+ika8ndlvkL6dh05IUXRp+L2hX48uvqZnwyv2fHUO6VR2ekT0p+odZu7X5EluRg
/LQSpFaY9hpM0LU/0fZYJJVslN1SV5wto6/q61Vy/waV8YhMvGvHNY9u9i8D5xwJYqcnADriB326
mysy9nAzkhktoZcY14BOMssbls6megXMVuCUm/kNTfeN4tkKimcjsgtL/EAL5gotbOpYHLL/rlZ8
oTFJgC44OAWiYOh9OoixvJfaJJ/PGLwwmvsXbkPIrz6Ntk03EYbGchhtlUDan4k9l3CuJtRyqc1A
50KNelp3RcjObi2oY75yO/dHaJxhMqskucPDcQKMU/0739Q0thfA9Q+Pd5nLWq1fvJZ8FMwqhXD0
LyD7YshPGTZFjUg2rQF6K/i1U8Z1Iu0L9M+bYQZ+p7hQ9PZmXSMD9Vp4veWxV0hRB7aXvw68IRbi
v0Sr1CGTrsTR+rZMp15D7xmGRCcDzUyMirGFRdbDwVQshuGH0YRcUyiFsef64w60jQ3Cs1iZkbti
HURAOVCXz0VO66/ce6RWSegtGqCQJFExeLjPZHHlfu6TtRlU9YJaD4omjXDz7nj3vOoruNelI8QL
kGllsRyRpcnHH/puu5cv8fVHVjhmXshJgXizuUv5vTA466elYmzDRmpGNHSWPAnGi2235IC/XoMJ
0XzUTJ9gIlQzYp2YsbdgmQIEx48UUXREVaV02WylmH2XaRXCB3XR+g82a3oykooOIMAx2sYaHqdN
HjfEMFX6pBBTHU/atNsQ/fnofpIkS6+pU06SIgdggKkmYqrwzANlPruq8uop3MT+JIcaKHH+Vps2
PHFCvGZFAcE2aUbe7bl3tVhpsZyaDofgSn5xMRJw4B9HkPEQRtiadVxBG8i8cpTzOCaO/wydizNR
DQdHGaojPQo1CSauOPm++XzEiB68Qyafj1T0DtDTwZGmV+5KHML1KFbbC62PDFy5s5LXQi064y9E
4yzN8MZnMPziInRs47ExYunL/xiC2ZdtLqa8KhhU/zYgWMgaQqbEdsVWcUyKZfvs24BOEKhMyB8k
nsMJ/7Q7sAQ0H0ud7YSjyB4cAEtlLwhOR3cY8x7qIM7DFN+Xsyh8eBHaUiLuTEKBQjTsS7R2aQbg
v41ppI+oW3wZ7tzEqRNJI/6q6y3VcziPo7rVpCoe1EyCnaS6ONM6gbTa3e/+kcEdAW3gH8PQq6ko
tezccJL8arFuvY/sWqfhe03MI/m7UDocu/WfJPrV1/d7nEHJ1n2DkzxdXalXhkQ/PaZ+uqbVJTkj
NsWF7fWojdLtiJb1HQRfG75x9GWGsajeQq33D1C27XtTdInoa5QIkE9jdgFXgLNvt2bI3k6rwVFc
jYh7Optgr5PDdP+76Si0hlRpStNusnalcGE9PcPf9wqmS7WEo788a9nOyxkmqmrUlXw5jpLBvYum
5Gm2XvV4L4GagkXizG8ZaqdviEYOIMbBj9OQRwHDGKG4yzb2G+eyioWEfLA9rHkRJD1nmi7+JZEX
ckLks3KlJ49Ae48bOowCCgHwcpn4gHY3GzVjYbQV1a7F0Re3CS5O5hfn0f28dIferZeCue7+wgDa
rOMZ9VqueOHQcLIF+Wm/Wrp0Jwys3oQm9d3VfhFCz15zGoVVEn/sqkLguvvmsOAUcRUKSe7pB67Y
R72bFfi2agJzM4STz7FxWM+QqW+gpWiwHPiPkgyFu6X0+oGJmmd+jIXYJAgWBidwdpdIic7LyDeT
fGVWBiKIj418UwgWEKQeLGjaIkvZeyAJyjJYz4lR0QBQ0xeFTVMScA7ec9Ezrvqq7zgiYEkBEVTc
lZCCSsE+n4CZNovQ4f+ajDx9saAS5BNSXjX0RCNP5fi8l4ZWroMJUJ1VaS+WdCZ0sxF6PPo2Cgnf
Hz5P707vB51T2P///UrdmaX/G1j3dAgo0zAhpBtcNJg3IWq0iuf9ulImrestV56OpCsJp8KnGNzF
Xd8VJokbNMPNFd9W/N/AbheskPoIoBsBlM6BS8+eIcx+8cNhj1Zv/c5IN2MePNCeNFLAEiOoVna/
++gtXcez+2Kp7ZRUfUIt/UUHHvKjKEYP0pmEZLLPKM8RqQooRLfF9lyXRESzUWBry66wsaNr+Hhz
bBkT0I6K/UGPiZQ2scExRsqcM9clLtVGaPMLZ5Oj8gSc67v0vVZYAk570IkJzzZilQZ7ermYtOiv
eJtjhWmDN6zLZC+q9PQ+K4qmAWnwuxijBbGZGowRCimb5Ir+VNZ308yzLW6szx1cL1xXpBLTjTkb
OKT0OFEYYBZX2EDTU/dWiZnp4SC8tnAKGC6l8GrJ5df0rFuWVHKOZPxcVXnudSGzZCubV5EbWzxh
6p6b6igmVIA0nlh9VqPgMF7t31HYM6CbjybX30qjw4FvffSWkmp9MHwrJX9StH2r/+98Asf5MO5N
/Y2Jwq/CZqbwBoqQ0GZrczPKk8ozDqQeeUyNwwZ/pnS6LlpMN7AJb/bNzfMvlWQ96nf/ksNNaMd6
h88qGhuuYMaUCppWqTRHI8Le21Asv/OjCAejrkziAdBXNvOyufY3ZKL6j/p2SNB/O65Zo76OCZiN
I9EonlME9LrXux/O6gWuSSVvxHRsTaVUml217jZa6DTTNn594HjfGL60MLZtvPwqUf2NE3T68XA8
F1UGwIdVBrs8eOp4R8Mp08pkzW3EV8eD2DAUBHbvySrmGhRXgTM1IRBynynwol2+nWBwu277Q17S
OLhW65sD3htQTmaoYrOMKIaWk3/p4BdVi7e4WQCElN00VVmt7v/ZkFbvwTf6V7hub9D/05Fve1x2
2PGf0y4WLURwjbS2FWkhDrfAzmHbFfWT7dyZSUvvs+041Pi5Pyb60fTu7ejK6jT7R5Nak0HubBTv
xEfPef9dP93KjGjPfmvm0tX6J3pL5fzfQiWVZg0wSCm1Vf6WIZ/ChCZCbX2RdBcC13ODR1SlfEx1
B+adJJbDYbdfoLjfX3SAbm2MwA5eqoU/19fBYIMRSGwYMQzCFEfEdC6SQ3NZdymSLWK/l4hQQVVV
1smDLwT1sTlYrIFckJhVjZIXkwVsbVntCstQuyQaXM2XUx6ygdTt3Mypydj/J1EUr14/NYLgGcJg
aZf09BagbJvxNm/MlrWq1IcUBNHG3sxBD0UBhlST1ktSJREWqgnVixwMb1RUfTsAgSUafLefDM4d
Wtv90IeSgO4c0HVqunq0rMjayq8YjLutO0huPxqqH5VvV8XaC3kk5z2vaKaJtXXTRvQl0LbDxS3w
s89wDW5OAmRR4NOOJmRYLXqXIrSSPvFcxWLH4LO2/io2eWoNSKZJMrF+SnEgC02O+0XFHf2NcAZy
XHZn+1vbHx1+OdPQkdtDfo/bUr3t0X+3t4tlKIbfXVTuX2MLmY/81WQnQTVOv+zAjbIsMwHafsZJ
EFSZfPua85unbC6xaObLU0GlC5AlGDYoXp/9i0OvkD5ZZ1dPDd7YUQbNAeXgbQ2t8vDrq+V7DykF
Vxos3GHeXYvjHbF0+GRnu2llmTALHtbhJkaAbFZGGwOiNWbr9eRKWVjo4UHED7fJnFcYKuV/ybRx
0be0AYSY2QMoWFEzY1Vo6eWBfQ86M3BwaWscfuNrXH3PFUCmnToPGFZyew8eZnXDEZgDmJv0meNV
+JLjxUwo5gqGVgFqt2R/zJuNgO5TvY+fjgYy5HCMkDkVPBqXfuvBWq7HEHYoZqeAx595TfyifjUz
W/XSXXpi7/YhnLUIk9Qg/Q41L5tkar8St/wVzd7AwV2W0Bj+w7l9NjATtW5ez3d7PeatTN8eWM2j
kIGHkx1iq6xKloOtqIeKC+IJWjjxDoDsm3PrpHI27Av/D9wgJ8CtLoowEADPOHOzTJAcAbFijoFr
U3+qmjD9xdFX87slvZW9eB6VlrmXe749qFO1mktrQprz4hMzqT3Z9UQCfaBFrXJeeFE8oKwFGPfe
J/+X4GXjiIRCCccKr9KkuXb8So0Jv5KwJaCECAJ+Fdn1zlFuweBWXPTk+RQiqiJZyWeVXZ9JU55J
6i7ClOiFBuJMSw/C+WGYic7YFZbxoRtYZS38ibFQlbnfIRPkojRvcPyKDBKrMGzVzZveZIuazF4a
RuPu3ceJbHDNrOPefb/lRF+ScUZf6QseRbjSJ3xo0CZMUxTvBaiqZf/Bl09ZPFYwnYW/C4FTBr4i
NHMp+7LgQ/Uwi/Oi9srFHNCNsMtXQvjuk9uiuNUhkec3tNPpUuD7VazxbZ8Cn+qMlvzgPo7fDnAT
Jki2pIIh7HY50iv6uTYG3VmBahGP85J/pats14kIjZcxF++cEZvyXXDAP5tEj5S8NYYuGfrU/QdS
Oe+X+r8DkybfCNtHehusoqIH7PT5WxsdTNn5YqHK90r/PfYgnlXU6Sh+oXDF3XRpUZRZo2TVGyic
9fZ8VP/WEnCVg6SnOYh8VvvdEPKB54D0w80cqYeHH9Yh6RE8UrlCRcG5nLGN/uUMvizAZL0cu9Cu
7TSCCgPExlcxI1el1RIXMb4Vd8NEcG4RxhPISkKJoHhOcduft+a9cjqoBpLoqkrdYO7K0+5lG8tQ
wu3OFgU32QBmD+BxV2qgMcba7AC2zx9K1H0OYe3cXxNPK0nylMFKD2LAfSo99ZIU1QU74P8Q0Z0n
IRWqQMk99TIYhENQdnRvrmGB4xgRRCG6MlaM61/43xehkt2JbLkpstNBJekKmlntmyprNzHJQfiV
tCSFhE19poa5u+JhnRxSfS4jBbCwra7IA1F9LybeMJtsViR+tpNHbQ6qBcB/A65tKCYVDSs+zMmy
pytilbrinFKMnaAUMDgqAtkAOjH2lNjgEE+D3WLcvwNeP+uumRR+acYrFj3aMtl+GFFG95yCUngV
ppPyKje+3AfPAqqvnJY0wIc3tpnIrzc9VZfAHMupCgTIPnw8gEZDX/UeHHQUZL/eZIMYbZmQZw9/
IKdG+1DbczeJnnFrxQAumG1Hs3xMg/yzLJOxkUBlc4vu9CxM5976MSJ0K3vjBx4HIBC/gzkk0dW/
VtC1Uz+umj14tGLMqHpKldXQFnHoz4aCGWFigfsSdJsLzzSQyiB2RtOA2SYn0L6XKiZYhMr+TLph
nN9D3c0unoSXi5nNXl/aMTjQ1P/7aBpg+KuEkNVeBGk2MV2tAUbfGi8mYn7MDq9goHAwmKUyFvKY
qVets57evjG2zDxHlnT0bah24lm323x7C2kzujBtA+Icmq+OrG6UMQjL1e6O95yLNlNnncpbMwqC
29G69Od2oZ67uXS5ikFAupsUO1PIoefFwBppcHwI2QtELqfR74pN5BGk1QS99sk3yYqH2ZAdnEWw
A/YGIWLPrxxdORrIR5Te3Pu6hTWT1IK9VFA8i/XTyTAc30hMujwgKZLVBV2diAvDjJv2P0+YLjRe
vvhghFlssQ7PbmWzFIyJouY/a4SRAMM1HMPKrcuvcEX03clYHOhTD+4OEB+BGhjwxIG8WVbpdEvl
nM+66hrRCeEAORHG5Qpnm5g9PtTmYaAEmApUgU/kfpLdQSh0jPp4wz1Hdfucu3BXTweG4+EFcgp+
oGG8c5AO/mza9nszDtHXd4+NhjGOb42mLDgAZ/3n4HI/3u//CxCTyF+1lNqBMN4wrFvMh62zs++b
L0FelRKokgGTZZWJmFJpNHfzDQUG5K4S5BQUYfUtibPz7czUPIfC8nzERR4gq6mNw+YGad/fCnFF
gi2b3j0pqLxkZnlyerYfifga/VzQNcwVwmLChy8j6dIJnyrrx3eMxAg6wRwinR+rE84Ow6/0bw5a
qwHdGgz5m7JQUixmpv9sIPNMhnSSdzYW3iy3g0VJ8ojcCyoPk9kl/ztZyr8sbhk9oasLDUCz2x3p
yIlf43MS6gyZrxHeACxpmoIhUkkVAagFKVJjkj8qh96oTP95bJikeliPdUXY7VICLezctEP0KRCg
3lQtS9Rce6s2J4b2Fktzgzn1S26ibGhpSLAXJbSiWw0MMSGxc1qt9F9CXGRi4trbmVTPfPseX6Qx
hHTZx77omNqcnUNtFHxnreeRUnMow3qEdj4/XSy008C8b63yO85FWGFU387QnglYSUrCijo0B9ZA
p94m5K79tp6S5kfLxagJQ4uNsb/yrQvEpWAUGsMepWr8k4rnjyeUOCprCjF1Awp3aZS7RndMG7c4
VdXeVMPAcPRdpGbPZsJ5euyDRQ+D+kFgGveWq7aqw/1VC2CI5eT9wn/xsWtsr2bDt9hSPam0hfKj
Ov2pmJLS+OIJGX6j7Ay+ClSWvjspO/WALlxnfrg5rtmHi6zApeb/zS46usWex9Too34CLAtXnHEg
mn4ljBvaRWFVanUEL7qYTv2sIyGdE2hLVeqjY/V2EDi2XEEhGFvUPEbaLg8WBVKdyBsr7q6inBaC
u0HAHInby8/Bk4WJbMP2G1ZUM/GZrYTTNY99l0RaU3e7kCurRhL1AjHTX+PsXoArAWOgNqtNEzAx
aJ17evuYx+qJUhvMDdAArctBQo0YdMR5h33F+SPYvLs60GnR32Kugb4D6XIdE6PtdWl3QeSVnIw0
R0ssUN70cVxeEP5nQuIbbsQLURoetCze7XEfZA4YhMcSLERvX9TNJk+DLeQeoEawTduwtGbf0pH8
nAs1xmBpuG6E2PYscb8KIcZBqk7/xri3+8MSS4ImdcLrtsGvwpF1u638sr7y03TEm3dkAxs1YQMv
W7OW8Z11zzELUs5nzV3EbQsv+pbGelosACVfrW5LGCgKdkbhx6OxEMlPuCOwfvszGCdJ67Togvko
INeQTpsFFUpeenAMyzaUYQ5LFaRzVz5BR1LhAXxCXK4a/Y1d1+G6ETCdVdIbiruvkqf6qgcY7z+J
WTrckK4KR0kn3/sAQG1tUXQ5zBWLsw2hfTf4sWkySCM6mDlcqkvdEAX52BVQUTAf/7+mGGPaMVOq
VUS9n4j7WEmyUqTw/VRWEfQMfI23F1vmUYU830vuYbJy3NznKNfmnFJVgjdSQrngTTsYloX1nTXV
CzgIjWHnXmRrE+sYNaniVgOyasNCnBp+jQ0sQGxwAV6sG77w8i9ScPKlyV3rcUuEe80smSVTIPNY
NwsQo5DqNBroMQNFv5+ieeMZ+KuuJSyQkCOwYbHLaXRQO3sViSh0QryLJ5OWuZPfZduKl48UdSXc
nD/lErqcRYNtOy530mgoWHQ4V4xv2cPrJ76XlZO9kX58POmT+15kA9DwwBmIuVML1HHigaAUaLtF
xZbYdsXdSr14qDEFwH3MfURVLJUtkLEwAZ0rbrfGlzUrKkGlZcW8H0IFqYfZtFZ/YminGTB+nVvz
Fz8xYfAnvRLY/tqFBGoF7kneZf3LqEg3Ziqs1df4B4IaE8FlQIOn624JvvvpnKkk8Bv8MgJ5/GYW
kfCtKB2UFZcXmBFyCY1TIpa47U3c/Y+DYC6dQL83uAerVR6yfDL+PHDW3c9kU9UeG9nE4h7cabsx
+ro/pBoVLfh1lDd/4iV/N1ozjdGGLNnUVRC83M3mSqARZMNF+4XXRB7nkdM8UESbQDHc5g3ALCEa
kewIAxEVxqhVsRzHsgp8S6PKP/wkaOGnuLE/pXgFc8jHeM/eN+phpUm3b/GtiMq5ihPhmeJ/wvjW
q+0YOluNiwnyVzC4musn4N/FJLOXeXlTZUvLmsuG1txW+uSDIWak/ptrLXtacA+7/IPrQ87O+50j
WFVj6Jtp6z9ySJkmpVZspujlEAfE2SHjvA9DfDCGgc7O0M3dimYsD3ekSQ3meduFZtcEGZXZjoYP
U+K17etwMBUMun3codgoNmem0tKjtANTkBH1jlfrHx+v5o8yQZxmf8BBfcPK4dR9g/W1u4jE0VA1
vlOkeCotkNMOMfKJw/VVgzl0/eP9q1Cq8HFqF8A9zm2N1OEXqVI5rrA93QvMSMJfoWHb4pLjR4KZ
5bS+xoOVvFBtLR7lL4X7icPcy4aw8+B2G18VU6mSLWkiidNoskbhbwrnC0bvawHI+4jUUWwB5Z5e
QKZwXlMjJTrEWGaFv0zwB3jYQZYTyVDgKJUfKLdxI2Ut2ycZuIdhR38MKXz7uGieFSzse7HVji1Y
B3hb8OzQZmMRzqkUqyJOY3/SRpadVlXZlgvrQtxkKyTRdth88EIzNyhxwn5SylPadoapio+IPqPP
WIqFpR5bF/YxF0GdUkpEi2TE6Qn0wVNOH8n92wTogeGf/pDvb1cwb8O5AR/PaHNy10OpS4xQBQ4/
ADYfiiGxkEMgifntInmgq595XLvR9GkSLVU2vuUfeB9eZYwq/ha7nUAustzgcQqgLQw5luByLf8h
B5kO3tsGykcM5WfhMT/b/pjz5uW1Vte3xIMgosgd48MNe/u+2bwuqgCTr/MDCtWbtFAM/oTSXUhc
wkNay1wVmrTfUyHuIQlKSLaq+bqKPfEqOehD6QEwBzQHytEz11HRUwcFx1sgd/5YwB9pmMM9kJSs
PVoSlNYDCzI42Uuc7QYZPPxJtcnp+p/RSJmtVs3KIaDw+KdoGvA07PiRqbEnjecZ3Ow+7UZIqrXY
23jEqJ9GFCKUymUoh04pQ9Z/IFitMXSDjXdw2th3nabtnrAYs7AfkyD+viZ+eZFCYvBAO4uQ0iQ9
UCokKGR5RRl0QyEXhPMpzxd0vqLBlBlJ8i3oYCLmpAxk1Z1fMT6RlPWRt/cB9zFwC/vJ7kDHsL/D
027dsn+yPY3X+0fzHihiCn5sAotIxU+pEhHPm+pfYATOlZUoEQjJ+V1q1NVMBZ/dsP56GsMJs6fj
lkXgwAUiua4X4P/NxyKK38uI39XV9Jkvnyn94Ad5UYrJDtzqhqHV9n/Xofxg/oJs9/TESlP7X+pA
TSx5hWY+nQhKBGuPMefmqlFQqA4lRmNfiBjf2mWGN8ANwuVP05+mj6HrVHLxzxTyUBgD2+OrTuPn
zyFosYtFwU9PfEWULYYdcszTkG2upEL/cUZmHDALOe/g3PcXJGryi4EYtF4YGNV7ZKrgvhtbDRi9
BrPWODLQNfnxkp8+BkHEHqP/LG8gFJ2mSUWIAgNXyVuzIQimg7M/knaR0LiKIVJ8AQV2u+APwtv0
yPVzkcVBDX7qcqdqiVbv2Dhs4cRsyBJRmChme6V/oFe4zUTINdeGZdFt3AReOjD4/hFvTYIXw2De
IXWga+33v969AjdBpKuBZtg4oXCQWBlg59V96gPKU+GNR2SDg7gjjsWWUJfoFfK8OgM4u/3tPafg
xLK1AksDXbFnxLhcXGWdxC5VFfQBZUFq9pqIMjBFcQ79VJzVSEJ0/G7Pd5YIagKimZDbe0a/uQSf
yE5TRjfVAf/eLFG6wu9vtyLL0Kl221QRj/Mu0CzKUOyOKPgrnsmQr+Mhe1niIwU+Zabsl+Bl8IcK
Fa+BxsxRnB8QiD3To05+xp84A2PLBCxCJiDr45vKeXa9s9kHLlgrnFvXuz2u0hmqGPM0jn2guno9
FluK9JLlzCVOuZAgVs/kcpynfYfFZHebmGt4IhpHluWbj3x3n3yuuQJJhJPw9COE0qZPPVvfFcqc
vYBh/Ps/oMasz8PEjnsCK7MuLcpEUSavbWDjTbfv+SHvlAS2eMst9JIqhegnuUwBMVavNXvQQwFb
q3IfQfR1Pu6BWaQ4g7wwn+RH+GIevWh/SRW+2VlcrPwIwNznOVU3h7wVFiQFQLgrhTuKjGEpdaCC
g9bwGCPTS5UEGLYWlvRE20LnuLtzww+aJnP/vq1d3QZbkdAZDZjSZt8qKcVU/KaahPRWQPNEceau
oOYPe2y1bsAREbLRBttK3LYpgBRZzyzf22NyutdT4ZlgKy/K4DVjR8B83u6C1QBBx9IoiW5aaaVO
TLyH0uYMkfH6b48GjmPSvyeA9ld8JJgBvRBVaewsWI9qEB3Hc4dzQ5xjErB949M5ka6ZA7zkJiZq
d86JiE8EHGo0vLc40zm7QS51WcvsBEWkXP3HHRAIQfVqYjN44JTvJ2Fap8i0iJv6NslXfLZdN4t5
Q2AyMf9aU6b97dwFXclmUwcEA/PfqhD4m831p8ubO5HsKPD3WTj9BtHK1Nz2KYHuHBijm/8tRr4j
R4j7/7iYhwxHiIh/h4AWSpk0Vu15JNNMqjFVNMiwXO4GScnf5VUALAp+Z/FcTv77ZwN6BKeqe/iR
R3PWqNxK0owlrYixOdThxgdMjL0wNNXINUdb7CDRjdTQln3OCVJjaMyTr5r6TlqXi6IGyCzMjAgF
cY2EAEf+09mxLEUdsRhvxBF5CUDwo7xitxlkQnTm72l2XVFANU8tDf6IjJheiA81GBiGvOoy6PCZ
OeiN1En2VOrJtR/YXOh4qBEWQitrc6gxGDPVHsuBg43B9yIkm3skQJxiSlJGb/x0n9mEPu7fiIC7
Ks18//pzFJ17xmeWs/sCucFnLw86L+sPKL/479zjlOEs2/SHeZbVZB37duViTPjYpRh+cXCzKudu
C0UePLtOZbcNbAdyDLqvZKEu7BVPQFIwVLrwjHR+ClhfF1tZ/ExXApHiBvdVMTqpLrpE7jf2ad6F
K723dXK4VSWvDDU7v31nLjRRmRlcA1gKNQ1ctrlXmShN3aKG0GwOiCzegWvCpYiQi0yEfhu9CzPL
DjeL2W/e9w+BnjSky7LXJZBqA7ymer55YlFBZR/15VDlOrfw9Hyike7Ls79h2Z/A0KKnnuexG3so
nX6ho8BdMjPspLn857EBWCxGGHiEQzyyejJ6f5EihhclZU6n7OejrDb3tGfQ7xYntXAyG4yDMad6
m5MhkGb4cszAdRnZoWNEgYdFpYWF4ponPtIzkroEHqNd4Du1H/QGTL+CbvTwtfrWsXE8L2sTRTU1
D/vtQn/sD/HJnyGFLH+X29O6cT+mctQN4TPiyZ07I6Q9otc3gwkTZ6+Bf5eRReHlNk8ItbRU91oU
2F7emh65qZaY1bXOx8LA5rZK8vvQkmW6/SWHenvjedQ7ajUvGxgelZDyQIWV+UsNWmLmaRgj4hkv
k/6X4krtcqMlloECUZi3sWGSQqzuOCS4E4+G6GUUH3D3+r0rlEkshxLvwvc3Vf9YQay9m5t+cLhE
6BRf7jlvwQizusm9YSSSHIReIxWOel5vkOWFf92Sb5L8UzN3JEDHd3/f3Brd5ho+VKPTdhnaTKrR
tpFPhgRcfIBBeHQlKsyttHUL/Lu0GpZEgrIu2VLaA7Fzp8ONIDpBZQMJ0KkpKcxfBFbO6VJWCOSf
8daDeQUlsHRsAdCIhzk0xjwRERxscWu9rZ+HrYBjAyxa76Dk14ucl3foxAUuVmZMB56mkqsFbn8m
Qq0dJwd6v1jEPPDFl7hqNjazkdb1J31AaduUlQi8+8IoDuX3JPs+QJqQFMtTQdwFgXjjdUxiu3mr
7B0rl8CMfJdnkUKvuRhQGiRgAvvMa/rlqTtp2V8TyBnbsuq8l5QxXrpDA72mj0s/PhCuyMYa57TF
UH4sYqLCDh0gLjYE7Z0v2jxV6EQmu8j447BW6clHnoUKskR98JbTPKvPQeM1yaeZUdbb/13w/b9O
wUZKm0OCOG3juWDoO3jw2IwSq1elGYnonnnY7ID3ZsLTFrVARIv46sE2cw5niTvwpr9sic+vaQqT
eUmESctIHSkbe/nXtaPwO6h6l/IWSPlGjJsy9yHzfZ/9eLET3W7aDCkO32Ou+w204LfX6cjQFaUK
vlLoz9Jj1yoU5qpF5RsG+zuwKhZYH6vsv9tyrQvIAxl711d418H4Gp3cmuHnf24MtNu3mBwCsqEV
zSnKT6MsSd6LNNS9jGFH+zVXaL7lg/oHvMNRjV7msMNmjxD6qpyNvQAQOLu9DdjpnvyXC2YUbzYh
Ycmdc3PMavpuA3GUFTNa9oIed/zjbpyH/jIlMAG4Luc8EPjXITfFXYHSrV9FWxAcqU4OENE1eEre
kBavvf5yJBsDNW4LHugFByZcV9YMp/l1M8CkvjETjry6qOBz6K2yg9UiRh2yC0xOzvAhTKTQ+LTC
lRr71kFW49yZPD5Z5rfWRBNfxp6r2W1LDl+5yo3b8AyubiLfTyVK88qoY2gp6gueVy8XKEj2YDxL
gvugyq22FGTrNA5R8VzogWhVOXl0sAouFNqQ4mc8mdVdnJGue/cK1JclBMa6G2Buo308n5kSYv9z
QFyAp+ASq1Y7jcKcA1G7EWjpOeLoMoUeVkqANagdEVnwwynXDV4PEUAuE/g0ttxEl2EIxfsmqcet
0DBhw4VJKzzW5nNbsDdIpDXulpQyEOaQvN6YP50MR3VQgkkRK1fmDD52IxtJWxetjIi0WjxvM7Wp
aiIlq/hB81LZsPu0JJ0hcyLts8SRuJFYNZzEw1WmVMlyrHQWLsGIJ4ORzquN7Zf6C1JKgJtjrFhm
U7ntsfzZiKWWmD3XwtXb0tNHLhRx5OLVZ2zllUr+xxFCBSXe4Le6OYBtHrx+1UB+8TdjOvjnOUq/
LpnxfmFHgJRQ0GTEZuhbGO2rgqhDkkE5DM4f7RosmUCzLRHJlzpDAMQUNrLzvxAgavjNdssejvdS
/0Z8ud3XmgpdgksIrw8Qat2rBlJouryPmEDLh2D1lJUb9PwqtmC7qH6NpjnE7LVfVOaabTTB5M4D
l4kY4ezw/jepZUicTHQEksUYhqwAR+vp0hkN0rxhi3QnXnRCt4TykFGsMRD6vHTH3SITMb5GDKCX
llV/dd+Ro29Q7EtLDqDLBEg+QzE2MAPkBP5/+vgNV/q6hsRjPr0I0DPvaoyShNZxkOBPPhx2ZUvZ
Ox2ry0vcrVt8dREe4+mzT/Z5xNl7dhBA2/fTVLHNTuc7McLWv0vRrPEcwYZ/vNMRFc9g9T/YNgsK
hddivHoDhBRx3lQQpWt/JBkwaBPvmMJbrtqb3TQ3mMnenUQEGUQOKGWP6NRnTjpLnIgQH3mJe1OE
cGDXJg2lLF57w324sIc/TsV9SGVOveHOLGLR6ARkcz1QfpgV/ZEaCYxY/epFwOk9e+LHc4tI3QiK
8eV+1XQwk8cUIexBiuIEJMcp99q2/CU/bFeBv0/JBFt8pP+sJyGJYnl4lTG9XLhtWq2Sk0o28frd
GdO3fIqnRVKCtCB22rCXEKVlSMBy050r9zzmc/wpSkN5+vYLOTCiV9stmAZ77ByNXt6YABkWI3om
t6y1El4M784z+0WUH999aPnLL+Z1iWLcqOnOjzscereR6vzuQQgE1suC/fJXXuvcTaOSb6samsoY
GScpLs/b/YTsMAKt5qnc3+TgWr4gKzqQlLwlvQzZYaKIJ9saQSD4YjPjhK5brj7V4aLo4XXNJHQE
w77AkjvdLqteLH3yDiUXM6o/JmgzJH/DzRsnYVeiST/W6nPFVGYU5XbNsSTmpVG/iQ08vHU/IIJN
xlnkLOwizPh89myGnO3JGRMQFFLKPWVDZoZ0VYkS+Em+9kRm0k5JLxtFmoFOpoYp15IjZ4C/TvyC
XqbJung2xAbJH67E3cTA0X/2uVWXzeg/viP/zC0FPhNkcrupK47jabAOgYTXsMxDKPQua6qrOS5Q
5hXjVSTIk21oeyzoUfiDjItW37flRnCTkzc/MDNJgsOdQ2Gn6sexeyaUzFeQk5BTmdoQbtcZal+f
6h1eAZdxhJMGQC8VmAg8rxtc68dNKwX1Hbnkf3gAfJGErnvoz5T4ZceO0+vxBnzZfIfIgVsHtlFe
Xend23AcgxQyWiqLUc25A7hijT/i4/F/qWwc7p/j9UuJa7NnzgW9fXRoTMZ41jj4lb21r2s4X+PK
jDN0FA50FFnEfx+As/0arvY8mqbVkuQ6RyCqZNiq8H/07eKNrdS78She1wps6fhtOR9Nfdt3JdiU
EWzEv1R2eeUInYCkbiYWglnz2a+zsCwrH0qwrIHuaM3pvev1FZbA3yfGgCYTDpiXABEISf0xJDKs
v7b+tlPygQS6JdCsFSlju1ZlArOWempLuRsfvifl4W6C5/aNxfOAXb8mHe4bAm+cCfyCWg5KShog
nkky5emFShPCDoXIOeh7ITKZA1aLP4QClznFtcrLvGowGRX6+wnNaKB3qFtR44PcZbiu82bMEv8p
ghW6a5f8BRcBcbGXGanzzD80xuy3HIZZS/y6rdvQUa5IOan+o1jOhRyAhFW+k4Qspc/U83XJGjyU
oUEdQI/OSNaKBBsRrjrLeWCxXCT8qIbKiPkfT3Ksc18gSzp+TmpwjGQ5OCVPb6D2eDUiDZcOqx3k
d5fnVOnGKpgdoKmyLeMxkY6DgDaYLHF5neNeW6Z3DnMXZvr+tlJcerbexkevwPreQ8sfiWVqA5k2
PzUxfQiu0K/xl8aDAxKqgefZbVQlm00BtHdXEKV9pICczZtygPcFjHGdIwxkoIfZR00mSW9CzKJa
MHYtaeSRXlpC/h9OEC3WpwCRZc+gNj3/NRKK8SH6vI8CYjuvmd0cnQ/FrKfv31lS2ZfQzdK3zLGr
3IS/Y2CKU+Z5H528YNWYY9I6o/O/w2ALREI6tsEhoPT1W66mI0DKmYI5CW7WS81tOsto6Zn0HEa5
9BPMfA30nptnNPxu+bHTscq//+RuDX7LJbVBtLMB8dscKWTBGkN3Wvom43uyZTnHjz+zytd0oKZz
ssyI3qzj4Oz4IiCCrsWd8In1R4ExX4J6sJSUY/nlWqB956OF3l5yVd7xcx0E2aQguOR8wmHMwHA6
eBzKdIuvUyjdaesp6IqJEod0sODBLoztJfmmCuM1p48a1rrLTb8sZL56NUnYU86mLlWgA4gRYHVb
9qIwTJzOK254y9us734z3N4QcCPAZ/sBFCviNtWxhq8gAkqiCFPQFlsoG9X4Pjdy+Z9sw6cCpWQ+
GxVFsXzXlVhPnV0NJGI52Zrkbcg/QMgj7QH9yUxD8jdosBictXidvE6wvCBuTvitmbcG6EqMRntU
HIL8VPTDQ9Th/+oN4o7yV1gS54JNQ28HdfEBUrncM/HVBEdGSAyiOekCKVzrL/3TU0CCj92Wh5w+
FX3Mhfc3cH74+xMShQnOdes3pc1uWGaRi2EBqTjmVJij2Dru50TIiLICa17i3yEGoi8I8YWThKib
WYIxQroEfh7DFTu5o/jSTERZwF2ok4ZT/pkrfUfv3ecq5wIydYrJipdn5jc/T2S/G1MaZPuDh7Qp
jtgsnfROmWV34D66CDzg0Rz3kxHVMik/fuEjnRanSdiMUEW0i/bd6SIvDG9jcXdBIWv613RFwxsz
1zcs9qcqm6uK4SCRiWsjFz3DObQFosTZmQKDKLKt5KWXoEIoc8aePSJMA7aFat/GO7+EGVi2DDox
eBYJiEyYtiknLHWRoClhw2CCLUkCICOyKhlDJkNFGlbIzpyCB2llY7xhzwFod6eTnVXmHLQxlHY1
1CDVyuCQUft5M79qVYePsLOzb3VZdhTbmWTyVD2P5uulrZDdDOo1d7sZ+s7YyRTWLKUopS+bOE+A
pqgdljpQ9Cx3xyUuEMTpJ/GWRJv6Wc4u4pWlcsd9zOZRcS/CMVgmpmC1oZFg5q/Y5fJ7jKr3Doqw
kobG8FUhjPrKxNnGuJxS9GStWkg5aYwncvMUJahfBMbqZcOQ92fEbj0/zbs/e4bULngm74DkvDQu
l3LSTPuLMcPN0/l1AmLuDhga+HmAd/EKAksxaC/zZ1YYsoUmdhYMaiSVDkQLC44oWG8Npcr3qaO+
UdpZaz9JyrsvscZvpsMU4RKUUT1YRK9vobKRUKRUwuLwpOQWxzOdxfPn+NIf4lk3wkk5i178F4Or
y36SgWOm+q/sVuqI+9Wq+/eMS8Uqvdbe2Va4gnF2nRq6N4e/bHSxi38ZwvNhxrFXkEGBGbkC+B1I
3gQ6YrwA6rylnox1DdZQtNPO0r8kUUj0UYhqKl4btMu1R4VBrKKztUkcMvIxHh9awSdsyW56oZRv
PwAg4uOZaHolCAYMqmn3tSbIQueBaZCPCF31IS5KjPSqHTmRgXp4EPkv5mDtRdifta8iisRRJp00
DFU9lwVyjbJV74RnDII+qICSERXIl8MEa8L29lXtdMahk3qRETo2V7F+DD6N3uQcMVw+TOEwZD8a
vK5ZtXHsTRt887zJhBO4TtRWtaAYWe2j3+//G8JfqTcWoCwQ59BjiMAiWelPhPMkE9lLBTyoHFJw
DrP1LZLoXgLwpchBZ/blnNaLFf4uhTiSgqm8MrRL8mlUgXtK3gB5iTh2wyG6pf8calsSz+ZtKGE0
cGVK9RlEzNQAGUNVHBSBi8c2yNoXhmTvP1WJD8+vU69UhrpvKPcsK1LH21dHBubX/0+Aj4FiRnU0
wlQi+/aOx9GV2buh2/xwxytDa/cqQFTFbt0tMHa+Zhmm5cqhzvpCZz2W4CK8+QNZR6+nxMuCzvt8
PGgIUrOR9060NWacUQSG9EFmdLvQP7GqM4N9PdkMXeJZhxTU95HBmCbxyroSHGP/k/tKvnm/sr/u
CLNF0plJXRDSYUbcGLwODWj0l/Sz+2xVTuQUDHlBZz/U+sJmN8mHTCF3oASdQ5t49DyGiRDyDTfp
QOiOIzcSZznhaGZnvwNoosHbfFK9lO7a0deQVxsewHp4kpoLNesnHnWu1R3p61bEVrKZbRQij+pP
ccfvudEHxJALaA5yKTQihaZhJifLJ0+OiDhW79M1we0X6GfxgSPfIyGomYW1dRRi2FeMbN0z2CEL
x3ODa1Uv+urJHAyKzeylYKHS7EH/Z5Vqd67guRHsMxnJvrp16zxsU1S9rHxxcgQZ40bs2J3M1acB
5IjbT5O/6wpi522hNBvcp2AH+JKIReUy7TmeKdlYb/wMMVpAAUqDJqwHAMx42hBFUcsgeJEJWl0T
Wzsa2c/JTg8smkrfSVlFjPiX5bSQoejJXfN36kz9hBe5qQGtvqeK3YpoH8xmRiIg73pXmj1tvnL0
FK1Fcv7WjNSim2tPgh/cMi1Eh1M+c9qcuQftgDyDlZIb7pY7OSaxG3spXNRJr79/WNWAIo1wUD1N
CkaShRy8ROUQ4bmZrJ9tZOp9iIpLzS2KfBx+uGRd/yL9RZNz9DOYvztQfja+ohZv+xgzdfKGU3xE
+q+RC3v706l6R0sN2ikimPy8C7m6o7bKUzTGHGUFBPHFUGcpEaK0TEcIY7OoOj0HDC37iELaCIzJ
Y5uJauXdsk/4JQJLa3eb+kb42Oq0qY3drw3+Ug84YPlFi9lAOrdKGcyMoteizG7NdXu69W1uHVGC
MG8NjpoCIaBIcTfrCD7i5dxgnC3NZjK7Vm6DVLO3t3OJnDGX1v2/W9ci+DXSXt2v+TTJOXlY1OaB
lpFrIgcfvHvmpYACpjX4drjT9V9bMpKMLmn7LVnzfGxHKW+/3QtljBMjowlm/+1QkAAiZwKf3i6T
ktZwMe22LE2mPiYlXk3VjdnTIJk2NwVzkFx78nsfMhHwnGTTjDBlHlxiKDYKMKtST0BFyXAcbf0w
fCoD7dsc9KvPhQIbVxAmHHdeMC/KJMH1JS5D+3Nltrio1AUPlDZTfxMUpTJgmySbyCI1RzxiMO5Z
M/p8DqFvgG5OR63ofCuk9KFWXHPpVvd0DeDZ1wlOtnWtj1YAIPDBuvTYxkA8HNFo034V1Pmgh0Xk
S0+5ULIEA47MLkxEGjBnEZrMEt6zKNs/5CU/WnSnriivDsJhiNSJpD1Hy4B0dX2RC417SoP3W33S
/rL2O9t8/B2pIPNt5z+Eeqv4pbNzdAg5pSJNOYWxh+FBZihCaBcfAP8cvNNbgJVjsYgDe3TQoxvN
Mst+vZuIs3mH+0aFcnk20YhQ5ZrcktXAQUfyT8xgI39o894djofjIvlUzW0pHBiBhU4xFwMqcD29
sIdgIQD/AJmWFs5Ft7occmMmCzcg2T0vy8CfodQi3T9DtBe/8/u5UJYBJeIcvRIieFzZL3WAf/jh
l/bsI8nf3cK9LvWztLqvjCncYSHk4m30v5wD4eqNz3CCIGn7wfIK1ox/HD5spnQFVALtEVoWhINv
k7KPo4eEcvzD+ORliu2d1hwW/SxTprg6E0m6wS95wDjFpPO/vOPijOHra98K9f8kGOU9ufDOLE7j
zq4d/u0bjsPmYXTn+gGfQ/10kv05tKxb7+F7jTDB5zG2z/Wb5ORkRHhWkl+EoOxe/z8JCkcZL6V4
hIFT25Y7C+dLFEX7EX47WLzBxZ+EO+bPTw8VK2NplEGZYYov7weitTzAQ+vWZAi/5mEOSZ2tbAHm
OJyZNIAHI2jIfqWQuvWwfmWuw9jbzzwHoHAlKgBWhjHAsi4GVp1XsmLCbUCvuljKA0WxlbIJUFee
Rw0yuRlZsm0QtePsYfS33Z/W9ZdDRVN9B9cP35m/YtnuNSWYpxT8pNxu6mknNDQqcDZRgkh3EdhM
iqa0ns4JPs+X6eMpbwq6coafGXZDI3slxmOIvlRH0XRAY62+T/rtVnb6QIqSIZsg0xCALyRmiXu/
s/vIocOOyBhGnpPeHLD2LzACxQvyJh6lkSxdHY0yaYEBa+nuzZP9pZFKhurJdVCbIL0QMWbjpKGq
pL9/MFWC4XT/3Y/4Y5QYALhULENNcgzQdH87cnJzXlbmmWU93l7rHbUXrJXCPtgal/alCgLxYxfg
LTp4XLZj8gglbXNuGa9qn1gJvDiSZJYGAJuJDUgd5CsCQAF6w5nJkfV3rLkgXtN1mCTZKgnv90qs
WDZ3ciI9etqdkK+ES4cMVE8K1Qvd8Y+HIGmDWrseHtKuXrldKFybUHc7kn3YJlaPelEDZ1Z1FPLa
6x4LfKzHYrSE1K91zigMgIjiCTjEeT+h2i7zmjJ1NecawgMjG5sZap9hsyRqFVVBV4Czj4EyA7nD
xDxh/MaZyYNElWjx1rz9ymYkuSV6D6qWFUsolyKUvoEd3m3GXyunQ/oiJM2oN9zUoCn/FZ74nXaE
Nl3Fik7lqWuaSMrLEleDa30FQdPl1Np6GrmvJCQjGSQd0z62D285JLWIcmi/KNu51tBfI58hond7
2aGnIy0WurucHy2KFphb7QymPoeF9iC6fhJyCFoakObHTbPAAlbgp0A4lDrn4l2TR7PjY1tMjpoO
Lp0DdPga7x6Rz+zghppJMgG0zEdTnNY0g7sNJlNDofieO9g4yVQ2KTonNamElfbfmRb3MsQc0sQw
Dva9jR6W53/7FkU7VIqoVuvKhqAtnbtjuKQkiPOWuTs7rGQFkH6KZVOggB2AisIgDon/IARu8fh7
ZTKL1tLg8cT4HIGm2ffohWkdNtIcqwN/UJDW9ZJr8mVmrTU9Xi+1rrVDMbq13pLpFgSjSjmZUMtF
NLWG2x6Qokn4OUewxn2b+buILSDJCGzEIuKc5OEsFWiSgVgj9oALpCy3Rrul/DRzwXLQDRZCBlv6
LT0atp5EY3OPfZUpv0H8BLypAoum+bGoi0qRM2hLO0z/3FxrY1kMOPjft/aNFnRMb+i4+4YbyLg4
u1HOF+VRdi3MP2sheStK/wa/EdtVUgvk1LnDLkvCwwJ23WbDxH35IhXS4EYBZrKQCpW69+ttEz4/
DVqku0cKCeabyTAyVrrdys9TH7TDMZWErABN8jKpCaWTA7vtZyG3F1cfMUg6Z1JHP/HWaWLpTZok
z53zqkvgzmLFGWTUejgixPn+Y9KFzgvA1WISxsBpVoBvSFv1GnfB5ehxrQoSbn9Ods87QE0Ft47J
SXQjP+K4Qo/SOsGmYep6d1fnVi06MvYIyYtKzWQmM+K2hPSWjePdtD+NopFODmBISavG001BQ3uc
WmZxIElg+CRppNYbUkKj14PtO4UsMkUTcBab2dU+lIwvebeDzVVbZvdoVkc2NesH229XfxLuL4ra
fiYsIo7gq54BHziXToI02Jx7dNYvfHYLYocZlEGJwTaFROfJHJhXfafGaMJKEyB3LcH6y5MXEg0T
HcYbIinWcNcjyePnAl34rShmAkDYvDzVkwDVYKuc6jdTYSHQDIAKn1CIgshO9m7IEfEB7SClr4qc
fUNIGGriF9otC8rh6DkbVfp9kU4duF3dCiywYNUTu0zXVFTxHlmTgQcngcYm464doj43wB4rfkbl
KX9lPn50K3jLQ4m+3eP/BMYsyL/Dttj1aAU+188P6h+3RxBrtCvUO4pTD2/7NcEAFHxG/HAPkple
QuPsrvWB/1YNFywM4NTf60qMrB/AGl1F1bpXoNIIPSUUorffIfcpVAfn7NvSVpCx3UoTuA2C9W+s
PVbqfs1P5MIgxXS4vxX0d0+qV/uxWjZEwmDmtdanalh4qqa/31py2rezQ6SG6C/cEf0L8vcJgjau
viWJmtVHdiGgiIV3HVMOdxHnLH3M+d1XQfvPwHe7okLqZHFqX4NJH6LLh5Kk7y/T82Hiy7b3jxsR
kNqhGxQWU/wJsYtgIsHp6sJYf4iE+T5yovWTi+ECm7d1Kn3P7uuy0aqFYxrS2Uhdq2VejF4dc6mH
d8/sF10B3EgCBOKi4tNISS3VHJ8gDMg1B334BI6eQHqXtQ6WnfasKur0Jo9tS4FhBaJE1C7XSr2c
1aQ5brwXAaossnu1u+Q/ABn3ymz1IR3WMkatZHXLGx1Bf3fIdSbykRHreH6PYSdAH0ZiSk/izXpL
67A8lTQAQd7wbyl3uJfSgf2uXgR71cvqlYprJZcLXRd3QZrHPi/rafFvx/il+KVDVy28YfIA8FxK
4Op4C+0OykSNQ6CCbi/r6jI5EacBf9Weu0NCqCh7Yf2wttkt2XqN2R/AQhx6g7ZY6MujQoIFGiH/
Xeyp8FoXLOYJsu+Hu6n2y8N2sMv+4hkQllIvuPFrSwYLnXoFUeiggUGNFzAtBMo8DXk560FELMcy
UI3LjHYlkwaROahqOmlXys0c6evNaJx4A85UoURC+c1rh8/Kpx8IeEDcYzh5Pp285avZyEKI3+xG
mt/HpWB3lbnQESsDM8qWQ/0FZjNYq+QnmU3czH/ceOJ8bEroDgpiqdBYFTWUPWer0eWMPkZyQrO6
+Mo4JsY1X+xYFoPkCv1FOip2jeQ2SzLWejvmpBI+tnAupCv2YSYwyvRs/BNJpiRcYCMHjWqjd+gB
Y/K9eI7nEm5U1QoFtDemYp3rXzj34Sx7go3nyH66X6yiAM/ghISxwLiWgFOjiJVTpX8T9P9WP63Z
5ccGsERRAy/ubSbYqa7F1LysKkZo8n5WGkBe6o/c5UfEQbZEB2pGlId/bZ8+rbZ3ctrg6Wi58vUb
Xk3tFvrQfjzkRHLwpO021bhWFCOgf88+uuT7cW9KbOIxdU3f500LwG3p/Zoii1ZeP7GIQW05Th0j
KchjzD8sB68CBuUdlJHwhu9W6f59gHNylFJmQAZEEkxYdJV1L7c2Rzcnt4dTV1FNrYG2dd+MornE
ynf8Ss45rnU2b1HarRw33f5jVqo+7BkmvEh1bhgMeznZUPCN9lnv/sKeBJ8AsM/H4puUML9sol7V
57EmaG4tSdUChEmFtWQ7AF9cA3MhJIievp2DTMjYKEpa2J3A5GHecPH97NofBxjfxgA3ulJLdIA7
1ecpS6BoMHx+n2FYQxcD5RuUR3x6itS7MdElibdhM6rY6dNE2Bv7MCTIVM4gxSig1TttDZ63K1Yw
1uYahRvOCVp6K95yZwfSCXIkQqffEbnkchujOVleEamolvqK/G+IzNxQOj+jdykoMfSfm+ENYKLQ
z+x3O4pm5/KR2Cy/zpcsQxTEU7wIzDNbSE1Q2O/7IlY3DgaaYJ/ZyKsfJC7M+z6Nk6G1FQ1TWEH/
OCxP1Nk9xppF17zkYRappD3NcwoyOZTtoMNMcyF0XAoBxRpObKxU83ELY+v83/0ueUs+jHLsIbQS
4h3PT/XcsWQwKJW5KMKiCNlCljEesxFrPr5tq1UnCA7UJou056SlEEUXK8KltJ3mtWGH+wvmHtU2
WprSVdXMPREmgQM7MlynNI7+f92Odxnl/DzkfH/dJ34J/ApFJvGYestPYc/QiXscq7QmYw8VvtEx
JVMSNomS3gve+55sh2fD6ANOvwE6W4vrbbr42jfLnkfN4lXNeTuwlOVisavBcDNdJMobjfDll9xQ
oeN37tGw/7AE0jz9rZW2D3F98HdSHdBeKGyP74yFBBXlQNFAuRrM37i1NAnGDv0LHcPHtAMN9Ow9
p9g9uWcE8kTcMXyLzldaIXTXpMN0OMdetkIqxVbFQjRJ8sMDJCp5727lTFNylm5EzvelQeUsXRkW
9+CqOnF8pjMPcQsFAniKGKPiDsn0JRtw4LRVhd/o6yKg5flXqfo/paG9rAZ0uGREWcXlJVnMRT14
ikBnoqc++HaXCIxBt/hokLrl58oa+7Fe3yUX6itM7xu46mUY6QJ/YE72WZH6FUlLZvjmUb1kLYpZ
VfYA3FscPJwv2z1/Ol0t4QtMz6CnrHeu6SzoET2cmJ1J9OwvYhCWXeJTPHc0ZgYe4kQS8tl5imDP
WcO8/jGD+vpYIe8iLe7HJz3js/U2A1nbeD3vNj9RcgGjGWpdzd22cZtbvMDWBo9xZZTY7cBsj6DB
epeqvcIhcXaAcUtqkZjoNpZOhhGm+Aejui9dDR9PwcNc1Ft4VuKEz6TEO+ZDH3MesFA/E6gSZad3
qxs9jEDquyxmv+db4KpCMrGf6OCW/nKxUH5RdsdMzBGEzl8SBfrxXJqLqQWe4Y5x9xrgKoKDDh2+
qnP80bDM/mjQZvSb7i29zsqXZRrWjFjVknpIxuMqGnvlMm/OIT+yxiF9ajf7DUL65HD7stdO2z7E
C/cmTVCk3wPdjQH+ykdaIM2zeLENpXkEueEQLjphz/KcwJrtgJPcG/j4PO3ejCBbtu7ABqsgIPNL
CulZ9nMYtINUhC2nvWjlt+GzmFv5c13KFVNy7zisVw/iKOZwuDwJtxOg16B/F5lqihLZkUludIoi
bZkUz4AZqmitzgqCKRgCj49vitHTEY/R4jfiSny+EAw0hJT+FDl/+Dqlm/hHDwsG0iCMArKF8oHi
xCfpK2GxliIvAVIJ+3X7p46D2EsMyPlI25lKjEJpkVLvLB0R0EZ4EOjV9uLgcG6/3PnK4LNDHRpM
LqKiFhlnKLae1KrTGjXaIEdORYPtABUzJau+zvCxrSjVDK/KOqudDHrtvGPhR5SD2NkIa4YSJEJH
3hj2v8vL+Du+YZTnQgUZlClB4BtfX2cq4hc3EyJaPiEVtJzjxvlvbe6ZjofUk0ld2D22ZudOtpqt
aarZ/9JbKzT5nPqrA/eJaIM8YdlykSMZWHXugnH+WjfA4ip90vpXvXJPA9ghxsENSBkPKWfYMwv6
Ar6RFUqiF03HEfKlgf4HBweiZOYD7RsUs2NqqrRHNrKVeYj42J7/Mngos5UzvsSxGCAw2HNV0z+e
8YzROy9DA76S+pbdkqMC1Jb+HPG6JDsvlQ0ZwWwBhgSi/UfMgzeQ2bXh0oU3sAC6rJDnn3Qb9Qb1
OFh2ZlQMBKEdS3nE7zD4Cbd4xoKhSaGEmZvVbmjLMI1c347k/gGWV255kEXsBUiVAi/jIHFh6E3I
UA/0cX2en0hqKAo7vc2JggQyRQ6CW13oHkcHAYCdcihm+VcFQYMEVJAK9VcTOm93UAUvC2jffea/
6IzFyauRJ1J58WO5DFQHBtqtCnVpvg3hWjDSGelUeItBn6owCEXL/WyMb+Tdpmt5kWT8D41VaLrH
uhneAiGs+15scgqtgRms0ypqhtFzzpuvvVIkN2A42Ic++h3sap21xRoIzmlev3/4kd56fH9TMqTk
VG/GPTEPcIv8wbpCKJkyzp5hdSK/waOPAqLAVOl0WKoTaNzcI9ToQDRhzYU8kY2bnwccwtPYT43I
mg3Th9rKqHJVUiq3rbGSsCdABuEI7AEQgAcId7/c+GNPo1tdhSgZTaZeguEd2acI1E59mAlw7FLp
H+Uz0FuvnCux1bOIJHVocXBqM20WvhDa6nZrkzicoDb3AjQkSxgYHLn8AfpUjIOXMfGchkYKNMRf
KEa/y5owB38AdavsCRKMPiNIamPuTCzbC9htiNNKdf5XDRvtZyA9QnrHj00sApKQ1yhmAIvCJwZk
7EgH81WUTRuDBrL4qikhj2OTi4Rob1n8qXGOcbk3bV5IK04xHo7Ln9gMHnBK9kZGNENHYxmHRknh
pUq8JhEaeK6P+jDNaGw4X7DiNivwINu4sojlc2wTQpaznSg9+fq/sE9Y2d9xaa8YuTPsjKuBG9NF
EMmWdC/IGZOKpTcsRuQbtKqIpVSsQ/oTt2xNW+xynW0iJpNVzKv2xBSkLNQLF2A4T0I6Cv0J3gvQ
RER29wDB/Db5MosKdcaYH9/dQXlgr4+XreycEG7f0wZeyg37bKTWCuJdL5oaXAWCxJLGqP63K2po
1gqGlH+h3bM8gA/kDeDNxZpEOx4LwWHWNqzMenZAFz+GX+LYOYFJz3GoOlI8dIgeLFeEEm4CAzPu
u+LTTtKgjPMOjvFSvUNLVQ4DFcTBqyaZS/hNkOlAWdyvpKKEQxrJnLOY4UvQ9yh9yIbm/eJ44uvJ
pSAYFM395BGkr4/YcuzFVavFW/eZmba+RnZS0fGtsDQb/k3hiTYNPYimxobJ4ZePtIlcEj8uuCBN
csTG+S4afELBscVrQMqh3TO1qFnE07gIrbqup9W36PF4G81yp3nebpxWjpUZtnhKdP8y6aEGpfGZ
S58N4GjyQkdFyClaG0ecmgUTausMcFLHKhKdH1IyeRnOymxWsevc6Z3uaDuBMNUMAjbhH3omvBKk
tUZeBteCdZQYQqQlIz863KJCC4WMAAInfxnVSZldqcOfev6gIGFbm+AcmeRpCWnNRNsxySSHwRWI
Dd25IKesjBkT55cAjQymTTVq2sJUHo4kbMQCr6C2kzyZAsvUszTsGXQek+MNOCeQD9btLmmaX0OL
c1zV8lqx9uBflEeiiwp8814D3y6lrYEkuqGtoja79dZyQVvgD4pzVCCITNZpx/dkIySs7Ye7qqnN
qzceM/5+Ejr1AerUG4qP5OTuWnZAYFMacbdgj34WnKQCtWm9n+JTW8L1lVEV/5tJH/sx65OGDp8P
Izhp2AXOZ/wqGA6Z4tkoFzMOhFMJtrT2yQ6AJflKRol84oN8ikjnnbxa+8usrvB/UpoLi8PJ/IYJ
4lSiZAOK8N50A9iRZZtKIUZV7/AXAPkW/UH+OEIwFJVc9/3tY2yH8rrdp5/yR0FIe6N3js8Casct
5hZpFQaRXdTs7lxzTGhEYMjCBzkRlAQypU2GytkXTWTsIAtGhbJdnFVsLfhQ5/ySuZhAaTPfvJ1l
yo/vj82PlQqWstkcLtOyA32oqQKpV2kzRS5gU/Sd2mJSGYTbz30AIuCPxtdh4mx4jJUKaVPHnpYa
oyTq4kR/ixj9u+7NtlPt7HDcGhrhhPjJW5YYQArKnFzOQvuzACQZBUuXQy9BnzJQoGE/tHaAJwi7
897FzzT7uwLcL2he93iqVDdRU8ptt76u6ur66ALZYg+aAFFLbrojRY254O6NNUtubQN4pIRZvs8e
kSdSA09bAEiXvQawzfu6OfJyLaBb+cEMNV2hVviHTSoKWiQ1XiInVOwXdQMEbVor4m7YRYAotrU5
Ly3KWSNcN+NeZsT3sAKS1I9zJUYxClLDwSfZ5idro0CSZK8KIOf+u4IYFVddTDzwLHcY1ZQnDitv
+3k6nT+hBMH8Pyb4UdjD3PCOOK1MM1yCE6DlpHjw5udM7mhX+cXlIXwFOosmoVK8U1Bjvqx+2NQG
AJymoQ9t/+4VChH+L3ea/PiFsAfQMoFEcnsI/C75LOMrv4kDj5Qbbq77/pAzN8YMqrw0FiIUaQcJ
QhnWNMeeOyFiDWPEg/k24/17kzBIZUZCu+ULABIFicA+YQga6NfqkpgA66BmYUbmnVGZRNGiDDO1
dJhjxP+zVOiB/vVIKYvkQ2wfaRMDOEVO7D6CWlRCUK2fzxkMyMoGfLV9wOD5W+NVLhP5Kei0Agl0
W73tBifhfmX2eOvv1woOYWWeujUPhP1sX5KAR3b4qzDTbgwsyTB5E9/O28m6NdS+6iNNlUE7BXSQ
YdVWNJDpcn9J8e2kQAfVTliwfn7CkMyP64fQGpyVjWaF5JvUVhPiQw+Ttp1w1O5073ujJ+SCmWn/
IpxugnmAQNkKUAe3JOejL192poZLNz/er/iwY60m3rGi1CNAGZlP97EzvXD0TVruDtzN76dhcngx
Ss8wC9AB1oq/EZMzjQGrmK+sO8U1nL74lDOi33t7wq8QB55l1P6P2++kBYT+ZL4jsv6Q78Whh5RB
Ih3baC7+bas0fHAtGMLGkUdH4f5YsJAEVuiKy3LqIvwJkrBVNsWFnDhN7ISLln80YrnJahLulHFs
zeZDiSe/UxrBrIq6hyVDgW0pI2llR6MlERPhZuGD2tp98H1W/OY2eN4U45Z9QiExaLHl4kTUBdHF
KrZWflKbcir56DpPWL+MWDmcKGOGKwQy2lKt0P1XAu4bLnRMWU5Ed9Wei5kVDaMISgIoSOKzBMCA
Utu795g3LU//ND9FwC9GC8TObBGSr9KaS+c5lcI0lIlhAvdy0xlkclAc6l4YBihXKVg+ErRBOeKM
PIZQZcnZTAnJYwupejG8PGMx0ny8hvvTUWjw8f+vdDZwR274ZAwXzBt2kWT4/naPEFM24ySVVGGL
DVBrueCQ8Q1DKfTtqzXceJVgDCJsRtpQu4UP1iw/wYDju5AFfTqW05c2FjcxM4kpIKQcExWcKP0E
AoFsCzUF1hn2QIsW6+vaBqgNShce0/Zw9fuuxDspCfkggkUfKDQeTXXWOFSA7Uhcy/FlKcbFK/Yk
pe9QubG3tIKtLYNQwHg4x+wCSyqvWut+wX9g+USwylu2Vknvn6H5ucOM/2Ttmv7PK+FAqv3qUkfW
AWZiHjUC+XJ1CYsqddUQ5M0V0ifsioCjgcuJAr1VButNiPFB3Eli4Zj2OUm48II2CNlAXWPQjs2x
Z0pyZkdQpoIHHLbRQQ9fanP7t/tHL7MWgeXvVrISmXD+ilsPQNhOA4Xgt3X7T3QAo8DIsmi4/ybc
XI7CfycwST3i1doone507xemWVrBV+ctN/SivayNOsPIpevo/Lsx1fFPsLKiZzoYUxmjl7vYYXD+
bcZaRET/2c7mY7ur3lnC4m+AMDOQk4TBYn3MwJaY2MWmWCP9B1/ivAvanF+QdLXnIqTKdFyunOSx
M5/WHntiwNR4yjjRQIlE8elfaDnpt7JJgL6VPbMOeoc5950xyLDGr5IcRft//QTf2AqF7fUCcG59
AuSlrhiaAnECuMj8O/xvmU1QP/vm3H36Cp3hameLTaTUPsdrgtKkj8OM3L4SLV93kM5AJ4FMZMYJ
WUsxrOqVR6h1gcS9X8pJRWqBfpWau26jt15Gsm2jt6rnnLceucL2O3GMoawPYITmfExFEAobfFCe
no1FT7IrzN/kGnIVTqn457ZmCwTzgAH0isMz1s7/PxfCM6xwWPsceDH7dpwXoM2g9ayjYYuhySRj
3PXKxh82jgzq2xm+p0MCU/jIEDeKI4wBWDZBXAEWFRNkzrBImtk991a576EgE9dV0Q6Je8AmLn22
5TPXHQsstwM+uAq1zBZxV0F46R4RBEFDZWAuHGs59wQOUGpKdK70sdTcJyXEK4GNWYzHBsCmInPH
bnu1VOSgRk8iEjZf767f5LBXzKIIDmmw6/1St9E0bvTPzaU+eahJadzxoBwwrbrtB6nkG5qNvPjm
YPzUykuiH6KM2NZwfL0jH7lo46cjzHx7cxAEGBRfioEfd4/6FLxl2JvR7emDHO0vpqlCjz35yJ0e
OVc3dphirO4i6hYPgL7ul3p4gzGvHrGr+L6XQa43PMPfz0LgCvQK8wz1Tzs57uHYxkScit/2UWPI
tlXUsCOsKQLVbChF7EIG8CFQhsd4LpGZfzWNqLpni7ZeTjWVX6r+LmE+Q7PYIFk/WWmNdOEDPCGb
lEo1zlVNYTQHKdP2IVkcDUisZcSOOQN9gqVZuUj4AZd0FhEE/FMp5jwpFo10torG1bTzKKCUApIJ
zF1CtmBQT0dhClYt3IT8EG/2zwiBFO6sDYaUARXIV/mTk7qCTGV1WXs04LzNdQhewkrLjdU3bpjB
5fk8SUgOV7XvlAt/wqVh3rTg2VSfhBmGWPufXnDBaAZLwnt6F/m1S4R/KCjkd2Ct6wY+XlEG78dN
xDsyJMR9crj5QblhDjAVgjRMXXiT6xhc4wpVQgeEpbiiwrQ0An6OMdGg9cHqHDJc7y4Sb2p9K0ge
7kJtgdbrQN4vyIX/Pm7/HtfF+vJW/JBOORDVwaUfagLcOX3PUj74QPtuhkJ621Y7JoCaza5hnwjf
9Ewnql47tJ3/ZJ3sNXrt1nadH52VKgaG4utJes+f0jdThb6yI/Vd2xBzPsxutVcQGq0P15xiQEqd
OLer04bfKNI4wQ1nXZkbZ7X8ElnPGW1Lk+BUlebspu+8pRrmL22NudBaVrbddbShnevlwfXJEq8X
u200QZjAKtD4azW9YLSGy8jHg1k8W3iH3rXsvpUWlHPzCyosTNv2x8S4xgtUNetxWSTozqtzQI/q
EBpDcKsY6QFsZpXSyFlJfxvCoKprCkj6iibTmjwIOVZjnLcCk7v3XG8PfvxyG6/oGETLTBMufHiB
qmQ4sQeAqqP4NkC9eTSVLjSPCqQm7Tf6PywePPUnRxaLRfQZk95nc8cXm5UGbC95iR2hlA4PpuRq
ET/hi9nuLE95CvOf5cEnC3yf5wKiNdyxR0mxnCosEJRALeyB4S+FxIE0jfsA9VUS17CSEY2ae2HI
dBwg+jM4Jpcxjrw8ud+/IVlz0U2/kLrQvcBypylo4YogFoX9rI79G0DXlRImnWAC5jBI4qpP8yuL
Vp/XcCmJPj4BVhiR+P52xH7hlD9q6Qx5igr92ZF77Ypo88FAcXyd/DI7KIeD9uQoJdZA4OiLR+FW
GZp6gzfo2OLJHRlIV+wBKBLLggfKSrfkkXj/MqDmvmIZw+UWlQ3piVrbvqpqsE6qR5DRlNs5t4Y7
lJwNnfLwhhLEPikdJ9c+u+Iusk/YmjwD+XGn7TVzSEtt9OhA8rcnF6nNUbxHIz+/9MgyQGW+nHNC
j3dR3opEPAj2RChb/wT1hsT2QB9WjuNvHqCx3YFwUwY1i9EMc/szgNmsDLqBilxu6IP6nM/yU11k
BaHlznOwcpKKqONwJ9vLpyn8wOfGZNxWINd4kYnOtcVi82DqmokJWE7hF5Wqbs6A8Ayk7lPHxYHZ
jiOX3KQjCx+Ra1nEBA6H+/UsMNFosbv2mr51EPX0R8rJSTz/sTENsPopmlOvPfNrdEKfBBHjFO1t
is40sowcYN8R28oiSsCsp1Jxuv/fWt+1fkQ6gj6QwJeRRYDAFU0FUXZOQMwLnp02H9D76u8razuJ
RkKuVvjpbJlr2p/vBTJIIODE3w2v+FBOSREeT4fpY6IaKtbcm+OVUurWk+iN8mAz2P5WPkML/Tvm
h5FvX50rEYvfJHP8Fz0PuoRFNWCxkC6+CUfB/aR0K1C9wbOv6mZGt9Z+GP4wB+9hKwATSGgfKloF
gFoGK6wCgxfcopS3WIw7qI3ctBTTIzA9T62ES42dbS1JaV9kd850WVNeK12rHUwG1j8JJfGd/iQb
XqEXgbXW7a+czDQQkJ2peoWkDlfEbcR1YlMjcMFAFHgqWK7ss7Egmu/seOhGPxfFvYyu/RISa0MB
oMtXIKbPepy0+EHKt4VwkK9cKJ74xDfa25BLWIG6LINHPA4IzSi1+tyvvCY5WueSdYNaVlgYp+Jy
R/dLrdc+DdnLR1vQF5RuMp9IgDvXWW+52xj7MyIbxPTjv7T7+kMmeq2wd0FxDSJ49XGYENxsQOQN
yXn8UrM7jgOWV1AgSNRwAJSybNTq6HB7EHRl4fLieUVPREfDtP3szAKjbq9GuixXYeAfX3K4i7ye
TQ5gc73xVCaFuU9fmxLYkEbkSxFbllpdw/O3fukzAIPr2qoFRdY6JP25K8LezLTbfgouuO5TN9Zi
UBwvv8vpB4uUL9zi4cEq0UEQXWeInzxpQm4Vsf55RfRtKXO+yH1Vyr2aRfb2hpGCdTx2kJ82QR5G
EAkxCsSKDtFhR1i8bHwOKOtv03m8mhflzCnFCO+DEy8ebk7EJrAnoslw6DC6PBzyth4JkfpxWyfh
GAyInKXEkImKdVIjjDDA3reFJL9VFU5UcSnVHaxnEFVrGssg0SEppY5wY9JMxOtXlJsX0M9HdhsC
UR1FZofXWgrQhyQvqiDW378qi9Ebdj+2Kb4iGo8zmkhqPlEi2ASkmfmHi5l+DRvzSgwQsyxKwaaV
utHAQdAzdrc8lcTGdtBK2ZVjg7DeREnMwrDwVRwEPjEbhm8q8LHuywvi4YqJHKklVuAQjWieeCrY
DMCx4vM69erR/5kuZzJbB8CRU1HLEjSlReePxmxHsOxAf7HeODuSp+5k8NAi8/EtkpZ8Rz/LBpQl
lZzSxjMcIYaNGEQEjJabiJMa4JB3QOHFqMslVON3TuclLDbX5ecvEbWBVFakKljNEPYJ4mxbRlam
lObqDJldiDkS9Djletl81W79nKOTZw6hFGhYp3wcC6uE/kg06g9a+5WE2vvt8xIbcoP/Swc75w6m
wh6EQxY8j4lY1gM49nt/3fakEw0S6L044jxCo8z7QdFKVD9VNbtrVDePs7vgBxdn+Mw83KxyaNS5
rg0xqr7OjWYBpNkDAQf6p2C+9zF3C+KJtwaqg4q/6LYFkBTDmsREd2gZCjw9xRqm5FterLl3JAZw
nJgRynEQnM4wN31O1UVHrbpGO13M45N7q9pfJdJadZpgPmiXqB5lOuKNKxWv8fzRvvsSejRf7mvu
n7jg3aQ/UMl6jjL5jrJQtWV6AGOZ64P1V70Y6Y3lzUvb/iL8Owp4BV8mph1OALcutrZWL6RRsX4h
VhvAez6aBEs8rXaeWdjH272nLX8BE4EJIjsOW5VyygpXhK/nKoxhbWruzGFNWvY5jovxDAeM9Nvf
iqL/OH6FjVlJ+RvOXfUBSX3LSdArRkehwJHBvxDLhmhrhOUqfm2nGTkVDCsmHKNLnzx+NORiIHR9
1086zUJtXDN1n2961i/9y9lIhcQ8Gp418qRwi6NkT+R0Ldz5sI1FPma2fxvFPeY2wsM/OKTQfaxZ
AWPX3znbOMU7dz/66dJvLohX6yvcgolSTupRerNZrBKvqrnjtmhZTkj/bl5T95QOwmRU5IoMrgca
Zf8ko1Kf5a7aWfAMLYKM74hPtfGmIncrewX9Uy8b/ZeytTQCLhV0kM/wQPDOV41msI3RBXqMeUie
cnezZsMu24VoK+MYxEYmF8xBGjpW54/R9kRRKJ2GDE4E/lq/Wi+d3ad8vXUm2ejrEGbGkqHrQ2N4
1N30bbgNwj1fMIdCaac9NJIcZwz8TUEJ/TZw+hk8cve7LtoUsGet3KIG6+yNWDMLJvtzRnStpvvd
thE5dA7oKvA5TM6ROsiNTAishfK0QgMeMDgacpD+BkSCIqnBp05qJXzfeUb7+PokSzQ5085SypA5
6IOWiCsDgoLC3XixXIyEmLPyn08a76u8edWfEA4agrTsGkKKlL0NViCTMqNTSAEVt4Ob6tVTvzRk
hfWFe2JXoyovgcosOZCS52xFrqLlQywTs0fPvZETOPU0TzOYc2uuZNbiUAKQhSejuKJx3qHvYhkt
W1vhIgOI9pMD6WB+Joiruiig8AYk8Jtj46GMxaxWdYWOxq3zhBk6ayfdaVcdD7uLWDj7crz8d6MO
OItCRm/htECv7NFWCXK9oTP7XzydfbAkfietVMJdE8xxHsqBr8lcloD8+dgdk5VkWhEdej0LB8Kz
Ull95M54w/zooxzVt51XhE0kMyz3Lzt1ZcF98nMgk/bMDRPbzuWwhn+0hKHMgAri9Uxh45vqxI90
VM3PMzBC4nKWZBOOeN4BZOTM8NQ98y58Ex2l6BnChKpqytyQO/VFvaqdPUGkb0if18eayRrVdZ08
yJUgq31pD7qtkSeDws2dA5I2Jvt5DW1Xl+scmAWlXT+agE7dLOt3b6QQwZYMqSZd0so31DEYvFZr
9cyNJ5hFhS1srh46ouSLoaMmdJ/e4wMzSp8bQ4x2BPoufof8zgtjUIu6hWvX5PxiMOGmjfn88oET
mpecrwn8TaIAnSXWyb39ArUGJyiB/AgMjjzOKIKRbXK05ZwcQaffae0D0f2LwPQ8QrY8dlOhv51s
0Vw9TioQVquSJLKiBgJ2v+1f/NG3PZ+M/6eM79yg+Htk7rEUoskx8OQcv17em1d/1zSE0LdWzZvv
MuRJhxtFjiXhy69bk/iVO7Kgrzvw0MJc5uE1SU3gq8tgBkz9OiAC6lZt+oNgdWJeDC3x7pdFvSyX
ISf+KhldmSOWESA0Rro1u2U0USyuHChHNVnffcYBeIDBm6hb9noLuNDxb+OvzDe+orU4n9R6QRlx
AQjTZObR2G5OssAfgrCs8fHD+dUDoLyO4XGrP1Q3ONCE3bE5EqZhn9DThkU8ZH//T4MiudPAuRGW
lyrczDJqwCRxPIErIciAgwFY+SjZ2Y379Y1G2q2iaaRJAar4No1FfMhHI4BJgtEZyBudguvcV/J7
HlXFDvXX2+JgGmLeLcE+TkONp8M2sngpEfECafI2J9SdOor5MtLg77M/l9pXUU8i1IpoMuIwpoBU
XPzvy/W0S3v8jq8lTCmaH7hlnrsfOG0iN7hK28INzbXIdbe/rJWiQTjAZk6ayVAnkSQUiVywQ/wo
v2WFmc23ygCzALXm9A4lJhyYWizmHiGAESLtvnbN5dI1/RTOfH5+3MveiX4msPo5aBFCbjX5tiku
0eprpnU6And2vk30v1bjWAgbef0I7rUYMcI1bvy3XHsHealbOvq0nbQ7XI0ZupBT+LvixfEyI9xx
X5upGxmMb5OXJOWZPn75109L9i0Fymtzls9u6jp+rAZ5b8XTGA9aAg80ly2c7zRQMJz7ki371VTT
AyK5Tm07byP2ZRrYuw2V8+D6Pl10AcVpBvIQPSIsHQyIWfKXbMP4BGn26ZmeVo3ZkdZOVyA8ZTy6
O5Fv1qKA4xnaTVTdxII3NF6ALPrko77rDzPXpxxqoX/Zf7WSSg99SE6besHYGoNsubbdV+5L+r3E
cbbZIdia5cVF1Zzzj0RPZF9C9857+ESS4nd2Zb0/IAZCcjmUumh8WnCIyF6gOgz/Rg+8yMZFavnT
3//Sgga6/IfUy3KKKIt1NxVaBYyv7Uaiiof9dNyzmuDTXNJf46dL017LcGY8fNMsP6ZP4qvoqTuf
ceRGT4/JvNyp14aIfbBNEjJgZpf9jNCGFyp2K3IXgbGCPscW6n6fPaK3fUxGyeWWvgS3BUY+YDXu
G2GdFIqHs7wfL+uogAPf/UqLSsV5G89zSvrsQjoxGyAs0NKvRETZf9v0OKtUZFfbnZ15tuh+14n+
agjMq+qgtQbvkN9FTscsoo/i+BL7vplMkfTwTLR9j0exznoQL0rBswbcCMd8YD9nF0iDiegfNkbp
yaR+70elLUWj3jlnUSNGr7uNz7glD2S2BY7EqjBz+E9OYiOB2KM3p2KzWF1Bi4INcTXxv30JmUIQ
1RherRqjACMavLKv7A/PPENMpKSJfN1LEIJlGiHIuoUJV5K8NKXcuMUjy41NblhOGUcJQI4kqFzI
fzz8J91rYlO87uibHRvW/UhQLTgvFMSHEfnaxADoOg5vgEvLFU8jJzPXxCfywAIf3AbgbJz0lLP+
t832J4f6cwev27C+yxfakXA3/8N4tHq7pKgdPLejRO1WR9syVjQCOhPVNzmozRftajZtpNlHrY0R
fIe/n+22KZkZu/nJvEPlyKbXwX00Fn4DvDCB3FdvboQgPh9vUmlKZ9BSitTPJd7hMwaQ3TS/3dMe
JCcID8LbpPP8kcSX/Xd5mflEcpZMmD13P8sY9lcf7IeByHIVNzJncqbKfqX6UtnIAZCgMzNB380k
Qk3dHatYcC0K6SMKibFpVCCO2dWn6Nxxeey43peQx9qvZx+ZvoGd9LMRaosH4N3MLBSMyzaEu6Ep
ZT/v5R+D0vgWK+8PwNrWZIn9tYA9bBU/xSp+6jKxT+GLp9Nz/elycYZmAP96DeX9RnjEf0VsJJmg
OIec6nZZ92bDbRNk2wfKo/6Lx3XYADfY1o7azuqXUfCb1Mesc0kZRWwqc0M18r8Lh8K1RGA2HrGX
vZ1CiavpnYgvzixoJybn6RsAX72mHFp0/ld4VueD46QLj31VUKnVbM7IIwrwgg9DFbW3VdqmOE0p
RGqPmXjYYSIzcahsTxtNQ0DOjHF0f2G0wt0W4nJxvKlXBEIHgrl/k2AbGUA0aKVW6wtxK+hHhVCd
hfKbW8qkJBCP1vd96K0703kDO13DR0ZnBiqEVv1zQs/+uD9LxXmcaxqTF9VVC0AVTco8a8N5GAr5
5PMmz7/D+SLMcLV6/QxYOFb77UxBqXL/jCvb5yjAV/omvk3sLBCHac1ArkRwdYpIJxbxW7m/geKx
AU/FufZfgUX1ssaX19hvqxjbTU885Az2tmIOi5j3xaM7yUNAUYv8Rpw08f0BVyBGevEfywKb7Xo7
Mho5z22md2IlKcp+mKO2z6fQxTHc3TdhfeddXrU2feBy6jToYb22RhT+RdyqhDCKwGE0R6nODlEk
ogXQ508cSObTOp39jTUVAj0TtpmHD8MQ1WQy7/hMYfHppqS0kT45/0odmc65kJFzUEqylzYsPYm/
lH5pQKUXl9Gn+ldNUnuk0YbRCH79KzKSEQPpEoCQlzPhwNMRn4WSQySJfXG3zEDVD6yXCYFqkcT/
Y5bByqiYJNs2KR+EY18rzIu5kENAg6IPNkqJCZyF2uDAau2BiSINfXhFGh6GrLCnRkH+Uha8rZIp
UgftcU6IE9+c34SKa72ikEsV4Ieh8Up5NiZY++GiGS17JwDIh1yOdbj1Vvp1JrWgf76gRvJt0lv4
spvpp3AnrYQHxjbJPhQBfxxmjRQb8s9Jl4pknr89k9geCIyBAiy7+eL/WoZAf/PwaF3n7pX/UzmC
M4+J6qti3raenMkdt7LlIT5dwJvpZ+M83C13IIiH2oM3ZqZhkcxt+yf6ngjhq/mBxD7UD+McQaf/
XkFWu+7XgiDxXE9izSNTxxPnfgHu+Cq75TS2J+s10n+g/Dk1hw+vFx7Rlo8MiSrbx/yg+Tim+h14
F+m9kNARpPS5k1f54a1j3+JzcHBsdQWxQQO/7CvDkSsh3twt3Ba7957ogaSUh5yTnEk6LYFM0INw
pvODmGLSoqb5wDnVy7PIlQG4DBljRNXHjrJwMC4CgHajpiRzXlxNayAulrrcQRDOTBRBsLwDdq46
h1GjnIHsgyCSgyuaO4sy1YTLUJZhGFMfwa/Hec8H58PAUgmgEFKiyWFEAoqxmRuq34D8w5R9VKCw
+bcQay17NxZKZ0gcqrbsCAuWrhYXsIK3N5syzrPaj9JXiD1valZGfPdhCUv2HcEmwiSRW8BA0lPX
z77I9miGtBBeg75mYxnrWn5fft22PbCNmN8j6aoZJ4m3mwEKmOR/t8t1tQmjOfSzKf8UwSe4qW7i
hhjEKDgDsB6aX3HQ7GtxOnu09RuQNeLZng6KZNd4lPPHtQRIxk1gP5jkQnZHQszUy8YQIRl1eiLv
hkBfp3Og9wy5SmEYqd04T19+WGtBkswo2/JgzubCoGjZ1Up7t3LJ+iABof7LNTOWknaZZERk1dDD
p+I+uyZyx7eqEQjrD3v0bOybnl1eelwEs2lJzi1cqclqvFSWzjBzO1jEcvr2DsUYqHAA1TCRPYBB
7eUI+WEa+HDUaWZ4xy3HfEP9GMHPAcb6TBovrwzCuvHTSEBPGagYRZtr1PSFh7HRNpJj4iU3rsgX
0JpcGjO/HeUNalO98HtHIac4ejv/8nLgq85gGjLNgQOLmNV/hvVWSPaKRCSVQ/yfzOuoUIclSEwL
fdknZSj7cWYSnD3TCRIa3VbUI7HXvJFk3LZZrz5ctZoe2oyE4kZorF/932353RYd6jOCbFMDeW91
H9Wu1PT9NCtoCtfD7ApLBFOMEL81N/y5N4Qms363ttn/azeYHCmkt3Wt0ws9Fnxa3BeapjZLpdna
7e2MwdjKvgakzA8Uv46n5Do+ffZ/cT45y4f3nrqMS3mA0usvR9C+78PIiEDyIdejXE3BjKTGPkC9
JMH2/FixmF3fXDv1ECTIeJ1ku1P/8F7jlem+b2vJHySbnqTteDWYjCuHc20oTI0/V3OZwUPBFC8V
XOl/a5ajSmwzpGPMRFrwsL/Wr/MOFhh8nI03XtdHnOvZcu4PZ3EaC+Ihud31uRaZ7advyARLu/VT
7aBe9lUtA5PwfhgZmjkBFuI138Y3TlyUTSELWl6oewPydaVvWug2bmTwsq1ywNjWA3tVjvXuePmI
pIQDt0b6VQMXh1jS543RKzi5GfXP7h5Dzd43JeBpxcTCyWfnR2hVXwYUUgXwJlwOolCUlCZQnzQP
CunGTO+8d20TIdlc/AxMTSXzjCk268uYtkbB7uMf1JBF3gy8GHJIKSMViYS41ZS2sAtGb/iVUK9B
VWc2z3IkjxAUYsZ0JSQh0NqtLGXGdy+szHzQIV7KDzZ4gsVcOEOL4jXa8jW3xV2HaZ2WwKdMWhtu
7OMXgcM14J6ZDVYVIKO5ns4X16C30x3mAuSvkRl76y/KbpFbJ+riytc6YeMdA+0H5zq3Pmn1518v
UI2dgXG97ywVH501cw7cTlPJ5x+50qBjaIPKKyYjvCh3TVU6XVDtH5MLbm33rxzjMzGMYs/4xECW
BgAk72CTfRqvG2d23GDuR3KF5hEjPuCUP8tKOKxov3JemAxLtxkNK9L06g1tLvkhA9tzoIw5Xvhp
Uv3q++PjviZdraCFUjxbHKfcmAWBNfKOg9NpN/myIthO6GKZy3lc/ulnOfdB8zAC8w1SXF8zConY
IblkqBvwNu0xca/5XfkmFHleSy//PiYUZ8L26ariox+Ue6alAPXrRRlJgCKjJfiBeNqplQy2PqLr
IkweAy4/ecYE6uxE46Yki1rCJADhK7gm8XS91MUA97+RswQvo/1Wns+y7Pcx+o3gJK1CS7CX21/i
D8U8Agit1jjIdWxCVWphICXOJw2MsNlmkcaEWB5u7mu7QKKj066rdMLhF9es5ud0CXaxy+0zXgAb
WOIj6GCy/iOU5VhJxf4zg4T5kbZEMJSYc5yPRey9ax09O3kdN2kwtd3eVzGEms8A6lzv+c2qEVR+
upuXtqiCZ21DxfXpuNERpnY46OuoaBC2KjPPI4pibmhMjbSbowcnmSP21SCDHHV4S5xSbNs+asl3
u8LBY0xDlUq90IVtHEdZSI15Yn5zN3UR+wZJ2GuDPzHwWD9c3QesRcE95nOJ5pbfd40CljwX9Pyx
YX/e86+ntRtA8AE+gQ1Xpj2o9s4NacStP0eCCWPoTUd2nEKj2jpBul89q4/Z4MZW4faH2+yFE4Ev
S6DTBDQKUMgmywjSXgyrNUudc0OSuEi3uHVFSAMWFJCfbHYg3Tca1hwLbJ1PvuZG+pj+8Rq9nxE2
Yoe3tufrhTL8U17klRe23pSylkCIKazCDU3Dxnj0RMqhEe229HprRFIfT1M9QZKD/Pz9syrjZ3yb
8sE8Lu+dvGfZ/ANe/pxut+BLs3xFpgrcUpmP+Aa2gQURZ1wv2V+iJ2XlhFJG5hgEqrOrUusa3V6n
7irC5OuLeXoQhcoRZ/m8UFd1wpHT1RIh7KWFiXVFqfoY3fV2ynBqNpTXPkygeYWR00XvvY7KjjWF
JDWSxXf7cEyTWu2nduEwe5iptImG7gdhFLYCtqw9/Pnh/rSqMMQFDdXA8hDB91cKESrxUUKjmeFA
cGQocRwFdMmCnS8yKJKCLisHoOdT1bPOl++jjGO0PScAEw3PjsdlO5yAlRUc75YPUSIzjBjEwR+D
xaWbP1yypEJwirtF2PYnJb1jXu4n88JH32aC7f6NRMHfLYvnAntvr0QtlJEnEl9y+qmKsWQzFFbV
FzP+Atx9ck2IuWimc3vQ6KiMOs1WiEO4dyiPr+KefNDS3kuFMz2fU0BFRDqB6LqzWVo7HZ6luwnu
kPCKQNi4ThUUi5Z8j7iI5U+57Lby5xQFbZeqlw5GDoi5ORGZ9wr2k8vGCxXdyZmHbIuMQpNpNmbU
CvmRnIOEXoQ1ILTdvxBKxaGnMKd/cqpxl1a5uB+bzZJ+d9ZpNUb613fuwCQyipnm5WKH2MTYWepg
ICQZe3Ub8h5y75jZMp2NxoaY71IW8xfPwtzloIQrW8spK8HQR3uLE0VZz2EQPoekD9NEfjA3xHqe
wrArBvaeobnc+/FLG/cpY05fKMn6APwdNraPQFUTccA6zTmojLWAhYDsPXBb/WujyTFOjvgTCw0R
SAAAarL/ZsKcdFfoP3H28i4y//KAM3p+aYTB6WPP4ZCB9DeOFbpTyITiKMkKyMAPNu6jfcgrySef
Y0O8yO8OodPOND8TWfqE1WiPEekQLu8Fc4FuNb+U1jQqxdA+X+sytPM95fKrEwfG4gZZf6nsg1lq
+Am9rNXtwxgDFh9yxusLCjqfvhCIR0cDFKk8lDngh8efmwNoziqaPfmmb9X2NczFZQBRT3X+tVkF
bUlgDQpyYd7J+xx1iWPS6VWuwING4JLhex6LSKmhUr0TF7ZhOh2dULFS0snovelALFWMZ6YX1wYW
0a2RYXl6+XBRyPUgKgtYOZifWtvjccU2jrkpeNw+Ubl6xRbqTSH8vnNkWrRxoPu6hstXOLD69qxv
3vWNLH5phuOAhroPAHqbpm0UZlr91PXQyUbWnu8J43dT5yxjw/aPbd+bUcf3yF4KBso1LIIN78IO
ysZCj+Q/zfKJEnF+fOnQ3AlMiYU+ADKo18zbFQd2hTcFoUux+uVo9lioM88XXVV6y+5XXUDj2lYi
1hto96A1zy31sA28LVGhNK7KbuUnO5YhTCiaxa2MdHSCd2zq0F1deeQRwti7inwZDRWDklYNYj1P
F+1Rzx63jYxnncSiKt+FwnrkemKvPgOAug1Pb/9LHkMHFqDEl4OjMBlM4WdhWJHYnfBNMKD8CDkE
j/QnAv+tCgigZoQdkbNMboV7NhvQohqpbTd35mr4VW9oqYuka+kZp/yZfkjl4imdWZh11s75DtgY
xsCZiN3yo1SWAhnqAZpbWLpTFXaEDbQpaLc2DsOvNPqwpRR2zfKmQnhoO2RiqBgY49kjCDWCi7h3
KP1mXSsKnZfLF8lO2KRxB1/rOZwsDsavBL+NZjIMGUBFwvD50OXK1uloxq99Gcgk/r7MBgozNQ2Q
UlgbhhzD3OMnNo/pdN1HZRVDDnVOKm68HStDTBZ1SzrIMyA8eFO5AilM957n9Uz1ELSGXjKNRFQl
Di9XQx6/pD6FqpuUtZDGav8S4+l+EVuS3PzXak9tPQKrm3Ds0KJbYXEeQU1cassHHKetp1npWoTW
Rlf+weOu3T2psoIx44ZlUd8slH/j+ahNZEp17pUtrLoNdh/FTsWEpG9T0EcjyQJgVWWYDZHjPFNs
r7V0kgVNkPTi5H84JWYgd19JkryF/PqJgwmYqVyBoSOhZlh4O1qFYsnxPfALzQSTzV3zouz8JpVe
Sv4f5u2DjdUwlTxL3P0LF56etiQbIHgLw4A0KXdsFbyRENxoOy6aq+Uli2eMNM1TCiE3nJDag4Qb
m1I+naXp0u2cXdKAvjbvUz8QvZBVmyHmcyszFq7IGf5enKD37FcJngFw4Qu//yHl6K8iRSoX1yZb
WsQrUSn6uQK28xdZgY3z69s1XeKWHAVjepcq+WwHnE9EoxRclQxDpEFsqAtVWS9aycktNjQRAkZb
miA8Adh13j8dQmeN7zRgb92Gi2ap7HNFOr1b6GVpoiyk+jb6GT9ghiU+m3nYOOS6QvEyU7rpMC33
ke/I33QiBgesq2T2yxXIdASJSnpwtKyv7j/rxQggH/aQiKsR2DgCF1hrKi3TWjVpEZTlndOBesq0
QmNCJfMB6tk6gr9mKCHH9RHCrRHKKMmTbCLj/+cRI4ahY8VU5XjWeLMIAvjA4ufRzOXgLGBBqdm8
r7P9FZ6jrXObZVTN28oV9gzTSzmi8hHzpo1NHz+PyECK2939K5G/yXNtgkfBszxCA3J1zHtki+8+
HC0GQmnhshxF1+FjntG6eIikR1tOmVkdot4voRXLQ3qpsIDyeo9lRoYhU29fkrKMNIyuyEkEMCX8
POcvOszgVqA6ECi1D3OLA3WZSnpT798Jtoi5Xpj/G7HjKhAvyzWH6YuZtaGUfwoUxpj3QCSqsQxz
9T5F8x4TbHWk5LIGV7dK9sY1hpDsbPvYLpgWh6gpog9+Z0OTSoxaaZ6w498Dg6aL7yauQ9p3ijRO
JNAHPzkZaNi04OKza6WaMiJFl05WQJVtED4pM6zImh1x4jcPaz62MktAdMafR4VZlE1i2c8OJ/87
T1YyLp50C7y/pJPzrmo6vJxxvqimc3mQYFcw4bScqoSjPJWZRxzoyjSprzQ+HpS6XE+ETYCER5ux
1dKrH8GWFexYhIMW+jvQWBp7Eim1g329dMi6SomciMDld0ABSGYJ9Hv8DoHturf1G2WIhnXTapTO
J0843p0zUeEEqcTT3cufu+0JFg+xaRY11Tbqbr33jOec6kFMTPXkcBg9XlgmCc4Fd2TcTSsX3yjf
nu/Q51EJ2zud5tA9vkUUgGk1SmrXpykPXV9rRlyjV3WOR+Sf6OzE2P03kySskM+EecCryJEuispP
AaFdwHWOj4bl4YwHIj+Jpaswpo24/cwcZTDvhCuKkzMdUn0/ypxwamRSHi+hU4RX4VDD79mduzMt
62vfWTDkn2nuz9wXQNpb9eBZXciMKJEH7l0H3xbohmSjGC/mICtte3LwBje7Qxc0sa2uMHz9Jt1p
qfW1qUiUnWfuU98lys0qekUUMJsV0xxX6k1tFbm4XYJOUo4QYzFMtzUuAQ8yovve45uEMgs1PKHJ
30guLtuUN0vuTWLKEVXX6okCF81I3sIqSd40OLgaAmSk8XJnIDRdRWZUeYVOcLZPqg6j6kTZbkkR
T/nLcPpDFtiYnSDtfLaIQIbnO+jqEF3ICesUog2/ZXd1z1/OIVKMfHL4Y1Wb4dRDLbpoCDmJc0Jn
wNtxQqsr8wgBnB1xQdDpbMQBsRDRzxeYqZoTc3iW99swdfSndGxnIuTotjsk06CZlZK5n2J6Hsur
Jh5D3xziugyRO+Vv3zLgfNF3rj8cBtACM31in/HvnIT2K5dVPoS6OCU5Hh439UATau84ziDDvauc
ejLn53Z73sAPyecoA56khcDxHL+ywnCSh08je8q0prbE6amsHCDzkUyIP+ml95tvbSmCi5tdqvSs
3/ltLUVOW+BHS+OW2Z+LFolAqihKiXqt27vNjCS5olSqblTBVlVTIpflXDLVK5sWSl5/ePZymg8M
wKdzOII9A3TOzuRPW7w5syWiWmLt0x86+5mer8hu657Xd04JRjexaMBxK4CSBJmW+qlJn4IJdkNt
MhpuCc++YTWkfyxR/cKQe1B8ZuEFstVTDn/3QHaUa75GxDukdZBl4jVuqEXe2fSO60JcLnnON60x
DWuT4zjpiTwIDZGvm3GCiFlfLtUcsl/5xtINqYREaKcJ1tzOG9Y+DD9s2GsSFLYUqdKm7AlhVYyv
ABpzQJ+DFkns5ZzLxS+/ju7jAk47VIRQaDbaPr7qGLpRfwInl3LnY1e7B5xheTTv2rHe8PvN9RWD
sl+Rp3BdtSIisTg5oraoaXXRQx2XP09OmDHaQLTrRXvJ6CcsVZVp2D9UMJ7dNyRKyZEEPsz0K3/B
BHIrykbajbnlC9U/jLGakucF8bYhJS5Dpn6BgL+eTgRqKmeKsHDwvs4yzV1bbuVvK3UpEJ3y1T0C
b9m0KrEB8AFK6nRi+5E6JkrmODP5N/KMThn1jvCHqsUnS+r1aLqB1j/gSmow/RnN7IdeJJ4bjXub
sQ8Zyq6/rVM+QsewETmMnjOPjdGyVJq2Tc0miLVT8Iye1mrGrRXKARTOLmoJL6rqBX79HYOrRc4n
oOEi4ts3mT7bCn3hfRq0obmmPVCpPEk0dlakSvBc42UhI6b//h9FKnrBZiDKrWapS6gx0ZzkL69N
yCO69CWywtP8GNoVT5XlS2bVnZ5nzBI8fhOr9mgA7x/Nm2/0zk9N07hJ9+OGbAq510WpQCDIcpaH
YFf42v7m5lwh0AP/20qDrAWyCPexN2opqM/bIBHqA1z/YSpvOL1BgZ/vcqRqe+xV0rO+fdfF4G4Z
WEeEnYybLkOYAvV4HtbV/zqyXyk10k9da21fSucBP2+Wk7UwUGnwKMlzL95T5ho9FGiEHIvlcXUc
uQixpFTP0RWVwjgR7Kr1BYMTR6S/AQMASa+lQr76EMNP/eYl+jluFVa2R1+eE6MQBZRzCFCi5ZPG
JKqVfoun8vKLP4z6EpvhQjNgJ8F3iJ9vYmd+5CXDKwSob2hJfO0SrZ4BjVpPDinqotvyyEFduO4p
YFDcEH6ynQXU6jTnvjwiZRDbH3pmbJTL61mZOAlDa5DFtbcw0AKpaG0syJeIQ12j9XzvVIRVu6T6
jTlwWPqeUKbzzc7Vj9QuBRuhqI1sjRZLpe9SI5pO89VTFdFyJsMGpBq85KrWjdOOeUTzE9Enoq9t
YAnT0HdOlO56nJLM2TxAo67pAnnAHBopsg5xHGMJsTRptoNT/P6dlTKI4sWE0Fo3IIReoR9tR570
oAkZ5YwiLBu1lr2RBerB6vaNQaUAuCsxnl56R5sHXnDVOhbznrO+VB+urGx2eD3669S1VZo+25ez
Dif2BaSM2z7TENnr4Jbi/+kv5aS79ak7xQoe1FHCnerqUtqH1nPv8D+/Gr5nGBAr0LTDV9rIAY4K
HpIifp1BxNS5thWRN3FmyH6PlL7W9z6W8MFTLAvFTpwrXzjT3qZLWgX0Cjrr4oLx2Kp0OvWwXrGt
wDETTNC4jy+Hdvl4R+Wks/vBQgMtaIws9WPfuCYvIMrFhEVTu/dKCEtAX4A243RD5poB1GNMvfAu
Yc1dqz0azf0I2tEOmIdU7o+FrDDDyQJw+o2Ofw/q5BNRC7EVd3xHGxjyHYjb49PmQUCZGIJ3wWxV
d3I51Uai2/501KU6RuLppQbq2p/PCh9Ds5FaslsPZxZ4RsvJtajdHrqQ53JyCyEo0t7/tgdInRU9
R5OySVHc3WCo12hKVmlxClHdwZIpMSKNnFFwNNWvMC5J7fwbES/Vy836x8ibC+0+RA7rtMbF6f7K
GQyCVYiD2aU0IuBPIgqatuzNBtiZVGLaPE0Pr6tvFLG497TNxH4A0TzUn2tgJxEbVpbusJuw7rdm
N/FS8ttgcL363AV3PYwqTWXvqLdqFHx75XXU37A2LuQIi+Ki+F6oGonUdfQgu8N68Nk9Twl6HsYi
DmICwgiRwtWIfAPFVZzlagF8avtAupc8fiGbXFAZVSNPj2eca+c/cr3SqVVLv4DhF64Q7aSbLP5x
8GG+vNCTOSByg7tCYrxCZZ6bqEZ3C8BEpFseSFwbeiluxf+8yHFF8hS748Y8iLM/mKa7O2RIokrP
7yYKbiSNACIvhjJD4sKQQ1SjL85xzpMm/U1bRSUPzWrA/3hm5tIPhHCXzmoGq5kJBCY8DvXx00x4
HMpWvuBjHIg93YpT0P+2SLpuOIbk3UZnfQ68Euf9DVmWNnKS4o3SlX/YutUtM3RuTD/jf4CGT/d2
BczJImqv7AaC5gqRb83V0dVxXy0UYS4LBLEIEgPmYfQTtZ5k0Kldoh5WZiWPV2lEmCMXjAmJuFPN
tkX/7gZKlRX8YTgPaXqV9wzoILC6rBqqo8geafD4ThLSiCwoM1YfylyEd6H8BDz4ejUZWVMnfeVB
MKxCG1/gHM/bgB7wJJk1jLP7OgZ0mps63wqneuxXLaAYZb7rwt3HxviP4uZA2+4xuAAkAR3HsUIT
3kzW0/X1tAu87ebIMlgQiHi5PHF2YHWKa/RbySX9jgFfEOHPf7Rm6LKv70BIJblrKyWpbXxuQ8ck
TryUqXYSqVvqux1N97TLllp6DNp005mNkHouRfX0YjbLXmw8EP9jGJ+6X4cl7oX9+ZGW24ZrCYv5
vMolz+Bq9PYtaHhgoYT4hASzJYfdbu2ktPfQAowJWeT9uGOnvvFFE+UZwFVkBa48xq2D5fzTEtqK
bocIPsvRf7W/i0Zhn0nSHg7AUEV3f/uupNHpLUjs1Oi977jlN85X/iTAR4guw/78DW0tnGpaagif
Sg/3B7NHFEKPDOxea2jv0QvSx6h/Ve6FxwaUz1KlFh7AZmLWRjacHaozlLLB6mesgBJgb36u/eXI
+EL5p1nvwQCbxOiDaQuIc0S98ydoyd2NftGgdgprV7SqFb4DnTdnhg7v/eK9HQOCMgSpTbuWyr6b
QUt+3xhLmmMfaZlKyfOZwm9G3IzqJ+B573+3zETNu9CTWCazsufX+0ctav+73lE0Sos114lGD255
4oEwYA2FZ2Z69sP/50cFFziKPqP1ljScjVttr2vfYBt2yqq7pOOkxF4pYYRxPezvJ2M1Jp4rN0ny
47PC9D6T8OhVWGpAm0nicaeCO96x+1H8p34805/8ycaUJs5a8kMxFVitDxlgjHqxXB2Gb8/4DAyb
ezWGIor4ygJjMOL20r0Y//7V8Shr2XL4/8aSJuEpcg7Ee5wasuCjfRk3IpNlQV4wdf4D4EIFKPtd
JYlZw7cJ8FQFKiH2+mNd/np8bh5ve7Vv9EkCtomUv05kvtXbbPKKyZi/uxPS7OQhlEvyXvAamcqf
ym05rxI47m2Bbo543/ZJapgiEYbSQ6b+XzQblqkx2oU2K2cSjUcPPfAY98cCRortcYXDyKVXgghi
L0Yw2AE0kkQug7uTAg+w3+wxSqZzHgWfp6RJ6TOhs4tdb2HOngFrb0wu7EBJLzDoUk2mF4ii8KtE
DKi//c1YG2SEQlwGd7NROHGa68EdXv344lfx+egDnbO4K7bF+TnzqWT2Feom9YaF4Uc06zxxcP58
fgj5qxs5Q3HgQcRzkDF0sSxU6O3dM97EQv3JkxYGcDb0hR1Jm8FjClckJ3Dq0zi+sKN0VBWOey3H
ddBt7Ya6mG9fOagA+ceMopTSbnoBicQYANh0OuD5QT4SmKp/5Hj44l5aDcZJAbPPAZU64mRr8twf
l84KoT9x0+zMexSiaXMoLBNfc6YZHEL9Fxucahf7a4IuZ+3no05NnZw3l2EGLYUD6lZCWGMBrlNp
G+xYlwKhnYhE8Uhr0XutuHw3VLuYZ4heh+/9L+SaNU0uq90I+kDcKqzKjv7CdLmcF0BhD86qAkM4
a48VeMxALtYQayARRq/Ut1A7lRpYKOQeIfO846305/d5k/l6Q65ibPOjmm9G3FBJGOTaulwNOMh5
UCBt4pQd2O78wn/xbEVKR8qhDV/oCb/V8I8mjye8WldvdOTJ+QTSKi/LjqLBSLk6VwbAD68q8gkF
+yCjZHdcqXeampIMaVJwhbzQrEHAAvholuk+psKRsstUBo32ByVTcfEyyxU9SpzxsJjIbs4wt4df
Mo6NxEqNUkw3+Q1HXwWH/XYSKBWtx//m5B0pHEisazUjT4KR1pG6tvagVmutsbVqv9X9vB1BX7Ad
kbH6N/KgxxnfnTN7NWGEWqubPULn0c7gikKpn8d1Ct2mHfnqR0lLGUyiU+0+ER1s7jcoSdYvbKfR
OFTqNMcpl68WqL6dcNCrnGKpimBUR3OTYAcSHO9voDtuDHHMbRs67ksUCG3i5ncDgd/BZl4jRE8e
SoLiCc0rmm7TYo6gCL10kNxVdAJOAcoBwvL/yCdL1Q4jZR+lSyb44wT+PoxSBjG4qNN7gUtD1/Eh
QRPm39kkq1rXStG8YFANqf4vZWqeiMNPLXCXs8CiYXu6iqsRQrNyPWGTPWc3g1VIQeo9kCE0OYwR
QHYBonP5IITtdjztDW0VznyVxlwG9lvTHTuIjwE8bVOmCr/z0+Lhm5sYtJv7ZWLULyxogf39bLL/
YexNNpcV4OQ7c6tQxwH5ftMMr1Y9E90N7JF67zoRRbph+X/5F+6xg8UBGA1mDjb96D5fQ60IDEPV
8BwhlLJnIF1hnhuaBELQ1e/BP5ClUTIxKWYPZnYbv375wdrMnF9ZR0o3kJA7egMZ/Mp4nQBUFdLi
d/uxuKCwKeeseXqOFdZFQc3qQIv0VASxRr3U8A9vNnJSG76PTy1WVjtu+x7OPQmBxmVZBpgOaj54
4gdwD8osYGqatoGn/RpQWSbhfpS8yaLQjKNHX4Uw+Kw4Z0dDcIXkWkvTWBbTq5O/kzPatd4XsoE9
dWp21PAj3wAHLH8ArqVXmMUa4/wrctHVG12GMfAI/be6DyJOrajTrSfwoqGQ+xbr+z4vhky8GaoP
heVLIawaRyEFyBljc55k2F9XZSSOR4APw5BQC7DbreNadUJucT1PBxO7l0pIzi4ORrF7TufX1uSd
ihogb93VV2dsV14tCaOXJVR5U31yBA24ZsVQVZ8gPUc+U2vfZWQLyMN0lF47bTJInJ1QGtyNgfbm
Jz8r1YygwdGAOjHo/Hxj6KF1Jz12herAHJ+C7s/ZGNn6AojY1tpHdQ+WueZ0LMnYI8bRU2WgnZiv
L/odK6NiHas1LiiY72E0VfgfTjtyGNiegdqRk5ae6ky42ZRFDQrhX4gOzVqjoBqPv0Ivyc+rFHeN
gd6hrPd9hb2Io1XyCyEDPCumB6pU0/F6/cOwPH95MVxGaModlXclh4o8cl4JJtL+yYnxjTP7EIiP
r1OimFxyiS89Bziefn1h7r7wLL0lh5Seb/UphYdDKw7Y99lczHRJrxufzKnUb2JHky0xRgyXsGO3
M929EnyaM8RGyZC6yRV7HquFTgzu6qspmMkxlishWkW1dpLP4MgroPVPvZDDWp6uwAU7teoOJcGf
oEcqjgt5mhobXlR1hyKf2grcDM+VEparf7OSLy3ZmTAiGP4s/qSllHylHS8uivo5TA9VmOLsl1m6
rCONY6dH/Ky4Tv9aOXGf8mQJHXTU+RVoopfr7Qq4n4L5R0P5ap0aTHMYVGfwSVc6QaDixci2txMm
HgPyUJU+IDeqkas7F8pdwtIN1k+iRMynBhOuLot1kAxaEj2/zUgb/o/+al5L8IAU6D+IlAZ9qLmD
QNI3wqJYmj5MOge7ZEvCscYL1tCxFwa1Pt9gTi9Rg6cd4wrJUfK0WEpjRaqgsagDIKRQ2Qpz3hts
JMeoJ5oPqUyPUD7MYvybPTv/wHPxgn4jcmI1H34ohya5o27/fs+V/hdrQ6Fm4lf5syJw12v/Qvve
mTFFLkfXST48+Ewis3x9pKPHMrFYd7952337dK7YNNB9ZYXPxUJjuFcAqL5C60YDJ/zrLU7vBKWa
S6rPqiKRdqLDME/YAZdj6QuoiA4E0L2bgPv+oWtc6yYBa4xnycdoc83iVm+yjdUIxcEp2JmcG7Xr
BgbbfzAtknyIKwvD1ywPJn7jisfuVWab5nEe86Ft1LImuGPWNBFefBpKzBogO8b9DZELMbxqwU0r
JwP/WI3a11KadKS2wq5A0Rb52CcY+fc44lYELHAyTjvmAlKjlyPGqKxFhRqLj8u1glimXBtQQAnN
Fei2zQ9h/ifMD82ZJXB3ai20yd+1x4TtGKlBk/y6eOH3kJ63RGmNo0ZKb87QxPV8yNdYf1yCST5e
+Dz+9RqBD9o7KBqxa+cq8JkO53TAVCQoxR/U3lkkglO3RjdnLqeGnVXQutvadb4/SJ3z8IUgALiL
ZeXqy4QY1Efcm5HgBzPrXeGbb7fP9fp1liHJAGyqUhNRhxVkOym8/Yz8DSFeKdIj+lxrl2LHf0X+
f62a2MAu6hpW8fb0n5U3SkjKqnen0tQG+KotJYxwhG57H7Ai6u6bv3Fm6sIsUbvA5ik/8P1JthFJ
zhoPGHq4KcXJvJO9hkLF8MN2IBl1vKCCrNWrDSz83cm8YLOAWIe0vluqxXHwvzj6Rb496qzYnHC9
o9TFKrF07bRhNaHe3c9cPSNjKCYAe2bXDl0DyCsAeTHmaLR/E+mlogK20+S7TVGs77afSF4yAaep
JaQgwJJDGDtWCUhUwALthvU6M5Yc280OiP/akZ59GSbPWy6RYjWk98HmNp12mc2fNPZVsS1v2W6e
9OC/8biNXYrfgbsMqzQ5KKgPkhIfIsCQXgD3em0it8FNlk4R1W6q0+3YTPVxperitMLff7XyCnN/
+dyPPe+4HaFdj7y6Xn4B6JiVksypc7C9c3gbx0G2KLOm6W80XGkEzCP9RCJRrCBYQvlRLoUVYEys
fBoc8uWN52iXg0+x9Zu0GGe+Y/Tpm+DUEybL2Vxd4Z0zy0MUtrKeOWSE1dzHVNTlavINEepPix35
4q1Rr1vIy4PDS6N9tdXtW4oL4C8+SX0WpzF4KMhh7+YEy5vKKsBvPRpSlCbzlOdVZH53IanZGJt2
cw61V5D1dfT09oN3vRYEDR0pP/yeDjJvDzAGzeCCwKENK3AX3r22+IXPoy2Hat7MQ/Ny3UYQ/dVE
VsNmyyOloxIRz2vArgAnDmY0JZsclQ6OhidWTGFwpHvEdPx//a7RE828Hm1xFAaH6Jq5AdgXqjkT
NI7JqvFIrG2448rg9y1XohTHTegqECkExBy51vO8Dnr+wctZdN7oFnvTqcu06dTe1MchGaXKpJVK
RVQvw69sQP0b3drtwLJmM3ZRTJvg+Hw4D2KRD9+dGIdzvGPXmCKnKQOoQUwtceamIsC9o/Qh7LJB
CO0QwzOGGMT2vy81owtAonrZWva4jyCfq0LO7gJmV4bJvVhFrALoypIK88IeUc9xfXKXAy7V+oob
CvmDRU3dCQWsNJukOq7ofHgePHjaCJ1/b0cHop8naLGa9rgR8+A3cfUC5my/6GpzpIIAH37vNLPw
f3QJJa3ZLKOrKe/SmOIlLNuiZHGNWf6f5+rkI6oIW2eD+gYgmcoKfZRdBaWnxa1DC9sBOQkDW94a
KrjHo+aalcGvDMZ7yCrMQaHQWREL4xpdn1jShuKuu0PvEtl5vG5qBYX5T86jcFetoxyZyRY1ZDHI
XszUlEJDYpSJ5HAHswttERYJ7nGs6qzGH2jUHnAVj1ZZLK4SCtxL2fJl2RLzWX9KuhV4DQHXCgmS
jMdbHemz+Pi8LDfiEdr8J+o3GctIJJ3l8vL3aDiYxHfLAB94zGb7D3Zr3R9JQ4OctWzHwmFYVtmJ
uAbu6otK+VVSj8JeE+aRxEcZ11lC6lCD/1nCH48wzTd+EHoEoGFxZMApHpENrVC9NqY4IImYrsxf
APHagqi2xecdv/N91UdeJc5Hq3Q/XX+VhrKESQ49n0NHSke1x/2SNILtEvf4s3/LQvoC8TGoxgQQ
VRcG8l0RJOXqrdetxiaid6pjdMKlqUPoOd9/T7e822oOF8Y2we/xfqcQm1eeo1PoXcXCDuu7wfdK
A/VERlTMx5NRm0zYK7ZNaQ2Fq3vwK2oTdxSAjhhOw+8bgiuQCC/WUcdzPy4motV1/k0zhC8jvoPf
1Uuk88GDT48I7vQuvL5vA92m1DI6O0cq9RaVWOQLxcHKfFdJ20tP8XRkU63bfEoPmksM4KRCgqYz
f0d8Zjl+HCSNJvOCdgkCrE3x22dRJv6EB4JsBhe/3nuM2G1fmcQfalmp+l2ln7a8lFCzZESF7uCO
OXEp+QM1W7MaVgzLl24Zs96thPvWk3FPq7GpwdWIrWLjbP3ivf27pD5EEf/eJgkRGtlOCL8GfPG1
jZjmzX/1TNc43duYJBM7LlqLDitIHj/2GfarH8vey5HGnRw16sjVqs6zBQuMXgri71SVDveB6dc9
pMPuGJXyqu+QpYIbJ0pqUAKKcaIa5qtxQzQeWN9cXbCvp0cKehrvlcJ1JpD9vI5LjaHO9IqQh+9d
mbWkiKOFtaPyBKUvmq6QnpTx4wUH40yJtfXyPCHXqAXjPbjsGMyPlBm/W4NuqlvR6dPfurhSTHe2
5T7gu0VhYCGoISzDnBzPvSEP56BRVLSQFKGdYRvd+fKC7eK1uecaHLzZeCMiB0dw0tPUOcwxFkEy
dl+uOTbIvOdKaiZQR3QmHuaUVi/8zJH5LYKEBEVWFnckxQy2mmdACC9IAmMVDrUnQcgrt3BTZILo
Pg/j2BkAl93D4w2XQKYRt3chKLFXXp5NjcniqXRqi13E2OimwcdhRzDdebZSg5pY40fAAS4SNDMT
n7PH7MCu3c7n9gaUWW5EduFvXrD8/LsHonlOr9oAm1zT1CfhUWg/aTS+K8I3eL/roOMSMw9z/dcI
kZDU0pyjNwFU45oFyV2G1HP/chJPmhzP+j6cGCoq7RU8me2zt08Mo4FPbC+D57Po8EXJWTsp2pFN
ZvPYuEEAlqLjL1PEyVBI20/vsVBmPkRgLLcAbZp/DCj4/luswHQhHW/WtmACVlr5EKXmq40TLzRL
0bqnWa515be6CRM2JgdevT49NpMSpLBy2kQ+Oe+KgytyO/+FwjGKz7sUrD28vl43g+HxiNPOckIu
WU4D4mmOtbZzupxVRCgQCzZGEhG4nw7c4ZfY26C6C+OSrGQqqAzWVxgjOb2UX4KydoX8+wc6m2Jw
9OSra3xUtNs3YZNWWR9pY0P6dz0/X6VllUSKiQTBxmvbpAmGPLpLQFwT8GUXpUSwlMJQswjekmkx
VK3euU4Zojda0NQNGml72dbmb5cvbheJdzVMqOeQnhSNvqJ720W8L7N7N1qJsbXrJqFKTKxVlY+o
AsCNs16pCFRwh3mE514RA5bgvHvkzWCt/xmT+0fwC6hGR0640DR84xUJjVC6eVqCRff8Z0gvTI4e
3Ijru140+eGCDqiqiX0kRuYxYbWlimOQd2zK3/265gGN6O6w9YOftenDK81i5ExjNSV+M1IpdR5M
yXqpV6e1b/NjJTOWjSVZuYwkODQJTbvqU3mmXuVjEZ5RE46Q4XN4AHk8yg+TZyN59F0RWAgfCSDX
3uZSQOLkSAokgHczgDIBLJBToUmvNqYpPmGZblxBClgs8uKJcfiH3/F+7WHf3nYyX07wNf9JC9Ed
5vzyFgJeJUyPTIFusK5XZyHPQuC1DeLKl6lMc4QRchuAa6MuwC/gYgcyALTZnzOKwtkxx9DSFvWs
OQW+hEpiV85v3tvG7YW5aQ5VwaEF0PzZxGbsBOJpwdX4zbmblIS8RPChnFc4EWFoRGR9fPt+vzBm
zrfnYjG/KrnjAXYq/ekOpJG3oJxkzdVb3Ip7cDEj9IfkzmWkgmUos3ZvqRc+bXZJw9nDXBJ8NeAL
d83neX0usyXFpRO4gJPunMx+NJJCzxtIR0fdNeu6LGOwrwFo9b6M6RSebZxbCr+tRCzZU2AbApc1
dccVMJ+Be8Y1BGN7ZLB0UHHE7MDlVZXqfcO5c/JPKnp+VkBXaCwPuzqtE1jfdsas2HrDdQOvw1+S
fAVpdyS3DjBhFwEVXK859kLIjBFSZTtZs6pr8oV6jkP/J1kg3FsFQ00tB9ZOGciuR3X2qIfFCzhn
QQCQqINJJzm0VWWDhoPhT3YBYwHFk8V8pl9gskAcXISyNRoqusz3UHiP8Uf0trbHoB/ddtmufR+I
qUHOJ1ifedVxNp2uRSecrfeDM0d16sW9V5q+0nyyDG05KddtL5QN2LJjELMfmo/tHhaIfHvOpidz
FZdDQ9dIgTSXUSdAV9O3hH1NmwWAEMa1tI+oiIHPAVsjC1PFY3FXVMba6gqlK74ULrlIXOLbWWlj
Q4ZDXByTnKWNwoU+rQvCkJ8hpD9QfqpockMP65Jz3e8zQXEPxL7aHyfqtN8Ht3j8YrH+UM2hsYro
jCyA+UJnSQHcsL4QSe6CuH9dChii3f4kP8ZGDtPQtDcGYNMW71vRGKtvbKK0UECxg+B6fr6GtH6c
n37VV8P890x8giVje3UpA28wq7eZ04Nmrhcb899CXJnw5aezWhjm8utuUtVnctY3HSgT/rNWd4Pl
rX6YgKth3krXSLUCc99vS6o6R8XbxIQpfFDJGeLLoHczEXsx1Y+9pbLwBCbmHvKhWnlyEjlS+fYa
lhxSJkzMZzDkOXi0FI6fX1XdIBkZiXS4I4aYwlyfIg7+uaIQkiv98L9GbZx0so03tg4zNt3LcFv6
v+xYrPf16XFWLE0M/zYUAUkYz09Gun90chRJ5D7juzkSWLk+3IV2PZur7TaWDrM7wZsehF2O16/F
AjqskAG3f3SA4CTdBkphPl8zwNlWP25mcQk8l8jqljz4HXbss59kA2WLC6MH2i+vQOFqXSgIH8wl
8H6erxpmXw74+OOUVZTjEQntIsMRamTxxgQRkFNQ1uLYYwut7FHzZO9Ym0xyGxtJlHNU3dcspUeN
udExTPkUFa3+5EaopjlJKh2eXyz0mWEv19i+ose9XEK1li5/1wEtPjfuS0CcMn8I3Zfwr2eI9XsH
d1JICdr7PQfJDf7TzZL4afQ0x1t6WiPyFv6gxKRf5TXEqa6jqWVz+0+3R/R1s/y2SGuZcRVh3N6r
2zRJ0Puze8GdeDOfKNDbc3NzXVMR1oLvsZZyk9YTzunLUOil7n0RZVGw1vnyZ28ntRe2vxsvew5w
97nwrioxsQ2O6Ec7FiWUd7qzGeoBC8oMkhh3u8CCJHshQkGE1KCMav04dU2bBXgZmmLnGiE5DZ5A
fpxfE01akf3qu3wySkswU7UhjTH40+flHg/uW/YNa3eB1RMyc6rfHj7DoYT3Z+sN7Rh2YCMwE2Dp
4kH4RiWrGi9tK3cvnX1xo15wd1x7VmnzoNIWjhUSO93h2NBdYDRrRuu0SBMShfWSUpgXrZ/wwqE5
+95/ygxIKClbLk07pq+UMy/jdX9lPBD8pe72aOu22qpCu8kVzB7NMEQXlLnGPznzt0Oq1h8pgpq7
kEVaE9dHZ/e8Uwu9s48vjN07r8k+WPk0qHiDghZTVLloel53BTP3YXUIWuoWYDs5IgiCP2U9HmqB
U5IFNy2t5k4+gnuWFbTOFBjX3hwfyQo2B0ZYEjUR/Noejh7ZeD5ZnILvpmOLIb8MyWxziTOSUCNN
qKpHfZKnPDIkV2Br1LknDFpbnL1kXM7EL2lMCCw4RnUABXLpM7NpdimvBa/Gabl8M7WkBnzynLdZ
yb1M4YJiI7FSP1F7mKYjvLQ82QPa7RODm/NZv6t6Hm/IeCFKeA9n0ZelGDlW2Ch1bndBJLeLlHt7
RxZMDxJpBq0Z9ek7EUGDDj7VdM8vgBhVy9d2kbmu7XtENYbYoYmsnv6IlU0g5z/VuDPo3ChFSKA7
T+VifyN2Z9vKFqIvuVxrdy5A4bdbmDI2FezJPxpYhb0g9JUUgxETj4r3wQ90YDgWA/Y+Aoru1JZJ
9rqTi9c00WoeCiL7A+lGOoKY0OCNGocwxoMAHX+ohLzkbrBMcrd1q4gyWfmD/EnA44ek/RkgF+lK
JvfMzND5QQM4O/upuDq5vBdB8/ol6w3g6BuvWnLC41VOFyBLE96RgamVOyZ6/Dndoal7ZwbW7vAC
x9l+CrJS+kxNkEwhSE8da0Vuzn0Af1fs2ne1RNglwTho0N8sAJTmNhKZbgjP/jFaclNoVmGmtQtG
Ulte0//kGjZB2FwNimJYVTS8sFlG1Bp0WCfzaH2rk/hryhCVAP54sHXnQqYbgfAQGbj/hcdve5Vr
1BWwlwxXWNnVLcSTmRMmzm/Hgpyfzc2k3kbQwjtm4o5nQyKKD0TbG9eK4BWEgWVip6sxchzzLoYB
xP0yEvOjClpbMdo2YiFNQbjgtdScAvsa2LnrGyF1NREqmecgbQ7uqnEvO8ExaXoIaKxOsNFnH5UB
GwdocVCZFlx+GunJ+iakU2RQzqHnNb55d6tHVkvVtiLZo/WSfC7qqvpHsr+K9eF2v7U85yz3vjDJ
EpkdZxpqK/xT0LwWkpvkFSGd1RYbXvxmEzDgp+T4kb0roXNgPfaNldX9fotg7fmMEDgSuxukZgm1
nLW2LaF3eb1nLu3Tryd82IsyVcHJ8BIwrr+psEU8vCzsYQZsLUi74Brf9Z4+mdSRlksHWnxtXRMj
ZX3yxAKqCyCEliFk1is1V7ZtrTHl5PyBeZz8Rz/YgOGwct6gDF5vWvPkdf/q9KJullI6PX59Yywn
dW2ZCDDFac/cFK+ZEUpeyO+VwHKHFQcwes3D/Yac4Hj+BYO9BNpv0c8L4rmjp0aqfm2hurXYYWXn
iJmTPh1SpkTEH90jVAE2bRCTyZL5943mNn5P6NCcBo1dbGJm1D72FsASQvDhvoF/itLVsWYCRbvB
b31hWKKHdVa2B5bWNggWRbNwPhQXsOVaw5GLdlwHMWCs+Ql6t/P14yUZu0nCtRi5D6s6qjs4NXVU
gsQIho1lNf92VuHrP6dNKZe/XvudG6sQCu1mK2J3OXYuou9UWMpnUKJP33DhBNqGGFKR/ck7ai0i
MKSVoFL7OWKg+3WDt1K2SFejhISO5qc3w5HfX+i1npLMK93cKFQUmHl3/DARNNdbXvuju239K3z2
Bizxb4rjEkzdt8KGFNurnNl2TzoM4GiRCtVeDsx0oRDupzo66hxwJ3Mz+6cictt7a3YiH9vO9kDX
EocFiIaCmCpLxh17Gg5gHaYR1xQGpGguRaFMM3GiT+xYZlzcpXkwA1i0Bn6q5UZqCshw11khVh6U
xex1dPuVm+OySeVJocNySMPWkFk/EKfvOB0z+8pgKCSLGqWzSnUAIkJ8d8MDLxSIHeN4wy6hyRJM
erFv5uf3jDAj1QbfDxFMtx/kFAmDrEnpyoVBeVueitly77F9lRcmxeA2z4Opqkf89GAcoPf4fBQS
USVrNmJrtwScbOX7mOh9C/UPuf7Buw/WLcGDiNyXhQquwzdKJd51p6+ljepvTF56c/0IUm9vB9CK
u/4IkcRhzmX1HTvCZtRSJggUmK7GpsfmR9BBHoiodqM5kcTk8OKvilopSIrkbsM2kWQ0TtDVkcXC
dqA0FGLUMORKpoZxMJt7CrCqecZ37PS+oAQz5WTHeSQG54ntvpYpB1xihCJi8KmNRsBfbgz9QTh5
3kmPBpGgPv7dmHWqRwo8MXmwzEA95C/LZWQMnUhbL1UTullTh+WU5NGIRaUXGP7TSLyZa5GzBxJr
8MSgoKYrCadD1K9hmJftaunb+uSP6upEgXiiTEEEYkspeoBnQlG9nR4OFhjlq+OT9IkSyjsC/Cjm
uTD7RkcJnQiTytMSYRjgvv9QJz14/S2CBVY4cXUziIVs81olmVimJVqU3yxLNMiWpuJzyANwUTgd
/oQ8AT1K4PE1i5JXZ51COatu9K1y0cejoNVUoxHtA4ymbbWDlX/xFJfE9oHuyizxlme57zmLYYCW
u089DjObgp7MlQ6hmj6igva9jA8KVa/WQHw0GKCGleqN8nKI5aLHtabeCZFe/VibYkuIl5auliP9
Z9Yadbhb9cF9SSpXZGnWMGeSmQOQ91B+Ybu/PsqhHu8naI3fq4xC9E312UnNYVrKvNUGdQVM/5vX
b7MO8v0ZdxCs1WhkgCCZeBACkyG48ZMUABXRq+AiRNgci4e7nr3X3vpiQ83jX7Gk2FM1u5LbJMPB
Z8Zld2158F1hDNEl3Qu4nzeeORpbIltoB7ikbCLGyTjDAT22Q1FuFZCgdzbzR8kztlafAVJvxLWN
QLVbnYaC3BvZibRmI/PZYpT2hqipJl6Yq9KRXUMY1aP3hWjC5khQW0XIttHV1lOvapZatOUYPKyH
/TVScZaK/urrvkiwb5h7LoMvcS3dkUA2nOthdG+l4d2PaGZmwbKPEs97ChUXUHfWglitGPylAE2/
6pCSHKE6Kcbef9YphB3rWt0S+jlY2nFeD8ezsgdGxlHljf988ddztQgVeiR0VXqlbEkpl+v1YSMV
PcbGtyBu1eXir0kcpfdVKQuzy9ZcKqwX153AtcE2MJIYleY76wMqqWF2Pp7HsAFWrsZaQGLS7A5h
KowqUAlCmeCgAPfKLar80+Bp5mvU63nBkkqspdndsdh8pWQrA65VmnYZfVKl3oC71hC77I5Y/gU5
jjIAgYxK3nEpRj/86NdpeK4zo9qTlu64mqv7NhLc7H5MvUx41B8Q7EGaILSsU2ABnf5d4ASX+GGO
rgogQXO6FPf88HB+2/MHqb4vPboxq2jZwrGu0EVBslgcm+5yA480Hwa79NAgtCToKmWh6Gpe70Uc
BpZuEqm44TPqH41Qb/IRIGscB0TfR8qR97Nx9KTETvAtId6thOvaIP99byP53LhKE83MK283Asoj
7bqcw28/M+GimqrhZQQJpt+Ykn3mEDjtXPCU2SBLMq4jj0YwHquJVuZHJXTlWCmiBfUJM9taPxwP
l9HvFt9bqWdOgGvklsuNiqeExE7t9vdnPSew/v2nLvorQroIsFNb9B05NuVX3mrTkkruZH1KPHH4
wjp9Msft93M4CLip0ulfJJ38pib2D5VdUDI0S2z/w6S0u9aDMkWk7lqCAWs3xzc0CnswCn9MjkBq
fPraxqka/pWQPyylGQ3qBOwh6U9BaFKN13r/oReZvP4P+HB/lEdGcBgsv+cR1pol13RaxitBsb/X
S9Uj4kAW2vSaAwXr9FVubSdlizZMGiMmsCdL6YwyoWRfVjSPHLKue2Vy7EYkgHYL1kABCIvjzK9u
UIYZvBP8QcHx7QeQ16GGAi30t3OpfVYd6a9Z56v6BmmaB6S3Hve5wiudvUAS4SjIncJu1r5jrHSO
zNMdDFkIaLqYJPJSygqOQHMIQfvY1C6clP58EQzcAn/BeP06bADo0ewuGqImOalnFHCfo1PNk72X
XLFmxrgf8LBv3zPl7XqAXL/5uUV8EeYE1S6gNBpqmU6Kd1MgYm3HYYVVQk6UbVKk2zkvlMMr61sD
yGzXi4OdEa1q7878DuOybgiVW3sDB6P4UJ1OttElkpq3uD+Dp7HN5IRZFtXJIejyAayfqc19vBQg
nJFgQJJo0p1tiukafhdU6Ouqf9pjZq+Z5uTT/n6H8XIZSh9P7rO2pZRFZ1gdU1rztZLiVJqhdJZY
qX2wIk4YEwHhGzhzQuhYzZ3+pIM/29jct8f6AvkgDyOben6PW3YHIqSaZVLB7at1uwX6EpDeH1Bo
P0IztHMh0M3fC3eth4R5YqVTl7+Nbcr2gco9nbqF8AZh4aRpw1pPaeTthpdCyaI6ywVMJnUnzb2J
jL2UkExQkJb8aF7aouISOozitWuTLSwD1YfR8lPCoFqSH/A1utUPhTkUhfJwYll+QUx9Atve3PMc
RLJELU/1CPovM87KkBoGHrMn3U+U1kXAv6Rip5XgUkF5fsQPembe9KSPeLF8EN0EqE1MlxBiInkc
i7ONIGy/2NDaDTZnNu7qRVxQAUnkbsXwAEkzWY3IUv7B66dOw0rb2Q8fZSysa46xWL38dWt5+w3l
laEwRSj9LGCIr494rDNFv4TnIuMv54FuJbZOJaMPVqStm7qkiWtEkUdhusIuvPgRTN8MO/0/idkc
WqV+IzHV/bOzW8MplyWg4iposht6fQfkTB+1Wu0EREHhXYDEKB9V6b483tma0c9gPwetkEo+n7Kw
dajfaslH3NNffUC+DJz7aUzwekIlow8GgXQbDB6xu6IvyPI6UXNPfM0WcFaVNHMi0ytQI34akDPa
netHm8BnPaxMkF++rsR5x04qXmqUtEBJjDFvh9jgLH4yPfMZphEkBWU2ySWFXfRv9yDQ7IKTDmGP
SGHBH4npOqsIX7tcvgyw3TEjQ8T2tlN0JaKuaMHbWCuatjWhAf5YA2fa5e/Ry2iE7jtjphmZW6f3
gTqwYn/Y8o821vAMUa1Omhxw0FJNZaB5Nsx95+ZwyceORRFZFvPtVmohzfEly5RjTb6Wq6nZhDeL
rstMwMJaGWmcUmaZV0Vv+i6Zq/GLTHsvSVrB5uBDVvAG4jXA6goEaebnHEpZT/FL4tE7EtgpOFva
GmEWefHJOzlYn8n/KNsPZy+o7trfb903auQtO+fT2BLYeiHURwX9dx6r4GZuyqXoT4p+rlDnWO/h
Y72M1nQp8xlMJGohjEFKbuvqhpAU4ETnCvwWOIWd1RZf91JOMxet988mkuQJ4GzDQbz56Ay70Son
9EyaYS6/4Jg4NMjQJj16JnOGQe9TbFruV6hE8sHuS+G085Rq8o/DQnTNwKNgDj2DjecN6OOo95st
HBmPR0A/jfsDHQKIgHo01anXXOkAelMegJ6ZEg/r0vUZu8Ro7jJhdkgoEec5SCQmowThCFP3wxBf
RiE5QNYKYX6tnhI0hCrvaBfpWdMrCSOkI4IIvfL50N8rFOtiseZsda5RAI7FdTQry9OyXdEYtT8u
zoBX9mAsyKbPaFLMV/GUN6j8ssy0egRfCIL+xgWNUdunSPBg9AyOf9UIi+Y0kNGY48u7QgDYjoCe
pQ5GA+EMVdOe/t0HejP0DKLoEnG6Nszko0amHgH6Wo7xa+7WJsusn3O7AbLH+uvyqvrm6fwJ6arK
PBscDijQ/FCHooxoqV1+KFEU2yrHSLuNbbp4QQuae1fZ2MGua3f+lQt9xFVZU8sR7f5HrAmMJ2B1
OFz6V0R2/TEYPvXqJJh0UrT3ZskGBbJy3X64CrPjc9jdv/CMRL9u9vXddk9sbMOOQVpGvDeX8CHh
kfFgATLfzvL58KPmxljXEkSwSNlX/WHj+qC7OWgcNZxlMQcJb8hxX4t7WwcGlBpnaKXGIzpFoEwJ
V0HpM1nZP52sNEyxSvzeyWB3HteorbXuB3bU13n9KEl1aBWAcf6XiD8OHEZi06ToORTSqC+NLXFu
UipyDcNE1slh6zZEn7RR/dQvToxseI08706KUSPLgIrIeDIoF2H2wFt3caHw2BJV9f0uhtsost0C
TxcWbExgm5OtZ6Q3OcFpPeieUgcvxHcAQ2ffhwT3ICPnrGR6vDL2el/YWDSfEBUCSRyEfbZd3gnE
tgTas2qhqYVVczZdo/PSssru79+usymgC/0Ev1GkPBFBGza9dx9sm2mP7wBjhj1pVVE29+ZyacK0
ZPoljytqAnxcuxajySucpCB+HwC3c4qZ9AzUQGGCPadf60TiYMH2YnXqDib9LdTFKN2k8eDMzroU
U3yYnEWgkh2DGrTOxPKFudTkRc2hygBnkF1Gk9BzEh92LnPCC21bjURCQMeDJmo7G33KAkNqkE8f
aX8ec7Hm/9tbisdFDoaMjPVonA/6YeranxrvxFddm2D02rbaZDavl9gwYe2rBTNxdDkbK22xXu4E
rWNY0+MBgEc60Tn0o46Zauac/M85Jl6zTiCHZR7vMFE8eFSJK9MRQOL1dqDXYLlMuBY9ODP4vlXZ
LOEMKZt/hpN5t2hrKZoXQX2ppuY/hJxm36QBdfvCEe+v5OguGsA5fjKnwjDiEyqO3phA0I30sl6Z
SUuoGDPjGnBur8NdR+26suWnsWg7wmn6+IvhB3ggSjBC4R/TB4WoRnsIOpnTfcBh+kWbFG41n2rj
BQ96OpBmarQz9Onlm874RI3bzyPFyBOme+8t/hkUibjeTveeQ67gxGXScpRONNr28B53YZ15+iCB
paN8KmT9Y7AG+y2fEKJql9jIu/TqH7fA44WaeoVWi//zdPy7kNBm+1F2sz/1a/mhsbh5fZ1ct2Qx
JaPpD3GTSDS95BvkqKwxCuo9JQ+SNyzglUiFoTVKp83EfXkoGR8E7XcSAps4ZARPRwW6eVQmRX+y
mmEugboejwn/9DBp4xEPghnFxYCR4kNPUHpwAX0rwOc+0ggu+Qfs1osipuRTy3L9LTSn1P/GMqOf
qwZ7nrNwZh3Cbrr8v0g/wb7CJ4PMQqiOk5FibCeN+ms7Tu6f8GT7IvLuel168TUl5FJshVJdcT4W
+5Xu8pvHZEOb4y99A0g5kscXZ0ZZe3uOcgqjQG2Cvh7Cr5D49AGSQ9Ma49RuaLfNtBOPIWq/ss1L
ZHJOKfYGp6dAxihndbRAHrlr9ikc2X26G0t/K+ypCn7hBhqsNKryceZSTEUr+3mbqzjeP+qJQp9a
ytdwtispaeHud3zJO6xkm92ZqZEugm5tV86jFbaYl+uI7DcYTZOqgePdF2ivmQsF96RlpqcfywYc
kQCrl4iKEEBLgAK4qA3JxHIz6a1vfzIf09SgBzzTs0v20AgNkA+9zMWJv6YXx7SRdO0Y/tdt36Rc
I3pCxaxtFOl6usmFzq0uFp3e0DzKkkm5mofCMv2QnUFplGzZanEAlqT8APxgVdrHIGP2cuLVfzoo
W8smzw7ET17RoygIXrVWflkUtenZcG8ChZSPxQr9L1uNLbja99i/OVpbxP0iA/LHM6wUMlRR/JaB
Q8bqbBPIg3SAGZ6P/eZwlS8/cyUUM7WqSFHZD78wmRjbwnPHKUmVu3UMwOsZvzsJGJKp/pzRNCOE
5wpyhdqGIcmDsyFnPH0xBXgJ2WG2eIak7Rk/uD6ojrrgXLgJ8mZPY9FV8WTzV1aLki8cMDV4RKLI
BRkHWcJXoacY2XRPGwYlPEdq+OCapijLobUBWPgJJ35JWDshensReIryGIrf92FljfefMg1gNNIx
jTvqdvTNqN5Z5vag76co2pJXIKM9OOJaIa0BZR7eHCNIPn5TNeknwxQUEjs1a+OhpD6aqX+LgNXk
ok0R3D6g6BiPOBADQlY6jTTD6vBaMO4+exbsERvN17ztCYYyCm8UZeupxSHo8vIABQQL0PuCBfw7
SvWYRbeeD0/kChJwQunbWMisBxCovXRErPbuPLlh5K7Xz2AyiVQnh7tXewORHuyMyQtcmchnQ1od
jjW2YFumgCmE3SpRNVCf0IoDLrGAy6ZmChZnaLME9KdeBkTy/b9OHIjCveugLXmUhdOS9aRRNdkF
pvfbt49LPFFun2JGW0ruwMVESaav0LH6qPZuhLGB7/Uo2Xluy6Ut163g3Amd3HSvWtwC9/MabKlY
lofKpbjIDjtb3WXfnHXULzYFTNqIhqYe7FiFWT//XVAiOZhnaPTw2S7BCfwTW8LjiiQQotBliSKn
4yTXmEnsitf6BTirDRRSA07ZbBJVw4vO308r3NxA5Y/g2tzR2ZZ8CUrBPYv/PMXQ6xlc02VRabO+
M6aNfALrRkI2lZOUyStW2t1/DdQ/GcKOKFNBuwMM+CrfcYjvCNAnpJB7IcpWCp/jmgOKSeiWbo6d
oK60PttIioWjJi3/k8dYumAp+e9iLDkF4w/rxHCLQ95JIxhxsTw70W10hrGjU3m7SEaSBHdtHZVL
ucWI2bMXqAFGSYWZs+9RfL+Q9aKHWOJA9wKdg4J5RTQEChXNTAzHnv9PrwNs6vLSyVAo/mi7F9Bz
UhDkl2qTBVhuDbofdL1pHMvEp9Op5jzHt6AhxaAags0Q9iUkeZHDFpbact7qSwFIpRpxsStEw+Hs
L8acXQZwtUrbWNkVY5VbH8uhSw2PgjPSTTi1bgW5siVqzijgXOrCfZ6aNoRBaEgQOf7JViEwkitL
dftj4nNou+aVOrpp8GGYIRrkUbN7g1LJOuYi6TUu/56Y1lGVLBiHenjJsAVBh3U7UoMDFkkBO/9n
BjBH0FBO4uLRB1Ul39BDtJHKWoNJc2yeF3rYAsH3q9dvnSm5VEQBsqKPVXcfUKxANrwDdK7C7Xxj
AXJZnb1099Cadx87rqKGLpJtZkiGt12VeeLTLyUR0yvuzvcLGG+fvzmE1QLYN5J5py1w8DDnyx23
w2OAqGIci7KQM6eOfVQta9PxJenNdy8pYkIn7r6NqxS63RJyibyRKqlyLQ24FciYRevqafy3nxm+
/ntvMoUgjQRedeg/7i8ru4qXHfNq+aeKfRuN1qJ6vTSh9atpZKLJ6tLheVG822d7KsKLg+N7CAmF
AZlmKlNuGq6Z86sBQaUB+FsSzR3agp4OmwvFqM6rXTOC8C5u4xlrJFd9d+60trp/7bM6M7HxUXQm
27sMC964zT609347IiA4qIbnvvzviW/MQCv4FacFBOOzTo+eNTjwe0/vH47PK1iXItfYHUZdrUV9
NsVxLzTcU0uP0AwuT0piiL42Q4ezeijXNXfCnqmw8ZPKK73Qpgx13uiUJ6A/INK8Xw6y5YgbgZIr
aYno122Vw7rTRHJqnsx9YO7DNYXkNQrI3bNyLI3mFXtM4/u5m/s/6cIPjvFh3G6BXjA82owpwgLE
Az3MJPrsm0J48PZuUt3Uf/gfyNysK7RXCPLv+4CPqZBbWVoVeKo7okW4Z22nACFWMXguQa918AF+
QU4sRcZeaMmnt4+QvPVX5vq+ETFi7OGDBymxHZFdMnOYygT+lYPlJIHmxu6Uql7Qruq36Mwu2N45
6oAW2dmWZqW3Uc0hC62W5wOjBf52ce6UwGPegwWCNVDGoSo/ggl1s93WynsTW9zKClkji45epnFz
0IPRiVIwqnn2jPEafqpN081QkUQJULFrVAhXhJNjnHeeXy0xDh732u1YOEWEsbSIE9Q3lG1i5zLG
ovqjf07a1q8HEQITYe8FsCXVUId8QDpAuvqEg/lRYYHjS0//o5JP8wHRTSZSTpqM8jSamFS9OJuC
naHCrvS+HpLKcBQLlsRvIGMWwNSGDO3MxXzLNGJUHxsdJDvqs0vF6cKZhmxpfehrGpnSxaGkEZw/
3tG5fCNdO3GFjqsbkT1ZSEZFI70KkNAEiaOrtt2KArDF3r5/dXd4yXGF+pB1Khj+4CQZfy0wU68/
GHeMYFfMMxqcBg8Z9YwN84ClQb6KQU7zjfiCDIEv1zZd0OadzEM2U2YX4Wlb1Nf+/PnRc+YGUmeo
nRspm0A6rInHf2T4cR+p2sfMuMVghGl4O2YmUDwbSAL+zsMoxU27bB5e6uo6A8wZ9rwGzeb4d54t
4mQ1rlnj+g/azIeMdmuX9WysHG/HHam3RnKxlm4HhvtWTClW9e+OtD3HtACsMxMdDcV0xOixlXBi
44ro+Q/bf601z3SQjRTtC8Yet07tE1Uwit8p0fgk7Nl+XrNvHi/bdqB10zCfrV2BhdL+/BvqRkMs
z1+jlPzMyj/znbQLzrzWtn5U0zJrWjitNWGJBBe2wIgL88CzNaVc7cFfXRyXCqkf2/i9bWiQMRd9
AwlkcD5xoXjhYQAYDV1c9uW2/HvkLmG9NUp4MC62eBZpUdCePoqjGYT/MnuO6rFN/k00BCjtfRky
vVuvQyLpawql8tILqSW7QPrDXXbytH0K3K5hPhiXjHxN8GuAKp87tSV8pg+YOG9TXLSX2cSAqcek
ssNyYbxrW64YsftE0WShrpsZcFDB3wVP3R87X+BfaViAEKSVpLzP3cEOrs2PQcSc4O8JlhgSQMUr
HV70Zt5hShoZuodRDDuW6FFaGZ/peAL2AtCkqvi+78lHIhblDtdlPRBF4rjfOYF8o7SO1WVmkwQH
RLVVkmhNv/rYX3eF50MFRvk1MnpApgmym2IVUQxr+GG8s7wClU1WxaWZpmKhtCvxObmIhZ+B3ZiK
03g6FHXpXdg/CKNwswYseKZnE1wzqZEkAKfShie7QdytYISkMCzsIP9z5Ku8DfFu1mRI/06NSIBs
ljd6CERkm7HJlsIMakFvp2bTVHDR8F/+qBgroPut0ZhqY/0PgO/PugKuw97e8hFz1oXdYGUVHl7p
GM85lcGlOEO4mztccWbqMuxmR0dFMSevgru7Wr6pee8XVyxQAVlGkvf13HL6FgAILLnlWXjsHuIN
fqxLNo6GWXBam+2NBLKFo0tIageYRpV7wWc0qB64YicI2RPVJDHy6tZ5a0kVUk+Ua9RgQmd4p/lm
AWyK+zDxiToe0fsft3YHGm8MHkrRHPmQIOhO4HqII6DVuQgflCMtvhfQnmYYiKTa8c2ebds3q3yA
3gAuPC25hYdpYgqkkXDIRj2sYq/qHUvxC4avTGsSSCxnCbHABt9BfBREeqgWvSzZj5+mEK5Cm3pp
BeYcfxoEvp3Z4Hcj8CiV8i1eRY7BfzTjeEoNW/dRwRwBOjjhuAVOj7PqsHyRsdMxJmHqUy2Xpa2q
aFTjv2ELvXFtuIDSRxVPu/8Nmb3LTvsXaRBap0BreHpOXTB75bYbML20JxJuO3u8TRcTjfaGSowg
fWhpK1TuDp2yBLiWaFgeQNfHfWLjkEIeRxXsMIfkEmwv1Ti+v6qgVGHg/TrhEfaI/AaMmgxPEjbj
vRveCPXKo5hY790b4zIqRBVdFvZqDBOjd4JeOI9JcCxb/9o0KtMrE836kMC2ktA7HHYUPb1BloKr
tXIPEO9uzwwfAfSPoZrtThemBTnBC5amHiHPxzX6JBse7qe0xEhEUTbzM36pJ28RBuwdU/2mr5s6
0Il0yFR3KgbLEZ+TTRF987JtluuDta+02u6y0w3lhd7Vc7FYejwXkkJznm4dedBfqQfirJZva9o/
5SlVdfHnHnZlR0Fs7xjwbDmvchP4+BqSutzm10RHmpNJJ4drXzn+jvVYrvyFearZkLwo4A0z1sIf
xwPIQR5wIIMF41C3X+7cZ1dpPFGvS7D5okmkRlZeoSBBDlxGT3bGABZ3+V6b3NFk9nF8OgbkxubP
tsaeHzhNl6WoLFjSmZS+M8Gc6mE9jwHvp7lVnHEYdROKXSfBdWH8UaxSyKg8DEvf6JDvIrdL2mVa
NqVst3GbklXNU1hSw4DSgWWht79xvrJ1SImUAKwB19olVJ5uA4p4GWuQ+0jwFmWOWPOZURWXa2FN
ofEf6spySck1LZ2dZsaPsfAqw5So3I2y6HN0NhPDlDMv+WjAkp21BYNSUYTFQZW4xl6knqRFzZGo
NNz5gExxyH+Q2Iyc3HWREXxEYRjPJQqj8nGiwyiPt9xDsxYMJchYT3fA8LC5hT7OTmLj68CcDvyx
5jTsWmFSriid1Zm4Mh94KcfowIi8GaxEhWluXnR62LtOmmg6SdmS6cw47lV5VFTkB0a0ipNAuW6N
I1hVegHCZ+qw/ks/gpAC9JTywWnCQ0x/v2vmfleutwe5X02qdgi1q19/OgQf73KMT3FnyU/zTb4q
k5lbnlrZwOAtqV64+9xznyay0/Ytm/9Agr4+PRq4+aH2Y2XAZ6bVAsdEHKjCUTIlmMjrmVR9NgMH
Usby6mrSZDFsu7sJBYbHAwPMqx8eiWT+eTVwzNzaMS7EFcEm4xDUqdpPU6ujmmwayespMOFpuXuC
xVZV5ZFfrVe51Mr+dGivSI1zW505pHqa3Bim33t9iMFmv52C8YgbbcOuK8W6sD9/9RCECdqhofVA
OyWjryXLL6zDQPdcncGZ7sr3iHvpAvXR9hXO9WfRmVTVdz/tkLiQGxLNMNtgob/QnK/OI60EtJxm
16Rn6S74FyQHse3ul292tmb4ufr+KPpS+ZGEgQbM1Ti4v3x8vBNilLnWU2cC/dwgFchZW95m4Atp
EcrmSlJrXbaMNimHOKWc+wkvXv/LJNTQgwqfV5yDQ3ykMTtjvANf+V4JMaGo7jnVJDc9C0mtXCnL
GZl0lYoxtANivGQDgTiSevzpvS5Se2vNmsXGlXFNWTDxv+PU3Gy51WEmgLNzoy9EP0ogyqzmc/Tq
qhqszKxQRl63yGhHtm7PjO5zbu3YoBx5JLuykR5eGvNy0VN7uuYvvauKzFvJFZ10isKIwfbFDDcA
hnxj0UoOBLEgllN7weLoD2cJP6DAU+XslJoOEaX5KIlMSrgh1e4V3LMZtYtRzhaYF2wFXYbEcF9S
zXBJHDh1QJPMiZ09S5GwIm2/UAcVHL1A6nMHASywHr8WRg7LAvMYqQnIt4s0Q3560sFD7DWyP62D
uPtzGGfbzX73hGIVPh3K6QI4NdjBYlC4nzG12jd9lvzMvNlzWmtNfY+U5kHKftNEQYzqxC8E+HQ1
vcJfNx2MoUn6mGRewkEyH+cinfCpiZVtolgfBNkq5gaKIwELjIMOrzP11fRsdemFPe6ESEQwIcmX
Zwj71doRB3zxCl3NThfrrcI6Hj3U46ftK5uz9YZrPUKO+7I2NiVpOq7jF6q+J9u+yvDLHqnLNoJP
+7UWssPjJoWg1xJLZbXuTUNB0txprPWg4bgoHT7l2kPN8g+714knpsI45oV347eqb6reDg46xC8R
mnrfQSN4HN81GGpjbXJ/PuUFShQEFy5SK6XMCQC7zoyUhJbnSdI9WRVNg4TC15Nxpmny7i7ocAbM
NL17B+/juBMppXHCx2J+bsFod5BVLdSqa2GGGX8zCSOohMy5Tyqp2Oz2qPOwUm1Zks7iXGb2Vooy
kgYfOKAX2xfJXfRasP4G/kS2YK+u0Ltm7CNI7kWswOHjlT1v6XpqDXw6Wi1o844EsVKe5tChcs7U
ku3gg+Pzj73kksSv9LGPykYqrIo/lNcr6amDpPHeRgLWG5xxBGA7Vjk5Po5wNHtChRQFSO1kNdsG
vpAA9lnJy+agKZvFZqBQnZSAcuAqxVZMtktVx7JSUDCqgCGqe65uztc303hQfitnijua9GqT4cHE
kqjqbah04h7BjYyvQHGkaE69KZys7q+sN6bDy9+zhvFhARfSVxEgJG7qsOmBCZeyn9rrRMHVYNDc
yU71BP3YXDm4i/8nQb7hYZ8/htfJSU/VHs5G2i4ZLc5RWBgX4pMP2NBMSBff0k3WaoVEDIqDxcZ1
6UEniFoKoQEuO4gjcYxWJuYPvZglaAUMR2lJJVv19cn0EaBnZefyLq6WvXmnvZo80+F+sbB6dEjI
gxshOwywR/G9TFxzEQuViKwvgleyj5UotnCHi5hozc27EQMQtuUOHmEVb6pDw368R4UXCImo43Up
zPHOSacY/x/sq9CokvnF8yN1flvVj0OnumOKmbkYfI6CGv5+VijdwCUrEYcfzhjCdd82Vbh0MA8l
9WQRocssCY6veqiJ5qHjLsxBBjVLU4D/xh3Avq/j6PSQn8aPtztmQelJKS+FQuXfFSDvsaMJJLmG
2Yp3M2GndJ3NWjt6EbOGxKXVt4Q1a+B+JYSlMbfUHx6yNNSnFdoT12Oqm6t3OnX9Go1pExbL20rA
QPfpkd+MO7iUPRp0H9+pBe3WbClfaXhLe4FGZ8+spktakUjkuvyfiMROiLEeqFyfHlmIEID1V0O+
xk+zg1sRQ1E+suCXkqZ7LsXWGaloemfmrN0Do4QCBo42wWksm/ZIKgEH1eoIAXF3MRrEgkfpOBgq
4+NNYeHjeVV7Y4+3Fkiw8Sfe1IOz2TmTRx+1I2JMAaFJ2YbSvrePXFAIIV/iE1Y1gCN0zY2PunTH
WPebFZC7M96t9sFyIWAFaS+fv0Fpy4MAgZHRK+mFWwrL0HUPC17rMPMnxnU1dMbAGQ8rXmnFCXeR
4NTbBJ4+K9593A6XDT4hr5jmtGvcy1xgazbJiNUMtkWrfcePIQmFj9U6oP6vn7XbDDZ3RjZHxU7s
lGaqUQYCAGcdITNA22Qdis/u6OqGSe+GlQOqz/OwRwU2n+sTaPrWFzV1fn3+Zv0xe/sd19JB1v/j
VWrRLs/i7UNGUq+mxQWdRA8tEyHpzxpqLLxcNYCHXnRYZp3Q+B3CDBmQBruJNM6B3iWFavgC+hl8
2pi07FkPfwXYgdaYaJsx8uHUOO5PFhHzQ1waXEwxFZqtTeO9jg0zCAOdgYl5bwry5gJZ0hEpLHPg
RX7Hx4137mgvDP5dVcUbQA06OjVgNRXpzRk40eCi96jvXmA7s50tctcnPHv50LIbwXyOIT5jVjUm
C1TvEckruI0vvnN3Jlugk0qV46cK6IhxvvQ+DGp+7RrJGpUvR4lN5C1NiVtz8yhh0qrIG73k+hTy
kwPvfOzAzPKtORrH/HZUtbMJZ1XTgm1RfibX0IxEQSnuib097Qtd8B5r8H+WGSv7aKmw6fbxQzmU
JFzpiAujdT7L7tJvG6OgTOlR3t8jzTiHGejdtoYWcmZfGxv3UbAygGEfqGWgRzPdUPX4Oy9d3Uk+
IJyUbCQ3EjBNFguHbWFnupTwyT9TuX/0MvmWlc/WSziUE+SSJqlcPepLNOQaUwqL7jTKpzvvJKBh
Vk0Bfj1t/SG7bsUFb3r/4uH/1lM7bAlqTOo73fkoYoZNaBhjb37jA4rwj2NNsirz3PKssRqp2/Jo
STeU+Sk1NX+TCypLPjlI9kwV6/BeJot8aUtPh/TR/Jx6byrBPtD9GdnnnXB60nG3Z0BLDaZvRjGO
z5teusLXSnzTBbMMmo4nMMjibciI0L2rIIfYzwQoi9okkD5rT63EuRyCK0EcnEmErUFX66eP860j
iZNiJ0XBxpjB/Dpr+y00YbWbh4VFi3yi9iROxuKXp/GuEVTFfCHCw5tgsbIUwACfvdEJMxqm20xc
jMu/NVYfHfdcDpWC5cYymzixFA2v8Wjvp7i6x89Kto/CVmZxAU65R+3SXwZq/Y3slycfU3DL8XN5
ff7A+6bN66CIlKLwgGTf8JFXQWLa5QoZflEsVRH5zHphs3lRc83jzHred1U/Yv3qoEzAv9mP2Gm5
FQQT0oQl+CXUtGcV0n1mbYVtZji6SHSPa4StSMpS1VuGCZNwUp7XrPLFYNVW3R1yz5SFLKIvycgu
bsk4iQZOC4v1ZHiq9y9XAJzfU+FKaI1e0urRidoMb4YoJjzklf8rUbvso+OEOJo49bQNYAxEURfh
929QqxUFkFsGV8SI7zqvNioJWgEyFCZJafG9vYQ9Kn2YzR14b6PT9beIh0ve0tYT0iy3VNUIIGCF
qXYe5Stnogqy+dmgHU58Ij8/4lnoeVFayivyxEKf+fmtBBsu5DR3vArRd2yEC8fcyNCDrapM6MkB
G3plv4todK9PYSU9hB2CGOYSi+wChwwMEGX+TH2KX+oumnqTYfHqaqGPa/y9MB8/1J9jDKX7VZU7
YWc9S2OGVWtGtzNKVb5pMg/CuSAWHQ9kcdrXWABH7W4byw8jqPhuaYLCoWLAFfcmYp2hFhlK8Jep
TS7TxqYBQKHTLizLzS5VufbPR0eNNIIDZ16LleumYSBq095mQ1RDgTLH/h85LbDbblSdKAidwN1D
pZEDMaE3qQZjQ73S2XmxzcN12pEqX0CQfknYcqjcBnR4YM0srslZJj66us/hhyWi7EIw3PDcENyZ
509cIz0QslqYluoC6o+gzFpbmtZDTfPL7u8ngJ6eEE1jl8L6zIWb4x7TkA16mOe/a1m7uQaURZtj
eKqeBuNQRPw7VAI1Ok7eBNNtmX625/40eznDRYIdewiYQRMGvD5BVb72X8+09E0lFq8bYalohr1b
6jtgBYy5OgaXNxubr30R6kGqCn/y605WLnTrJ1IKoaJSg1eQTYLrCFucQa4o8+098G+fle00blRZ
QkJ0ou/1SbPlSQ9iWobzkHdXhHxa1QS99lhq+cHxAds84Ztvph1nLqs/dreOxX8XjbJejDsfMDch
c4H3RDC+HwCz61OHcwgkxjn4VW5h+GZbOyyHGKdxPSnaDvtgJK4nsTH5NRld1S4RvAOUn0Y8iEsB
gJR3k3MM6VZeJff0zdJG4qjgx4QZNK4P3YLVphyJw+00ugwcZX0nMyjodEhdue4v3mBoDA7KohqX
b9hsbZwDGIwuaj1psjU5exI8J6YD74+KuOZU/ommurpFhqLDiCkfaEvH5NUPRBFEHEWNKKEgWaSz
tcMAckTx5jf7VNVL4pkBn33yQoukmv26AfzYXa46XEAzIIyXQWsXyD+VxuRyZG7xQQRkJDVTCr8V
8dJWqo9NSnX0u75/9Fmm5rC0py+auumh+kc62U8MtqU8TczGtqpsi7gHz9/6NyH2r1K43E3RP5cI
8RSBsAqyk2OibXDfQHb7+lnRL8lUnqTpbxTDnG0WPynZfXjayPw8GGK4+fuzg5GxUtTOpqGJDUAo
0TK+MGjuTJJDfXK2RmMmKkzkI4zYFSrf/W0Iqy+6rSCInxhl0vfPz3T6MhzP/y2i44UWERFx99mg
ubg2sKlxAd+bL1pDhgq82qE/EnWGMY9lN6PHW4uE/Jn/Ql7hmfH6Tkfu/JViMrlirA3GRePZKNTB
8cpGUQXUVqMtUhtRBSClSNX1IoTR5nGY6uFx7qXx4M32D1qxF/tErAW6oWvVg2kmV6cyJfnPMBdG
9SU7hBUzculjpBy9opdPy/gooddexLYgEjYp4iW9gNZ+CqQf7VHv2JNAki8Q4R7+gKjl635p740G
JIkIuBQwp0T50UJctzgGs1AkNt2N+gwcg0kcRBg5md+ceK67SLdqJLmAxhri/D+QHpvvIMwrvF0x
ixckEkzbt2gmqoGAkgGoYknZH7358qIs/5itBPKE4s5/+CHP3Nt4A/0kW+IE8UMXE9hM944pXSiw
VDZqH3nwejGkQH4ISaAEIL/VEW7m8WmptbP/4r5rxZHE52UdyXJBa9htOWK9ElLONhbx21E+ub/6
GbwygwIN6oSDrjk65Lz3pkbtrkchkkQHAbWNJXuWun+6K268H81J3pOQ6AMk0b2x493K7urU43/T
cKbbypkzKr2T/uGfXidIyiY7CUIwLg4cfrcIXLoGoA85VpOGCJ+yFnKR0w3lofTorYpaEGAE4HOH
98tp3En1jfLKahcL46R4zUKUWuszzdqUE3+bPkWUiaZU+pwVDYAsOJRQiVwJKUcRDYncrkgwYeSG
BXVd43PDn/t+k+j9jqibjFgWCtJITZ9h4Ae76JKiMNMjofRQi7LXUi9BGwC0vjuF2sUjPU9e6J/l
6CVLYz/sWe82XXt17AnxVdr7Rr4tZO/37qz3XzMqBGfnGZbM+C6r5k66OaWNy+EMzkVA1X5oK6On
ApIeZMYI3ZuJAvzcv5yelr9+fQsUzWrpSAQKZI4yBPCDsjnS6+bcOmN3lNgVPKRhVwd/ek8fqkRk
cYCLQfzvyzWurr9XubAG5TF5rqqCi6T79VeHj/hCerQXRxQs6CboIY5lDNWAbPAH/3NKFWPAHyfc
wxmz/m4eCfmby+x6BojTXYxvM2V20JBfYrpKng5XuWp2IM8Uk05s9Bek3+Y/xSWEm6jqcaznFLhy
zXhcHQGQhTb1O6PAYzy+iuTFrundnW/Q0wEEG6zfxI4Y555kpvr5WTWfriwk3JyfqVWGo8P/iNmV
SLxjWZkZu/TSiroB1WXCLG0JpZjxXGJZ/7XrChYOLvtqcE+SbJ1gYURJP8UT2/LXnR5BFrJZSJri
YZbPVfMBL1oIZidL2ArWDkgO4BDcllYNV1mLdw6mggpcmp3uG4X4hNF3qAoVmTtc21sQmdTtXlMq
721itQ97LuF+8wBppEVwhXW10+GexKWO3GdRCF833Bt8hCW/KCsitEU8Nrlibfbx/ZYKuIazCd3T
UbZK2QsePqkr+l44CSVlR7FIIItvWQa56pEkTRfDtT45fuSKJZZYrjcu+CdvRG4lviR2nC1xd0o1
TI9/nrJTzXldf1+4jA6YMmL3oVbTf21U/0ztHXdEjNFFDaC3LFSUfsb0kMNHi6yxn+Pk/HmjUL66
qGB5St3ZwJB3U5TJvk1zMEBFlpw5HCgJlVZFyGcwuraCUQWWXW5jPyYqjeyxL0ieGeoG5npwltXC
sYyXv+AM8kU+bVfXWzwWCsaXG3NIPdJtUCJn+m6aDollg+BSL9vmtCOQ6SNVPQt7EUcff7BMGDUo
hOesyr1fgA5/VECkNSrkqrh3xkJRipyZYSbTYHz5arbB5Okx7NpGlCjCNKulOc4+WGQEs1T8ixJY
wN33OpPRtZF9rpKA/WszGEFlfJQWsnyW9V7YS/304zZBJibz4619iP1MJcwSgIgPY51jLV8R2SW6
XmTbj56WM31KG4gVrqWnAdGn6JXcUtubwlQc3eioG9VoJ1nqY65piOXcJmIG6Ku5aY5FJiCmREaf
qopoQnJ4HtXUar5wY6V+Iu1sctoVXxun8qvmGHokNLwpS+AfwUm0CLB1GaY03VGKrNABjb7e7jIM
3QmTv9fl0joQRBVlVKd0n4MGThJxmxTj7+py6v/ugGVzJjTHb/sucCIuvjNRWkt6KIBxMysaDFJ/
LSym+xBZ/wEuDViG1TfE9S5hbboaJq2lAjDwo/LkFpQr7POkK4MbIBrr9zMdyRzP+H7daa0P0R2J
V0DUNDp4VrGoBfTKMP9OwZtz923NzKVwOb3ARXE9WdhV5cMur2Oa1Fpf3aGKLaUHEf36Plb9joUs
uzNAIZHwwGsH5zVuAYCHO8vg5ZMxos/9PX5GRxka9eZxS9cigvCKEyTXbLxzLNj1BqZ8Mvt0w15C
D3l69v/nn8gfLVFHXQuZtmHM1PaBSkR7ry9c4jDstQ5WG7udrZ/k1ZcqRXqwmGA/rxk6Iu7RZw1X
m7kSrcEcAN6yXoqmbLE2w7+dYMCk0chALhiMq+BIamQbNfzib+ahBVIbLFvtfm2BS29CJdIjVgnl
3+60kz7I4vNyJGOhU4GyxM4R5hWNrITs4YQ/jvfeS6fWwfZtZGnPe+++Cc0+ybLbKtI1ynbyMasf
vJUuKiaDzwsT4abTYEda/UYogfJbsp9ckrhgRCIZxQa/MirX0acfs4ncy4NbM0JACqmoarB/Vnuf
K68zvWti3vMcM/WlT+wxsmcP4omdyWCgd03sFpP565oDtmGKIqZDdEnGV4uZdu1iQmXVamMAPKjv
1deyPUETD87U5awWFMiH5ujL3C9XJmdLiOhxLhSDi3YtZjK9PyFiwZCkQOXNBw56bk17aDloROHA
8F6wJLYXO96jWh47n5kZjW+OrLHrqoE7QF7FckpXbSwOXC+luCqaZzWENsM4LYkWenA+QZ8dSDg1
xd/o2Hr3utM99IRjuKzoBZeMXC8NAbcMGl4FvzqpWXM8rZAz5L66jBiOHww3HVAFuGDWQ0rVTkWE
eQXAIUB+gFSMBYXJGoHvImmD2wA1kt3o0FNudpJOcBO9gMTW1Jx7kG6IQidt1WQnCDNBJHO/vJAu
y4mjg3fqDxgG0MnfKz2iI6CdFNud0CMj5ydccf2rtk9zrYEHryLeBvZVl/askz+apAsWxl1vdcqv
PBmIgLHj4GtPA2JleE5S9YSiuWG1AHtLTPeJqw6SHRTL3BanGJqgxlHDzr9OjlVoK6UaNg1ev5ze
7C8BEr210Ni4oyKuwpQWA2cwNT5dOX3vEplNj1bslcB5u/jfD65029vz53rNz+MpDXKYGXUM5oG+
fze/4HyqeVoL3vvhS2RXm0FDuxCCQu70rynDB+ONdEfO5v6CYL8SUC4jLEz/2p8n0rY8UbInkn7Y
847rFkC2IeT36gvzRPW35JOc/+7KnDp9dX2pz+BRPf7y7aBGhopRP82Fr9+55JC7agUyJQBLoMzV
uJ04P1vqY8Q6ti3x8zQMjyQ47MbE7zyt8GAZYfcwE3r/a4GpHrJTelKg2XTh3wAyWuQefg/bXssB
8E3B+Jbm4//MuHrLX4cOSb66w5zn1MYz777MyybTFREccXvPXUQN8l0f1EJSMO/ySlv8ldfnqk84
MNSL06oAcp2YMLJiIrjKszvbCE4ejoOcgusqAEPYTDeypukpMupUEZXouFRjss3lM4Hr6aM+e2io
uogd3NRIv6XFaCEaUz7VmCDMNZ8n2EG32x9jwDJ7kWTP+Fz7+69jeruqHajjcLvHn3TpChOOcpvE
Uv0Sv+ppqYNQuHY1V6GqMyjhW909/OpUnKDD7gfz1Xf8W1anUsOyS5lorAbEvuGZ/Ftn39I8/CZX
VZ+bZvG48IW/gV2tTO60mbJxKW8x7YhVakINhmAXeH2ZMa/5FY0QLy/oY3AzH4oDclA+kvz5VZgj
XaeuQ9Bi+tHrIiwHByTUwxiG+9ewQxgLWyYvpfYR+SoJfm60d/8i1TdGzDPp/syDgpImawu0kB2X
wwJ3QYvbp25RXlQ8OFcBhuNdMZcfcFV7uYmB1cbaLcy/bsBu8icHMQZRh8l+7MQB7f1nLWRECOXm
3GzJHVD1Z35MOGeyeaCftAczugLJAvzVdwrkKLpmkHCJmuyFPJB7un5IRjJLMuZigECeAKJIrTeI
y4nVQfpEo5RQ1ImrQqh3u5weIpwNHSxwSLW7DOf1n8cR7dTBmu2HlUm888MzdpKpJXU+DIGLLO6p
bA2sYi7ZtsCSsmy7UEeEVHgFxbmAqsXop0gtusVbipFEUuHchqnPVbb8H/Z8MfZ/VkS6Swl3FrG1
3XNk8TVfrmdTFxZwFavf95LwfHocir5dmeaAibbBeywF5WXSG3zIZYB6DlJqL0vtuoi7RuE+W1mo
tVVmA4BwfuDuYGI6j8fJhCRNQJH1iauJ4mWLDdLCbHx1YXoL6jdNvhpacgFXGZHOoXiXqJrn4BGK
GmdnD4fTiiONxF3dzL+qQQNGeOK43TmiyZepTnnfJtmynhngG007gnw8YF45yuM12FytRut0kgW6
Ba/5ANY8PGSH1a/wjm4Yo2VeHwIoRfe7Bh+TqSc8XNlFxOIYkYEp6Ns8yzWDag4/kMXUw39AtQuT
ycn55QWylpg0anJYY5wOBiH8/R328Taj1dyeBcNwyGjHKDBS6PK/sq/8W6eNSLhwSCHYkjMagDK2
AePRbZZn409M7N2iR+2v+5f3orR2Zqx5TDSY5PmYc79tArsK7KXT4io3DuKEhu1ayso7JzSWx4ih
nfaimBUfO18qwNIbUT6qmo3rbDPuR+jACYOfNqVTE63tFfjUq0JN323kue/TUbCq496FoYwCBId/
MTd7Gb9ZYl2CenFmUBa8JSOMF5RWTzUqSBG1ckIS6pwh5jXbVr0NlDLUKu9InLDnbzUVaciia10F
QDJafEFrTIF3Z1putuobrblKCJNDH6aMlOU1lJwcFUt9/AglekXwC2ronqjcsbOIB2vfk2ZZnYyh
kAZn+keiQjFzqfJKaGTDC5Pm3m1CgNUbE+LGj9gb4I67iM5fOk/xarZwL1bqhV4gNv1cnHp5j4fL
30eaRUfOLxeg92/FrTU+giBcvZzW2MLMmVT+w7on5pGEMmZXl2F/1/UbblsY8ylBEcc5WAeTLJMd
C4hsyYF/7833P/9ZUA9Vschgu1Q1w/eIJgwxqtC5IImC5ytzx2MOJh0DbmztI7tgXibR9DBNs15Y
agiuGjIRpnomdhkiI4WCm6ZEEbrWoPpMGzl+pXSp8j0Zm6p2xEqztZJ9MaStuHNR8oKnkyqJLWvy
++Z4VWKVLytcMybt7xZ7dwGx/kzel4LxLa1CsoCrDW0JwC/RVnR8BjYx97NDZAgpy7voH/gQlmbT
iakQGh2slO3cCnaMdDbh99PS6WYDeRGryLNsChY4nbU2TGbEFekib5v9p7maeZeF6JrTaaP+eHMz
Ad5+GWKTd6tgM/yvNYPg2PGMD4UiKU3gEDfgqLVOLzxhyu+3SVMd5+E2WAgzbkcU5SeOq5Nokn6T
LmO5RvsZGzQpBcpB5ESYE8cZ6TxkKd0kB1IRoRQkOzyP9Ku31IQ+zzncvc9nirAUwQQ5V68ZGgwe
oXPkfg2HP8gI4f3Aj5g3AtGd9AMWTs3e3iGdgXx9NH6fY6Iflsj2WQ2MHwFx7/CcC2r5zrdh7f3h
dE4uyIfGxbsowszUxgXDTBKishaLpVJDiNw+vZVQMK2wJY21HcHBz8ymyEwCCM7k1wlog0hO2CPH
eVj70LOthwa7HOsxkZrZr+iXmws3bzGsa/Nr42MAvaSZkAEs3fWISWTVTt2yi+wJWRs0h4cww8Ss
0uTtVHmrNnDEI4XEylwhGlvc2O0QAV0UFMoyUUGct8Ym3s7GrxEeERza8Xscn28Ti+/XWtINUxGZ
R8PmSg4qNi9c9jngVTPidm1cGsEwI/g+kG5NI0sUYsg0ZaLy38KLHU3ORlnjycrW70lflwkt2m2q
GTNlFgqv8W93RhJW1OQdRT1jp5+ALgac/kfQT0hvH0EKn7xBwQBuzt51onM5SlCX/V/4FK9mWWiT
yEqxpq2ZITcd9i0B06sMUb74C/J69ALfqVeDuhNq9PIq2hiZMBJiQqexQVfxXbibUibudpffsmbg
Z5rlCblNhxNNW3CRySbdALV/M/ml8YtF+JldJ3v/pFP+BY2iNNlMF6FnEuer5ckGL/yJSbDCMsiC
YQl3GuG067pySQalay6EsWkbhKfORT9GS6/y2VszgVkHgoM2vHSi9prfKhDEgaFDVyfEk+d2KpeQ
iX6eE/4W4ZxnU2K/VYyH9VneT0KVbeS6CSOhOG7q073VRUcypeDCdzBsBM4sBigjA3J7vS4Po8ay
PXX09gDNKUt2jiXgxhsYyxK1kljNejQkgCJlenI9qIEhDudt90NIYGbG+h3mVzSrfvOE8KrG3sDb
EE696W0diCbsK/LC/3nPkNIYfSrU/O0ZgTRPEeAiN0phmtp+336B2o7+wrQ8sOK4C36L0FyYFbId
xkPiwG/1BKTfnoZ533+lhHRh7Yx37kxEtN7tgUT7LDh933ep2XySUAMwUpM3idxc1Q16CPmwS21w
w2WXzG/apKc/+AhhUblI6x5BoLF6r0n1wZ0PZ1UIDxI2qjDYabZhRQqUhaEH1Q1sgiM5tE734Yb5
PuUUVsKjBoDfR+k7kSn4kT8bxY+tBTcoqCnNVuFjkK0zMo/GkJ964UGRdiB6fiRjcWvEQARSPBF6
YO33yc1Ea2GbhzQTFwov4FgvB0nnfbWAOJG7YcuE+9514KNz7BzIF9GDtutO/p+huc2SVu/KderO
g0rDLCk5UF7YgFMBikBntdZoTb/ubCaBdnxmxM/TJSF2ZXGyEwXyaBqiyDAlIP1X1lGPTlOt2Eln
0XIuBOJHakN6JOXJrHGv2s8bLLTZJ3niYQnxNPLnMXfp5dYhK7ndj7/wxIYX8251XFKyNdD4OaAa
DhUkMujEj6SD0/EOdxeasrkzQhSZD6gdDMQ7uF8RP1RKg38SdN3YshLRsKGPascL1X2JBl/SUbk6
8U0fuUjjhp1VXLh7wKJRYbblsREEdw1JQ0mPzySKURyQPI7W0l7D5tn4GOg+IX60ASvBsGPDSOZs
BormTaRHNKQsQilxa0cIliIaZeOaNDeUmZPWTsRTqK3p5zkFoys745B2udopuse0GA7UuwtDq7+R
h9FY1bTLA+Z+4XBJFhXluNg8ew2SHlVyErpraU5oIqXPvsl3bpwPQQHarcwTDYxyeJ8rNSntRowz
/PhLjt3qKLqs3q+QnhPNuwcBq2q796mw0TjrXwVbw0Gy2lI2Q7GLNaPNQSvjBQ3TgTeBJgSOEjSI
EYJKJwWBLiU44aq3xC8kwg4f+Ks6t1itWTRm5Si8ESDVZtaisIzS4PxfRrUwnOjrV6VCXXLczZCO
9X0f9A+8NinnNjkDKgJV5joBjbGnZZ7Tz3sFfmw9DDKyr5u4fttxyoergELzB7O6idF7O15Gm91g
wE50zxMtWgYAZkAYu+GOMJXGEkvtYzdSdhe/fq5/nK+WzBdgQAEU81lcSzbdpzjvWHvubgfoJcng
7w5URAnKDPE4XdaKYiZDIWSfaotUe6bA/SRmUcoFtsSVIJCPiorO6TnHPL0N6GtMlRBf+EBCNxA+
2aDGjh6F0cGUwLc888RY9/znGUh3ZUKGAxbnIwByayE+54+i5OMtesSwC2hSPUfQBNzZR5NgbSJ+
sDl8ozG4vvrN34a45GEyBXn/SVrb+1KU1/svNrA6MTb93Xlo5+cKihU2aK/nyVGQSR3fzse1juu+
hs4CKvN+HOFl1lCVghix5FcnKgVt5h9EcOhG9D2ag2/MJoJJf5zrSKcBHW1ouRJRkXBlcswlyIL1
ad//iy5Oqe5Vw3PRfPfwUPAeLNhb+nRudV1noWwQjGByPzWc8sV2xD+6lg+rPpOtXfXfcY99En/T
jnHJeZNBL/klwiHRilsHHhPNSf+8WNOmTur25itoqZalmB/kvRVWRoxSISdHYLXSDaNMPD8eYHef
nfzKSjERhe8cglVv8bReiGT2Hcka4/0aqzeHWiwrRHGzYAwi/adFRDMRVq40sQToF4nCJtE7c+Wk
9VSlvYHZbbhnkfLLfn72PcxJoxSes81Eu0BANar0sNBdtunxWZGEgo1QAtl563G3RNAKtv78+mbV
ONPiIM+XFjf/oF9H1jNBrqOQwMzObc0LF3ZvO/JXswaP7SpWe0rAdtmrx9DvLvn24i86hdBkVNZZ
cNd5YaPpYG6gz6/9ds1c7xvCwk+QxPVo0j6WzAXEwhuT8DHd8AuQrIFiWDbWcTjnv7Nx2wDae88c
gipcAksKjiwe5HlQtxQaoRKzbFq5oiIfm75wi/76DBrzXv7Mf5F/KPOrtYcN8xmLYgy+GUt161ev
vwzcPj4yWF8+LnYvj1mRlx/GrIDA0Fb92jk4hkaJ9kVbWQrp2KnjjLT5tcm+TMw/IoUoqqkEPhUc
5MW2Lzgr4yHHut6BOMRHVCxplIjb4PZQ4R2BSBKDvgOIYGLTsG8E3TmCgLVu0xqQJYamARrJ7FPS
ewl9izzwB0PN6JueKjDPw2SccxR0zAZFD41OWlSLYh9SoV07IJX4gMVbgk5B1lReUe1q1wrPIduJ
ciWQC334OI1NDTqTxdpimQD0VVJga+T7yQn/lcKBIp4zTo1iVQQGOwwG3+hHX6bYpN7nYTxETDA9
2S4v/3JV5mJad0grExDddr1BahgMVec+b1zSv1jd2ts34nzJIi8pFAR26Na4n/FMyhSQaeAd0RcO
9SLXmed27kScqXnSr/iMfzBn/PjFzafu8xKv1jYIR1ZlhbpAJ5Dmzt2po9c6qaYdttjPW24fSRle
rK0v5bWwsQl6aZk+R+CdLIFALf6E89YtHWnuiBfJviUB58V8ZO7WoENRBfAc9IQ6XxDS54GZHkmI
GSwqIdHt6pcAs5Z86ugK4a3SmcRTssAcQaE//+Mcet2gNrN+qneczL9GWYAadTwW90jutDqYMe1k
A1zp0rmZpMagiEXuXEn1UX+mqwPg4NcVPdl4xCQoZX0J+W7ENLhWyjDgBpTNiKJ0LrtXcuu1dStn
WcEinu1Gqlt7L2KFgmVoAhpNGdSTZQ3ztzWbN8Thp3tBgkbsZ0jyGKMEl2oa+X26cbZiI22e/KOa
Wr9DWeoqJKGqBa2cKBpSu3gUFpy2VN7FFtVyFpMQ44nbyUkflDKsS/u+ph5/54fWnihGHrypBN/U
blZ8tKZ/sYpEEaHBbbbjQbFDp7iZLLbdHVPD4zs9gtY7CJB4SN2Y7tYU5PcgKvCZDGeSczNjq2aC
0jLCRIkZ/8f26ZNeR2gYbYwIN9wFcQexxlySEkjb7ylunoIdCIbmaSjq2p5nEVsxDepTvfRGDdhl
Pm2x+l9Og99HihVLk4FvzQ6NK76R0+yj8jIQLRhPXkIaFIlK5OmGJLL2kKbFhXB2UzPpNdeRnb8i
k+Z3Gh/bJsMqmEACsZELP8mFIC8ZDn4ECY8SzPQlP2VyXpJCCuFBV/gRsXipLDglW/zL0m2XBtMV
vJULqZGfWVEVg1eorV93cfYnrDA53BBeliwM/tM9Y6jqh+tJJmTIiZwoxK0NqkVBzhcEvfC/zjFM
1xRfelM5NmxW6u/nu66AFV8uUj8/s1Dsmp8+U6nbjaMIXhaxhf6ohNDrXWxeulcr1Hltjev0vune
/5oJZwKEbmO6wOzW7H8DXSD2gQ2zW7mCCaErQBSZFtX8y9ngNpLj1kFh+xL/+kAxG/o5618A4Ctg
VzpsRFkwVFJSb06E/jyGtwdfhw80CGUmzp781/ZJaDeJ37T8QqOiCNyX9llQoIgwmQ03Et9FZTGl
g3c8cGk02UQgBMvewlymo2xCCzQ1Oe+9nUbblcB0T0M7BbOG1BXTicCr6yADwmvf2mPmASQXhoi3
AtocLBCmNzJ5OiKrfR/wXJhgIE+ckwwwcBxywH4s50M2UXl4ofPIoklsc5FNWEKr9cdmEhcn/sBe
X00C0giDT1kZpBCnfnXqyLQDsRoNZDPBTxFwg93BkfEhHZN8rGSF2/zSHaZweRQcdWWN0jFigrKI
HsUe0sj+xeDWnmN+zCuzqrrdloB/smDJ4si6ZJ4Cr13v2JuO1lO6Ddj6mLBxiB7Ca5w25besH4/o
u5ntk3r6l+NFwix8dNm5h1TDzGnQd23szfwHeWm33TM36xiz4/FjNb3Bp7nKWUkdkaSAUpppVtmV
pNw3+EwWGrIarum3r8oQfMBvH8vuvuBJz2p4DfE81fxgA9pH+jSmOWe76/K2d1mCI2IPZDMxQKTv
wOejtEgzjNmhEGk5LhHcEXfb+PGEPTtMClx4U89Qht6ybASgMMb9amWLOb/5GlztCebaXjrwjsA7
Is4GL1jK6xqdxvMBMdmSPzho84Cg/24J5+H8WOsBloAhJPGDP7tVBhowsy+L7mO6NjAgq+41JJGZ
dwqNQSf6hWtXMCW1gt1BuAqy+8DKxJA6mYdbBrmnRcvrTVJTES0rDmKRL3Y/q6iOkq50n9K02ML3
8+DnJf/m4lyzLrg5cSt/Lo9zS1QxAxIxwyb8iLfjCRtUXVDcB9dKkk51fytk1x7L2s7Ed0R6mHce
Js5X3z8UwqBGB/6gFAQcsDee3B4f+KgLcxausH4SzyovYTtr6aX0fEq1M1Ly4TLgou6eb+iR9hxP
p3N1mahzFpibm6lC+gme3+jnJJ9ShS5s0lRVN/27YZfZyzQ7mSzeMYxZnhbkUOLdvWRh25Re+EA+
jx2COSPybwc2C5hr4A0YJYZ0l0kCo5sfWJBQc45vonOP0ffJrcgnr3hTT0ELNSl9Y6OrXfdvSVsG
uEzH4qoPz1XUTnK8ZmNV9y4MUxfgN+YRUQLXR6TznvW8L6Yh7fQYyr34XCyGp+inPnO8CtE26yrR
Du0zWCFnTod8DRHrGs5fWzGpnHoyDOhJckpxl2HsN5DQbjFw+XTeHT3/TaxvjGqMMLL6q86ELywX
Wyn+Q6Jn5MAhKtXyeNzStFBEjuheLXLJRHdG+e6NBc9rUp1KjIrj/S+pKfQZ/GaKsQopoqsddc6z
QxZ1cNLiTwA4Z75U0VqQj47B8/LZ/UEJP4ekdvGxbN+ITECe2gFw7oYTFWLCPunkzAZtcLTBphUE
mayx4KFOEoJsUaljTTwk8wbS2rDgOPOyU+eGdiMfgaYHJQ9/kE1w40N3DZG5tsMy1B8BLVZ31xLz
XXSwJhfrO6v3xRuQLaCm84GGPp7HUNfzHW9f3l7B6RZqJ2M5mQdbkgsu3DvbVDpU73B7yguZ+EQa
bBhldEA3bLXIvfY+zhclBcyaIXENur5okZ7biLaINbGOM7gBB4l+/HdK+AsOe9WELNrkuj8PDX1K
Wr7/xa/MZmB2D5SIoocgP4Kn9vTdnfqfaGNmMogA2Rbd17dCZSPJNpECaLOOlZOFlk+/NZel+Gb/
ozesVW02wn2jhLWRaHpnCcL6FsiUKKaEE7hHGeiQqEAYRM9hpgOgU51SbjbzYNR/V6weVDFR8Sge
8Oek0XhtIGsvUUJzuKduzG29CdnA4t4IksYc1Gk01w9pCRg0OxYgykHxxWP3F4/iCpoDCA0o02r9
0DL1FtKRjfTTRCqV36XoZ8bkitjsjATDVrWfaq+ftQBs+WtCAgi3TXl+2UnBicDs0l1AM5FaWjOe
0jrgpfbCd9Lbk+mmMS2hviNwEzCpRVMkEH6PRmUhryqRj3wrQDgv7+SB6vMSmDWvJmpxnsvTcIgE
2Ow/81bL+6B00ZvnyjOGuIpBOcMERUZms6QwFpHL+aosj9nXULabPLS3MnozZ2QEnaw8pTT7DHFd
WwMpmfAPvrzOn76AsvVBKHhIWFRDMQpBhubnwnfKzFNF3hhOYrmML+a3lyDaltNpGtl1xYzfleOI
oQ6Rk9BP64g/sI/Q2+1DvJ/wWWH+PXfRbWXf7Pz9dYj7qyAlIfR1WDswtLtNMIqKHqMlFOOmFc5d
KCPM9LF/WhJD36D60xtpi3Vo6JS9DhmwrpFdzzaw8FxAzkZtdvj+pmWmr3SxPp6LC8wjLPPrqVR/
g1eg6td6+9u3KueDL+nLGpE1/tfVVZw+OOISGD0Qmhe58YJaDZPPzNCyCzUd+PThATammnYL5+xp
wRZO0aX8BEbOdDlk8ddrsJzEJWtawLU+1TDsJTqc7/8haeEiwD7MHFhUP9AGkGyfTM2X4KU9F2v4
VsUYdEteVaOX1gmyN8tipixDF45SmDAhbPeiVYlhNt8umU54bSDZJXuJMZ67hMIcNEJWmm7otgUJ
3NIsFyeETgeWqmt6m5nts+eKOsaM+XioL11ry1XJMIHsg37/jC0rFblFOUrXEtjmjy/ODlgCI7B8
m9Wzo74Vtt/PfFZ1lMlgok3DcuJ76Y9/uh93pyAOqwlmKObX6urhikJ0I5AhfE2kVjmIIhoGntx3
o+beget3wBHKUcckdh28HxXzC6CZVxkT6aEeJ+Xw4UXfqTSB7K1svGu0TK/QItuSvqtNYFIl8HNR
slukt33gCSRplrTzQXpwABQCuW9zj7kSBgBjycj9SDqKiFi1qODAvAkln8LgdgkwgbmskAj0M9UG
sb0GMwktkR3uDGsIxH4alqaZKe5+GA0KbRRP0jWbYtYVbL+vT23am9JH/DHxtfcJVdvQcIKDfLws
ABx+DL+Du0QHhNy6ycSmIEg83jZnyD8qJpi00SfJK5wZ47J2labo3gR/uZ3H8R+sKgrw3VDDTyUq
ITZAbuS4ZUhcHmeZPm2zb5O5l5KvsXhYsgmFmoU5oxPd1nVVB3T1IaXVkrlTJXPU+cmUq92EJa1F
I5JOntV7rtk7hHsNN0BBvV1przN7IZJMeouC5eY6gvnDz7/6bHplpq5yhXz7Rky1IhQsP4zfTBIk
vHkBxWz8Wtoi01MWqCbAxdS2eOmPBgzzfaDOxEmHEmxKk5cJo+EpSyAVVafXBjwC2btNCCgtPC+d
x1vLlEJF2wULKkPodjEbiMG1p/x4uTJ7PqoHTaj/5aNYhuAgEq6wXLp0ta5maFYpj6gGTa3Yg0YD
YiYHVsiLfPOK7wOPApCcRjaCvWTJeQLw0v9JwBZJ50NKKGduWNAag03pRaciSfemPJ8wMBfOM94w
4V4eZimXWhsSKB4xgU1vNxOmsBdbWk6H5KcSoomTGyh/NsbZ/EjJfFGqr2dKxy+d6B11QLWVdWlh
akGDdaIbBECdkQjg4iSiJCdmRCQQphfLuWNH8YpDZT/pRF6sNcRIzfS7+EjnJNYaD3oOJlR0kO4e
K9Q7DOtp1qF/22hOfcacJVoBcjmN/PaxoQfPAJGPD43ItOVQVKpmuUKp+VCf5u73NIXdoVnX0GGd
RJnKe2exkgII6iMuU1eIkyImQ6YBNmg/cMdGjsfvmvSTthq+Z37IMmwxV/bcO/ymh7qoLbMBBbis
V6tK9CBWlkEK+wlTaX33/pL8xNzNRwAh4wLq9HM9mFxa1jujPUlSDrQOeesa7CX1PjV1r4sBkalB
/aX92FFi186i3YKdMct8Rai2UQCzq+95M4arHExkE3bGATHOOGy9vzRkEQIvgt77mhC2MViyxeus
Zn6w6tx7s8PQ1SQTPWtnmxNwfHa2ab9WC7/VsSJbKYIo+4IgJ6XS+Q5ZvwDB8DcLAcG+B2B9qGGV
RJBzPOFp/v7SXJj+uyz/46kqeGOt6gAp56+XPibRvTEjehHDH2k3YD9Tx1jqmbl6JQX6ogoYmhZr
o/TXe9JZH3xrvYc5n7S7dZ49E0hZMBOsSb2y5dkSbmHt9eZ8AaoPLCAgRU3rM6ucRmn4HqUIJTYc
Ycz/QxTyt1QKV1m4AfuqExQlxbIt5bLJjulfh1Nt9gm2GY1CpAC3Gzu3m0hRBTMNpGeiTn9hvS24
RojShiH9W33DGB2quvo6BPqio9j0cfOwZWl5xXLLx5WdqrY8TEHvk0yJZnmMBz0CJ6xVe+R0DgrB
01z+MHdzx4YYzfZkjeUXwA1YieT9t3HfBSa6dnUZyE94kvKTgBJhjgYYW692UYufte+V6EZrowS7
WAdxJ7rhgVGJwg3o7sVGaqOYKbRNiRg5q8g09uB0SBWgkSBQqXLHh8kUlNzww4YMjdjn1u5Omehq
fwZuEV8nznBY6qa0+AHCb5PcTU7OPO+cGk7qXSiK5Pftw0AG/rBtvVDiN3dMwmGbyiscrhk7lUBm
UZ4fMFSKFVTHicSeFvdwKUDjU40TRuM1FaU42ZHeOP3ex2DQZ6M+TwbbR881e2xfQGeCkN0bWOgY
9D4Ss0xAiDnLUDLIBC+t5na3bPjXAFnW4Fu+ubWBNLaovoQPypWKiyVVfryJaBpqdy3uP9L9RQ9R
B3LnMRNP+QQLXWf6ioIP9V/cbi46NxFgoVTN8Z2dJEcMm0cn55hszReNEUNiLuh9g1sfUo876Ls/
oOQpY7bcYHwXpFKa1I1ObscadrOA67w3xLP9Vn3OwcQerO72XaZ24W1QbTj9FK7QnWxH9GrynQiM
Tvfv1eH7Tk57bHlOcU+2ejN/qTodv8rUCQPA3SrGLjbcBtymskxDL7ZYz/0ERmshdlDBCvC1+JwQ
NCinuCLMrL57nP33xERX4HSOEZL+oBJKbd7Dwi1xCzdyV3tX9nr4wkRmHb7JhF+EC5Dej1A0isBM
TPmQgv7+yosGPoWPRbsatQALOIteXo1cqbh6lC2lgny3O7Oqlpv8xcHuIG3MH5BvX1c5lfpXEBad
1ir4MPO9PntfJOizNY1O1Iu2FTQTg+pFleRzQOyAuwJXRQYqFHwvtWWApOHpCfeqd9Km8Snfh3Lk
XPtQ+Q8Dg8wUMaPXOcSDZmepZfwXhxaMbs5sSS9zor9wwExi3YnXSJMOgKli5JpYkPfiJwYq1ic8
eIor14YPBA7WrF8oOpqj8vCDwVGIka3sLqAMO2FaHWwolq0QeCTgz7VWvIiJws3Enmde2WHA7OnA
cNJqYxKdK/RpRWbeusUawl8w/M3J1344QDiGG56vbb9K5Jcbzzi6L0UHtK4x0ZUpbStbz0Rsgy7s
D9AcPandrlZ5puioft4XIO8P64LuwvddJ2Nc9ijhMO+0yi4X+ZRcfiRLyH/2dhSXHrYg3Q4pqCv7
dmR5IX5PjQ+maVO1+jDzGtobDZ/K4TiewJh13GMoBIFJZ3TUuoGrcfj6Cy8r06UueDgPmajkTCs0
IHZ3kmo68aE95dC+Ymxm2BhbdDCxq8FBFFY9D01wuZIfRuW4WripxbJ4hDtAZPkw4ZcGCAUGiZTr
XZgaJpOvUyQ78NYy4oAs95dh3tdRttsUnUOe8RNmgf1t/PYhkpxsiKF7P8iv0UAbj7yZGsLgIr+d
WjvxmYmkLpzKDtmyaFo/MC3QWGxAVjDvIgEvc+r0bEzXPhPsRmTI6xfd2ixjC+K8HRnclMF1MIIE
HpGDGDJTss9W9kHQygWpulV0Q/582TlwEF3psCixB7dBjiMJEMHn9MgLayfGDFy2VUZKkQHo5C0s
SJe8LMk1qVtI+EB1CaqoVtaU6yZofAmeCKfibHMcWdm9aySKGklR6gGtvh0FQICSm+AO5/7mKB8u
/sYSc8MNd8rNQJPvrsL0drZ7DwzqjLTvy5mj2KsaukTHlzxX5s30SidaY4dKXPkPwQcwEE2Kyfwl
zN18mxHOSLpJ4qijz8VU400BCQjpFZeIzOPpvhFCTiLI0VYrMvoWwyCg7el1ScMeBdcz7SlBZGGU
RxNWhagCazxxqPX+XL0SF1PG1ukZl/MquUEiZBv70eYvSgVtyrj0jg0bwOdwMt3Psv8fP9bWf+r5
S6bixfgL73FrT5y8Ghu/bwWiSFvezwh+uccEnDhzSzjKbW/n0Di1IV0GMlJHF+jZ7V4ERTkO/M2B
42ncxisCv3OPwBXsNH3m802ATIviAGLQbV5jhb+OWNcIa/dmV9rMYuNLpI//em2L26j5xeYd2qQX
UF5n9vghrLHIhGxgdV/EfA3GoXYHWa+gYD+WtvG/f67FRANpWoUa46I9zIFbx2Cqmd9fzgwSCUKU
gm4fs9Qwr7ZeR0v6yE5k4Ht8Hy3i1Q9C2hrTrlStnA1AwLge1LkDMaMGqVicfx/7wnGciq2I/K4t
b8ZFGDDTN9S1CnOTy5dNTxXoj4xYd0fieazVUlgYDYOl7HRlywkvd/VxA4wL8gHRfb5FsMGIA1Kh
+hZ6ugAcLd4h/st4EMGMLDCO3lh1NMGvTMzDnqThwLRK+j/PLWNZMI0KupnbnVvj4lyyDzUzuSVm
6zeozzULtYRvfhMBU87OrG32zrOPl6u0vLTL75m7pomfmQPttN63yPgpYyhm1pKjRGFK0FVM28la
fa7gS7RSfZ4QAMAxyk50IGFOO7nOxDYY5t44zEscV9Le3owucX1JD7M8a7qPWfWA+szHFizd+OVg
Z/PbgUT8Xno5AyklIA+Ohz4vHbBehPNLo99JTj5WmfXAH+WADUYSKerot7Zmu3F+FqE+hffeJUCE
bhjRQG+0cmIhyjVZV/0VJXJ6yllinN6QH65JvlZLbGnGMl6pIFNGJY7sVFfagd5uEGmlCgK6sbvB
IvGFJvZmb3Z5vj7WPcLnGggj30QeAPy+eRbtOS75RvoIuUlhbUwatZWNtU3CEzKDhyN2sgbjU6z3
cn1/ehTzgr4xBrZrDJqiAD9C+9cgc7dmF0/jLgiFhhNMf45Dg/X95QFH8kBISWs2MBkTc7dPBp/E
1IzFXODUvOTiiTo45YveQ5AEOCrFKvMcTjakxDDnt+lsPAIVD3vFSsnGB98mPlxmw2inrlsjQjDl
OsEmkkO/KMrTpFmWWiln3wsVAuLB+rWq12h5dt8I0XdUv7LjGRsVyhI7e4RtIaFo3oy1u44Enije
96HNTrIAhlAy+KHXit8zsHgwyR7X5sEbouGl42ZQJl5vYfEE5U/d0iRK/x06UknoD5Gi6k1piWtP
hiLI5Tv05DhFRAS71Bk09cZy0Gk3KaEfDAwlKnQjtpUJo8gaJZiz9mu2yYBB4Z4X4cugd4uA3aP6
ZTMh+HwLlFQczc+2oizKvoPN3iXwjKWWAVsMkSExXQXlld1APfS4ZVcXBAXsrK5EKX3/yPpYtPzw
svy1DA+qKr6QnNQ7OiCa7X9UL9A4mDxF1JKbdeVdzWv5B5SWZZUPtmwGfIdQddk3fJEbLj2WU8eQ
cQT7uD2sJrtvmiNv7DeARVo+Z3gRgNMnyEwsmxfm5Wf9NsdCDLEyvpUYii71BmyVS5cBi6zJ7cMI
1ztP0HhTnpJlklkFtrTOvjhwEHSkd+dWiXuHzB8xj6E9hvY8YB9zsRk6q7gAUGXrDFTitS/6nO1d
8xfpIytFOOILQzF0aIcTpaPja3tV9XIlEqsyWfs/H1Sv1z5mzPFDn6AYyAI7B93/MuRAicz4VZBA
yr9UpKe0k1YrCSGXdT566n7UoQaXJJk0ytDE0RL0tciceQqFbKHKAUIe1KgHOiIMzZweNdJl9KSN
ljFDNTlvFaZSC7kBD6ycxXxj2v9PdbYZVfVLZh+MICo79I79+h38aSCQRw+eH+3xexIflp6ktwRg
7taXXsZbmIfd+hIapS0heWIMvdxpk5FGaLBxtUeQ/VXCTYmn+nBTlhhKG3+L+oLeQSNfAiy1xA62
J2gO+V2Auogkh77yHKJvylnxvTih706HKCyuzGZzv29K3Di7/3aCEcFedwA9s2RdepLqKm7FAKy0
Jdg74UPMXmobpPP7ZLlvn/UOjpW5fI/dctIrhzmeLpLutZAc+WCdYhliWTYMHEzC51ES5wpu1677
vGwBA94EJ5An+R9fm7mLf0TcAZxB/21bQTwXJyvkKeVmZ8k/HZTfCbO16seD1fxM34zXainq2A/R
SM7fEYDujYCSj8bwwYU4PD/MQR/XSsPPZcTPetRkiWc/lZOKygsR7L6x2v62xrOVt8inBM4U/FiI
NldMWzVskoFRNX3/vsde5z6DmEmgV8KXSlmbUk9oIvOIHeWbX4ThkzNQ6W+jdWHkdjqqeTAmhzbG
qC8/ocNtNjoRsrdH0UEVsjLY6dGyu4ItcU+j2Uc27YzXG3DMfJxqcrAvJFPN0NBMV3nNu9wVZ9d0
jkYy7R9YNPNyhJ7MhaojL4nuX1WPm/seK0h8g9L1UcNZ1d2WciMLO0BUp5uFxa4jL+SKH9wPx7NG
hlggWcNjoHs48YkPA6cLlYSmo1KAho0UO3d7dW17g6ZWQjf4mS9WuXZITMk5EM9ciy2mC4raX6sf
sZk/C9zBJmmQ2y5nFw10FJkUQi1TTXVjKnrMWgFdSBQVnaZ23s8b2y+I+H5lB+2En0rY0g30t8wg
AZPdSfVjtDsp8Nid0b62ZRbMsFcAtUheT/N1pDTLoSTu8ULDgNrxuQDVrJUtgq5FBImhcP1ukEhZ
AcVuLZvAs3Bta1iTOfWNMUUxWez0bKNyHMylfwqHqM4DIF6RdBqK/drjd4CyKdVWCm2VpmL6gVWP
p96P55bAy6B9Fateks1DrRAJhMxk7hn46ifU6xNjV7K3qibhDV4nQAOHIIe+eVnmtUmp41JPJJrA
/QFUxBL5ju9+NT5YrpZZAT47gTVIWerm9CCLLUXv4JtueiyUSRBUgW56HSH1xqqD6Y6R59kW5x4U
bjtLtJ/5dPx0Olsko1P/iXPibpiNUFXxzx7+LSkGu2MSmfedMyzs+UbCNRMxTwYFunOeH9ogt3/x
TE5NaLhwbkfws0ALP5IASapIRNfKKxPJDPrRr+WiIcBWvHQKjdvqg9s0kvwc9PSEV4425Encwk8D
vTUHcyy7LROojotkiW5KejQfU1TxQts2VNVWQEGkMANmgJjZ8dEId0qc4N56L88Cxo1HwrPxsG7W
36JPcVcNuiOnSsaTx3aFB3uHmtx7YdMUPZf6UGTG48ahvPAeNaygQknDglyu5CYQGYpHaIspJLTr
89mKDvJodCXPszZ/3DNueLzPy425JvxOkS2tI2JaReEYq6nS8Pb9urqvTWjzgIpv16bNrQDU0lv1
QcJBok9Q4/GLuSTWVYIKbAdDhwtL0oRj6oEitOl249vOQ+BRaLjy3nBqvhtVrXkC5oKel168GIM6
w+q8JBloPHbLtkb2Zop8848eOfKpKoWKIVc49QY+d6pyJUiH5iZ+Q1jLN14iCGGepP3V1Ok843yL
xsRywPg5UisA8fHo08FIYhoi7R3Y60EU+m6bQMG15DQrC0oCNQ1oaS14VZBM24MfndtLCKfYtrET
+R4XJBKRf5CA2xmpI3pfQiB99hOHGZOebrhnTDdDu4B6G6YJbfbzGTSrEPl4MloingBgte+vstEU
H8XHUd29fIiH5Gv39+XikpdAc+a8FJ6n1NHzhEDIeC++5nS7TAyf3ObcxQkUsHrhj9GSCAcpiJfz
pQy4rMqy1RiqcR8c6qLucp8VTIP0M+/54tjhMLrKYfiQu4nFio9xXMzDpfs10dNxELAEydIdw760
YUlq1Izi50DZZtnBnNRxIoXpBvU6R7FCBEu978mWSXtJOXRvjRnMlhuFUx4MNuOBRM5LZaxaHEfF
klzMU3n1OwB2+jIq4cFzPurK4r5Uy5DtCwOM5czQ7wap7qWIbum04r8etVC7GzXvT8NkHLaqpSKr
AllSQqvABV6Ips2ieUeBnDozkKPkGzhkFD4+3umq6sTut12dGBo3pDEvdLbKmZMqxjaM0754ChJ9
EqTJ5/vFD17T524g+ImEJkEwCfQhbE7x0pw/nS8ytZxHrXZJqHH+/hcjTnyTWaNCsd28Q5THa6F2
g7HIkmHBoN37PypcHNx8AAGMOfWS2HSYZMHMKBXwz8EtJrcbDalwE5PWDSBQS4mVK8A4UW5J1bfm
dku3XuUO9NF5asILyq4rzcZZt4r9mEldfS2YFa5U6E4uBqo0m3TM9DAD+TXCLnVduwRH3zN422Gq
XR/mzzXF5XRTdnunCSbitNoyk+h8GoRhOxb9MAtZpYJ4g9jzbeX/QLsuCvBQSc5shxjOEQGTCL7G
525Ii9N8GJCo2GwhgMTWycZwHTmERVdjlZQkYu7SWSCSgAkMZ16zYGIyKVMjK3OMHEP3xd3KYrrW
WFY2ZUP+wMBEJmUakIf38K1P4BWFV/sx6LYITLIc3shNtetzNb2E91FZ1tUrSRRCMUBAfx1MA4PB
Fc9fR5jaZpXu8LfmKgSD6VQHJUldzlSLQDR8T2zeaprOfUBdqksQhf7LAp6APPnnUDcxdJsBI+l9
56iXX8LKW9xSJtOBj6FYasaXmx83mO/z3tgyDjCJgZRpchiHC6oXgE3bRTn6tgWgdaujLy8e+NoC
LDCf5dWWTyaTA1cuJPfbwf93YfMQwaYWxCQLB/E7e1+cSNIv/8oFBlmFaxgnEgoOIlblohaXOUQq
Ro/SAltGQUlwulaaIQuau60vNzPPx3OGblG8nA7gNiTzzNoy3hpjA5Q4kNztty+VmA8VeKpqFHmh
GRRoKw5yoVN7l01uOWWgAYcbnTwawjgxhc+RuhxyL+5nbu0SQ0tNuC5WuLkHNqKv+WoQ8b/nEM7Z
LoABKDgHu4TXwjfkNOx5tb+lX5WpdEWICVcWLdY7byy7BbH5btc/kOnVwYu7ECZpegRlC1tSvwbU
3h1A3waoMMh5L2G0sUmULtEZXto9qnvKAgh1yfPjHTLsKde/POwaDT0AK39HkcbJWWV1PbZywn74
TX3WVggxG2LEdLyix+OOHoI7NWAx52W+g7N/4tFJm0opYrwbj5n2XEVbUb/h9O+i/ggM1e1PbWzD
SLxSbh40Banc7/B8Qq4IYQmANWdyjVHr9bLoV4CNVPnTG4B/Vm/gsyE9pGw6L0FsxNqHjCZ+vU3n
8gYyb6Ulr+FnUXaSjvpd8WClBs8BrjubWNsIy7sqhtHLs1tCe7Kb87S45zwXXfzTA/VrA/8+kgJC
w7UXHan1Wc/zPMBFk2t/ECngDJL0nOe/Blfl6LhzYHP4Duw1Oj8Rl1r7fAIbGn1lofXkHiIcX7pW
kWqgLPhISDGj6PSUHR8lZYP7DBhQw6wFKMmfh6Tx23Nzo1iaKAqUAygPSwKPNLKP4jcsKtQ+wPHQ
VDjApvW8JoWskvbXGPEKsOTzPLglfHgvqL+2W00KXX37Hat0hXH2ZRM+8dUSxnGpBwm2pCvcbwTq
9cI4icKznX/C7oHidik2gAFMnxeGcGSeNo3xsppXfuFekesH7sAw/lfqQJn/ErxVb2NJMFoS2oS2
FMEcvYtJw9Hmst1g+E3II50viRq6hyU48fPIgfFA5qutcTQmR2UQ74lRrSuj5KW9vprlA98V+zwc
f9pj1UWPo+CQ8NQLOdwj/NMRuwQ6ca+JbjbeLif11G4G3dtA3Nx/x99a9kRkK4vJh3snE6iDwo5n
D8EWzmzGEZEVCNj0VQwMlbpwok5gfgyHT/fbrImFXOw5jpRDtL0iLQQVHWe9SfOp+sC5TBiELO2V
TtiE2ofA2POLOY/Z5y8oNDbD9AuoZrU6gxCxQrsANA/ZSj5hIIfthM9BwiqceaM0BOnivEiD1Dlu
e2TdsqzqQDAA6pBB5iUlKGbgqXiwpH42TbF3qkXgSz6SZnHy7sgSw3t1AJ9HjSpcobdJ/m8ndzIT
/5zd4zxlG8x8aTXWiE3pJaPfxOwhTg+QYNSVe+rPd8Scixm9mYWrrDxaC4aE7LikZOvFzf+Gurxp
ARBRg9uG/S2bm061O8VwCvJsustGmBlNKRWXPQYW2Orwr99QWcnm0FPoTXUdtgyWKbSUlkEb4BvA
tBupJiPu7TWhe9ziPfB8qxzEwVxBOfQpu5eMKNjfe7Fhj5eakYrvNBIn2L51kZGuCpb6AARmumGf
C9+YVrluFMXhtStXJBDU/vgy3l/xT8cU0Hxta3/0CziCZVmCNHvIOYQ1xJ2dbfU/lzE7sWj4Thu5
Rqv5K4+NWUN39v7Z6Ah/2u3sF8whb4VRdNeuoFdxStwsbOMNsUrnsP5kYGhuvqzEUaWdB3uZR0kz
n7Fi5OQLiVdIicY/WSqAgQrC9J6p5cr2DPmgi8kNAZCYlpDnhIuyEN1+CuLc3esDQPsf16qjT3US
5YYsl1UN31XvIRqncBtITH0GfvkjZ8TmoA+lO3OIED+7XfuY3Rn48OQWL+8tlXQ0s+3FCvNUro9Q
SsWmPc/bgoNsL07NShoeKSEZa0dAuh3N168rSshqqd60pfvO7BY5rKq3qpbHT2vgJazjJ9wfby9z
/kpxRX6RsXo8bFOG74qkTRkVpMzLrrSny1MfUZHTROXUSHZi7ukj4gh4/E/483Qr58FleS4h5jDV
6kaMK7zupAqFfsC76ygp0h5H/F8WJXULWOfENM40To10KEp0pybtpJ8jmbl38KWOXBykx5mXupWs
BwZJo2c6KN5G68E4UVqJHWPKSSfjqtvhS7aMgM+XMB9Z/CPI72zgAccVWMmhcWcvJc+UkMVIwkOZ
xP+MJ2lUnh9vTvK6f8N768aj00kTbCFfylr3Yx+j47pWH0QzAL8kMVEL8XzS1AONX9m6/u8o5c6d
lp8XmyoHX/o456arREob8M5mOplCbSf0v5n91n8FsfFaBqRlgdRl5qSnBgdkefpfS0yRmzXcuzsd
rQts6hNtj22IJhDb0a4H/Ah2JqT7zEIO+POgnrCx/y6EtaD8ITbjrq87lUWdF3YZdCVSQIqI1Fjx
ORpoSD5Gw5kefCdwiJho6yqAjEXO9RrWkjIYvTmJ4a/zwG62fBBHA/NMNSpuSh+2Mc83UWq0HVbt
dPCPQsmmpuUF/3rrUqMWOgoV781QkOl+cb/K9yno2L8a04wfnO8iTaNWsqCAp3V3/naw/dK7PFwE
DkoG5nhJUkfPn3LLFvaqBz0IeLsrb0xu16t3uTf0f07ZMwqpstyW0eTc0pbZTb1HDeJZ+UANZ6zY
BwSWxlf/tvS8YuyLCa1qfRJyLYH0ujr7wIlNbSP9dhWdH82Z1g2WR57FF3wzWTKr37Z+8SBaQOuY
/o2ENjd6XIPi2D88FrYH0PkATfJrajJV7mqaWdjV6r7SGKIoDriQlsnuHdTuF7POqrnor4yYcH6J
SR6JZ/CTz8BBJKdVxCMurNSl+VWJvtIUkD831tkkZ2K1vKPuh3YtDMUnwWhqZ28sz4mddfxvZBET
KMHrXz/qe3qiq3V7fnKdRKFT6sesBiEzx53sgLWc7Dr1jwplGsb8wtkmQ91f1jDpjOlvJDCcGaUb
PFHNd9PLg0B9c1vWLM/wP47QSDcVEagYksy9OjqmNbIyaek5uw/COBKCBjSi/XDhPUKwXBzxpQf3
z7IP7Wm+7C+UcqpHf9XkyVu622O0RbV1iss9eMFQsPMfiaY1PEiKACg4evBgX4sQugwuTvbXipAB
Lvtkqp41ZzKZNBuIikGHOSZjaUUTdBsQw7t112cb6MSKF5Ydnh8NNI6ag3bnh5iq8mAvReoGdDwd
olO5ULj56DNc2iAxLImOD8t0iMkqP/2JGxhCXQhn0lxy7loVEw+r1tJq/a9JEp2CV0jGTfmKEcmp
aOFvkDhJC2hlAHO88bhpECMnvyQeUmqn03MDvIlqpy+zpDdC1WH9dCJkW4iS4KnA5ogwUii3NdBe
cIsa+YrG30QDcJYA27uxbwbr3CRb5YMRxJfm4GxowHIoo5Fp40xAgMXgzTEVgFqiyKXn2xcNeK8Y
1W9DMlFC6R4vhnYW9KAvdbObJO557FVpuzdg+WzGE5NA9U+o0+y9PdmFU3WCKdP9/DSfYJ0EPiwV
2TxBDEjfJwxZ2zJZxT6BLsVg+BT/M/H7HJg/8y6Zd4ppChm6pQCZGY9SQ4Z+25QDScQoNikANnW7
iDvy3ETqicmP2ZdgYCxzJgmBknFa9UlVfXvDJpqBSgOL3b1RlBTrdBHNSyGndOrKvGgZJIGbWX52
9Q8ZKjYjDJS8C0qq+DfiQBbcq0ITfj9ZIEv9yTjNzKPBai358Ci5HRh1RA+dYSwfCdxNWxwZ30Xn
5lfN7yH2mjk1jXcSLEpD1/ddAQfzrRfx5VIGSsp0sTn3t3KK1VMDpRSzpB7VyaG2CtYrlJgkdclB
LyCgRNerfZoTSmo+N0LKjCzVemX1PJ9+w+Zzqb8XbVnhfx9b3jFlXgv9sx064wxKTv9h8xYp7r4b
vWbItr1bUKawuXTM65ULO3EN/Ho+imUqXV4S91xyJMsFelRajTU8eD1MQBV9icEg3N4fmRi9eZHR
M/CJMGM/+7kxuP2Ht6v3tNd3nFbbL8A69lMfDBfDN8PduabUp0kZoq7EYexSWEmr6ivgzEAXmYD+
FvVmoHNYtLhtJDFtqHRtHs0auZeIfXYYXJ4Z9xq9k4QqfSYDeZDzFgnhB4rfIRVMpMA3yRGEEcfU
3saE0hp83ztWhGyaJz8maOzQoHAQHXmM0obOc7Lcb5ZxQJWw5v2w2cHAf2jxjC+StMXbwVfsOMEf
+wZSZA8HJACuDXHD6cUCxFcEbD+wsOfoHVUN9+iMuDcz2NQfCvvCVjpP18FLvO0u6ombiVSQndiV
lm+o2qjhj2zV9JjqiDn2pe2oT3XM7ytmUlPU4IGCoTHNRyLQnpOaqpcBkrtAGi2iQf8n6Phvlmg9
n+VLXc0J13ceNpLrIrV2SUQpeg0MIMn8GYf8TQZ497yHWfmjdQRjHz6mDJjjRMVaAMnW9Z/QMpUg
pmRg1UMXacnz/8Lr1KVOio7OxM3CcgKCcnyXtDAetu8tqa/MuMp/lIBhkjEPac2+XJVvabvManP4
uUpR88kJNjXfa0Uq73knF+RWz1RbJ4l/RTMrvMNxIJS9CLGjevW32kNfwNGFlzTxW8ZPFLOijQRx
vDaZvYqTnrbkkee+ws96jJTmQPDP8ImtEgcILvLfc47EDtS96sNAf33ki2HPQEKIMO5O4Z/z/ORF
k4BtebKNxD52CqlkC38kNxm/Vkospk1rlCjOK1KoDM8pq0nUgdWovAnu5BjjjBigUVl7usBugAVz
Gzk0Nas3Y4vYBHhXKsnf5jpEa+brRLV71QvLIUo7GpINFiChaR5Q2T211X8444+0Mz12HXfCJJVX
0Y/IK7AQe31SMsG75BrFZcyGE0txNs/Qs+2tVbU+26uTC7zqKzWG/a/4JDSpCZpvebG0if6DvqXE
dBRdRNWmgL+Ibqs9Dk5KoTj5XNtSjtxK39OtYGs+jpZbT9SQq2g+/wVJrRWADw9Y3ksR7Wmc44kb
FyBaYSd0BeckTFo8Ea39EkUvdgb4ONGOtT1lpTftFroqktAy+uLUuxpezEhZnfXfIM9Segca6K5j
n0fM6Xe01Wn+ZDw5PbwfjyTUhWn3xpCZbpttyN99z+iqoL1e0CIhdgqcHSPbiM+lsSKyn4r6Ot3i
YR6d3HtQaO1bGzNp1jzaoa9P2HIsR1doBwTcoqlTPzIHpJG2RmkWLpzS5Bbensp5DL1cGkrsGdya
hI4gpzZ7JcWwXxhvRaooInG1KCFgSkhqRyhu8uNC2f/pbhZ4T3hA8vWz+7FGNuPi+iuXgC9vj02O
PVISytPGcKo+XT031jsSXo4WYCu2AQVYHbCpON7Ke6Y3OwYd1Qyn47bVHF1WRzyZ8KvFs2YTsGkx
lVHR8bjrxDRgGPVihl+AvZ4ko2XlisnXdnM2XyCCeJDBoh4gpz7DtxwVoU6tc4T3DXLXbK35xTje
3Ceo9+Bx4g7O3MLqcMjhiacuuzYYoKEeWyYTJmBViLTnqI/vxVB+NR9ESqbzS6yggAuQxhKZGEgl
VswVXY34VralkRrC7AfLPACWuqRQ6mosDyVyXmc2T8I+BR7bq8hzqzr8Jm+QOqkstKDozWhiIP+l
lZ7N2t8oUCjNpDJBJW9vTo0uA1zp6X5Txaa4mXlWAZ2kOTKSo63kPDyU/dTHEMEPZ01cYGZOlWMi
b0a0jH518DeRLnqiyu/3w15rmTUmMsnzCt2dsBlo0uov082n73IGjdCYONTuCXPY+lF+p9FANzut
4XlhB6slrNrUf/TZGo+lrvvRgiPe83t19t4g5tk2xV++UNyIM/OAhe4eWQg+7vb+eLYSmpn7aAyv
y2ZYY23defz+L8FLvH3L+QPl6t5r++ka1P6n5J1jqfMBhQsL1SqdKBZhaoWoUD+LuyrRnx3gjf+I
rh9LXOoDOVNuA2zxslOOyGVL7udatiCGJvEcFg2zX7+PRAp1JzRc8rLW/wrKjWQG1Q69qctcmAUf
rOjw6lFKosIHoz0ca5sRgflxiekZ4v5HZNYOfBDLsSjMLg88apUDf8G1s6zyD/FO/hMTeMI2yI9J
Y3OdMWiWSLK0hkDjqmCccK1hw41+VDnvqYDh2gaPnIA2cNyOeWXz5BtPKf8a3g8MZTz0/nEHQXTc
odHnQSkdFgHjE7MP85g6y58ZF3BzFGKengznGYoywJJRXb5ejH993AcqBm+UU474R6shC1ZiFTzJ
H5omFprDmJfVMT2ac5syQS33+F0GcBQLYznJSpfzNSyc3LDXgamITCr4jddPja8/LvtlyZMVzCsx
bhHjbq7c7MRYD+nYb+EKi7hNm89CFziiGl3LhL05uIHmGGWcaqwzMqXYZ9RJsTsqAXI2gvd80yuf
G60QdvG8+IAHC1Z//Bqidjzg5/bsN4neGw7mDalDsxBf8nFYXjPrqiRdfAp0vo2IlTn9ahcpIReh
0Abbh3PAL1IV+LR9nk8b2ZSJjPVWbxtju+Ir+gFedjJxJ5FC2LXJtnwjU0BiLpkXxw9P/tSjcN6i
UZljr3bEJdUXZVXPu6iIshKVJSGXGS94yLROOwhPTId7LxeslMRO++6dPXRfQdgTZggPGnsZQEcu
qX67Ear6Zf7hEDyU7M3eAvnz92AXQO+tZKv89xxhT2W/7HsfIAuVwwBdEz4OuC2noqPkCWeer6B3
fWJGIbgxrP5GszRjFoRpRlUIO9FK6jVPEOYa7BTybhUZM9SQxgkZRH6crOxBa7UBbzIYARgOb4WL
MdJOc8FIaVKLxoRpqNLWQ/QefmlxODRmkC4sz1bFH2kIQHUnPmlK5jK0uvuRCVsnOdUk9GesStC9
1WldCLHbAvuanTM66jScGOz9t943LJlR0HM2lqodfF7wOCqfi/HsC8RW9XI1yBUx5gYIDfJr609c
R3WFdTnjwpIVb+qMNezZjSCbcK1OPLsacjpUwvr2pXlZPAGrGURzJ7cz4XDHIIvWYHLFuLCNXwUd
/Og9DblfZCQu08ERizuKp24/SzU1MEJK+KkNK4dG3UnG/6Cp07Lfyj9k9dZhn2YkUlUYlbufzdut
tp10C4mfg8WIqfEebqe9iZKHOp3iEc2cBTGb1OYleTF5Elyf1pZyOdGJMV+mEkH77uPKxHdQKPrC
n00Mc9ctYj8YOyCdt+JqBuCOsBStPwSfBUQULO21/UuDN6UEfpLwjPbSODi5sgKwx473wshg0ZdS
yPrr9WmNznzTIJi2yAVxRFPNq236+1JWTM0JvV9fZXjn9N/iscgFB3EQN4Ko5tBOQmN8KjIBbd/f
ZE5HT+lBuSic1yQltR4wOxyDdQMCDPp82QTOJNpJI0Yr17wb+4TgodkTWgQirgBhKFgQqBnCK1YC
ysZiQlt5B20hH1vBmkRArXnQGUl+/Dr8XM1BUVhk1fcuJoSCP2wYsDOqXR9ammEgofazYIzgPdhY
je1sls1vKMYZ7Y1GWRbnFQuBynEuDd+EuKs8M2llmpplcscKne3cmDq1ctdJMO8I2rFJHmZIM9or
RIPo9euwgOLrh08BBhSNQZufBdIT4ttmiHPtx4PWZU7MAzYdGovKSmsTJFneZ8xznAO75zwJYcV/
gU0nTLU2qHr96ruramM6IT8uxnbTvyhyHOSM1MogsNh/VH4r4pqNKwEsFawee7MGCXiJesOt5BgA
YGBbgGplmzW7Ge+pnEo0lwk1QwhyJ19GftYE9z/ytRFDQp+WRFCHktVZw1Af+PPJgcJkFzmTaZjk
h6uCGmU89NfHkSXdtYKD9q4hwcP0cifo93fWvGagkNV8IDs6MBN7Q2UNk1+fxeL381oEnwIZV/we
p+p78j+1nwbBylWLX8saIy1glSDOhogvVXedeLXdNmOMjAURzoJCywaYYtSkc2nKnwzXPDs/UDlq
ceNEDiwFRdB98qmPZsBH/Diq3EO0/AHPQvShqJP8nzrynGLt1m3auAXuHLYXWCQdwK2oCT+dtmfq
BZrEoiNIMltcc/NsX+u4R1bXaa8vmAzNP3Ml/klrGhdbeM/smHw77e2tX4Gk/IpZbzPWSWad3iiW
B3apXnykfy+OLWRJpkutqUYEOHf/hiCH2s1R6WGR5+eXq+KMoCCMtWxaqRyobX5N4RUqt5/eFeYN
f0ZTaWjZaeKL2AnT+EcNFDj06uYWvi4Al4+J5azTXxKrnBVPaEhQzLvbdnTTXWP95RhO+/FATz6R
OiKIyyoQWjY2bYkqSrevpNKIjGHObqE5jd1x413Kd+L3DW6tgCMnnF0v1ooa7FBwhtxVrH8IPJbd
LZKEZrz8CaPmMkncYlfr0e9wmN8vpQu+BlQc9SKBxk9Z+xzHHERLTiY0EARkcX31jlWUmILxhIwJ
aAqN0xjluep8/870FniZtvOLEcBs760DWoRFg0g3xykkJTtZ3a+jKpDfqvIDNuSO54+glq4zbjMu
UUxan5yogP3gZW6l1Tzx0RjstcdEI1s/5QwQClqTCjmaYDEh2XiOJBGIpyrVsBCCKElZfQRWPpQr
VMtdUdX4Nu/Z0SiECsmT30+QzlhmaMwKAcrXRfJZN1ZjuRMzcyj2F7G6Q8jSAUPI6bGBsDIQeJQQ
+lXu1njpxDoXeq6mH+L5Ah/SeyX1bDmJXh7GONE/cArp0FIS1aC5WHUGCx1b2EyGRHdOhOeuZWfq
t1jEVMklwpL9pw+vL4cHJVryWf0BrktQ+5pfmLdRNIsriXt8NJtqZFuoQkVxmVAoddhzy9yv9fCx
m57buNtlBBg6B8zUN3zpZ9zAupdlre/a7YwSTurkdm3835SSyF3sBnSWTuDraR/P9vdFWsxKpINQ
JC/aAXHH0ZBCxQEqL1C2Zl+8eo1afew6UQ8I6JHSASt/EwayhSn3lPUIb19DjmHW6yHbBRodt+Ld
mvGb/EpZR8Z/KdsDAcyFJGiTbSwXc1rNyAmElvjZnorYK0i4DdZo4GLbJPFxz1RGDC+C/hV4UTw0
saIS+IbVkBFT89O5uxhwcz4Aisyd1twRGAoJYaQRlcFSjAV9mmWCpuK4t+Bm889GAiSKrqno7X28
DUViyKqmMdSRuqPfcccJ0r6Q86RBMZ2cWHJUg8H3W98r4hxVbnhTR44lLwGBKOH/+3YhjtQJ2XBN
vWUGoGyUaQhWs0/cDNtz5LWTScGW8cXYuJWrSE/wlvGmc6DrTIQ+cPmYcw9by/VZKNAD3eLkssSr
8dR0zJ4/QsSPD7zO+2aALxys2HrMvA1nhuDsQRhVOwRvwPK2TQvDJ7Uuwu6W2G6tz4PaJLHuR8st
2q7/6pU1TYxgHWIIh7x1hk92wCQ466qAOHHgA9iQl/flcaGDI7TRtHkUllT4ttnO4N9UvJHlmmiR
Y4ugDm1GkYQo3cpmxVlHe8Cw9mvNIsSOQMMIZpZrX9QBkxUXeUjZw1tgEh+TZTiewGWNPYnuhAH1
CsWyMDI5kjx/Du3fxV16LA8/wvhQhhZMrqI9iITWELhILBgdYXR69fH8bM9XbZSyXcDa/5Qs/rhH
H0ZkBlqw+wGW+3C3AnJMZ5iPCEUSjUeFWfGnJRHxXA/akX5LmAK46pNijm24oCaV599pM3AxN2Q4
lhGY5VCZoAVtaL4FP/S64AnH4EXAo/hd5yndkdvcySji3FQMeL0RJfO/wBNnqxTUw41bWimDQDal
qGSDp6W0NsEBZU6X3bc5hhRX44vnS6UupOWmmoj/KCGX5uy8Wtcsxx0XU/ilh/ISFmsfBWkMA2l7
bSA/WXQwAPXUh7VZ+YsBj8SekKMCm7X4xRmDoa088TgBb89vYdipiNCQ6VRE/RZF8D16TzpLkGRl
EOvz+KjLFgX0lu7EpcA7VI/r5+C/2QNmGjxMkA7AkR/i07xhInk3nzrC+1qnVQqmN0IFQBspiFHJ
hBkhcLEXmcoIn6uZdiY7RJDsZ/N0HxcBrq1y9mm9XGu0rSf9Y+LYDmTyzDkA07mPFsPhmnWwcwBz
2FKvCp+/eN5zbEWzJFPtkTJKOMVYUb+B2fs1a6+TBkyI+0oPmRDuWe2FV/YsLGSbAzl9ysfPT8YD
z31x3ZbtkojAhpF43xqbKh93AXOFJaWf2AQVM2Ha8suHvjSL95M/OtrjAs3Ds9UnYMTQd9ubrC64
ANZ8m/JE5ZtxPCd0GskNvZJ1Drblp7LrTLLsR3FhxuKcrTPUIDigtF0qLcMF1XVKVgNGnAj+C8m7
0OHl4PLhmcFK2L3rVyDyBcYG5qz2ubai0+WTwUS1ZFbEM6dSOhunL3sIKpXOCWVbaHAG5i8NXVFe
higFwpmYMDgLt9tWHD8kKltpYGRr7ic9tYfdAyEtKRNH5IuD14bUBIe0B/RI/8T/sxLRbmj3wWrP
7nlcCIqsx49wIfmGQ3QJ1PWrzmEq5hhP2iF77wUEn3ANi2/snFZUIy2kttQVPjKuBD4sDLtXUeoK
U5cr2xy03ahPHOC/xfkDygWppI3m1CLHKZZMB8he9C4vK/Gcax66FIfu7EfEL4hZs6QlBVLd7jUY
OoRSrG3oBXW1Ieaj6mjZ0XYNwtBxXAME0sSxcF36ccsC9c2R96azptim1gRtPmbWFC7CpgEsQ6wt
4VtmE3ZwobdRYISiDmrR38F/+IvB4XNg2mRk/BInQV53cI+tNkf9TzF2EtAkBBi5yofhmqE2g0fi
Xop4P+d71URp9Msos6WTtY3C9R9X7PCZeJS3mDHf6y1RBrGSL4IbhonvYqEMHpjPI8ogRuBxCYRm
StUEqlfQhhC1gM6H9dJS9hCfYgLB5elqVz16yUiGMlYR0G0mG2UBm9FC9To01SmPDcK44pMy2/YD
aMitUADSwQNtlmSh3UT2MziLF178kL8iwODo0t+8qOsmTUSLRHQgMz1L6SiSVPX3FeZGVVTbSZdY
X5uR/ALGUtmrI3dilL0LmD1AD4ddDxkrXwcSYM1Pds5ULolEnKcC90eYhP2x+qWg5tOrqzkyY6ZB
RkOV2QluPXe+RE3GMW6oMx9FYP/mgY1ce1z80jQ14IZXtndDk0FVAhLHhGeXq5WMUrtS8kX33Rl6
3eIKHGNbhku3kYtI8JoFaaCfvWprM0yDHK72vi9hhLrmMLVBIS1ieacGksjkjenZy4KgoEfYzKyk
19Z3JbVdVmsoCid8I5ttCKzb9o9lA4ERi0tF0JoNm5qPJ/cycz955o6wDQnEiGKF13zZo8+5lFAh
RTKWuvkqlHjGMTVdTkkCwCfwflG7Z8oE0HLEcq7NbSR9QxTpseQyraVVh26CZULgZrPybEuUf80E
jWBWYaXv9TCqQ1KrAG+E5gTH1wWaixG4YpyFfITW9lLu66cLUff2uXHsT56koU+AEVaNxzQWbIoT
/t0kivmCCeDA6MXM+0rKziXilyQVcyfOefV4DRZ2L12v3iiD0FmaF2y7evnylyyiib7NOlE7O9I0
QMageDAA4l8Md1tzg0MxLhcBwD8pB6o85ajuvHZuI/+r9m/3k/VoiJ9hShvWJMNt3+tO9TCqYXaU
BsWIIoVAq/Nl1nGx5gTYUEbaIifUXPuU5nOhMY5L5vaXGMWNSW5BZW8IZ5NlNhADthTC5iqw8bUQ
uIQGSVQgBi0kD0fCrXmubWry7QYbntI75RT8GAtcVN2HnbbRK3MPhF6mTGi0hOQ5vTEnofSIauas
YlXlXzyTaFIWvsRU/4+BYhuTFTkYF6Zv0u8G2k3pi5LQUGNXL99bWcbWoRYWsCrXbKz1okg8mpsW
h0DNYLSQXYEQJ4BHRAp6BDhumWM+wd3BUJx1VqJeQpsDlMePtjgwlOQstOhBcrjmwIRmNu/14CAX
ADuuG3/21KSC3M7IDdrUY/PAgRSmThSngXyfqzDAOcBvxyIEtUEPxQFfqvvuZUvNQQLiaAqbMyGc
ObuoCHagOu1lLsxrzt3cCfMxUEAKEawKGIxYImgD88SPc/CveSDq4CNF7SOEjonI0cvjCkNC2mbo
RM27miCWJDcHtT/A1fdMpUxTRwxEFKTiGLEUSMLQTo+stUMo/33rnc4l5AZXGU2jPqHsNrm63nTx
o3ZjUJEv+OXciYH2n1FJ5dbsecLGPhWhgdb1y8z99IT7oqku+7nVPHS/p+IvTm3GWeopuNvzp8n3
pJK1YYsNzW8zyckvTGhEbmroORTksvCvxiVUrXwjPIhGjNi+sCTceUB2P9BQQXtCC7F8+SzF0hhM
Lmd/3tsBlBX6IqXG5AW1PtEMh+U95myMsASvrOIRsG/F8ugxlxDreWpF7G+dH7MuiJSx53ALjHyB
6m0AxS30pGKxxjsJZ1uuQYTlMR1YEioa5ilX3rTdiGsO1vTsAsqJBndLuKg+Jgr73T/iqK6Qf6pf
u+u5vgPlNS+zLR4hqe+cd4hWBCVu0hZH/WVYRzUp3aPBQZtZe9R+pbbWUcfOdH34oFZlgfxV/Toq
W13GhxRMF7bxwanb1c77LJm9w/R7Zh/sJjLs/gsZYlauufFIQbCCnHMDeBfPxNx+UUFnOmOF6GMr
LWukMOgCSt1Irhm6MgcBTbeiyEhbbFuOLdJsr8AH6adDRBRg0xysLsGiPKzNmdhBgqs/uii7BPLV
8dnhpaBMM4xlepJYyJ73rXMbnvjLQSdnataVWCxR1sbObGYueN7rZf581ZbpT13k2Fhi+zqezI08
KCzQRRtrILSpPu0AAb3rWmJ7FuYByk+qPSWGFiD58lRvOtUp1j8tZWvbYy+z/XZW4gb5knrhq6ku
39MVzONL4Wji19kTIxrdToq30RV29/Hwx/09xGjIA3qoGreOrljNK7yHsvnTVArUolGEfStbzRJY
Wr4ZcUU3GXfT5u0Fdk9nkexx6XT21qLqwbdUzoqM/8U8b6TRgzHVKT6XjWefdxLH8ao7XkQtn7/I
H5G1nOccTwZMXOJxGeMPGVHrYeBXU0BzDIDjgFTTULRt1fv6ouDK3sO/zIF3U2uNdNWfHNGyIpm3
lbNN0HK7QdaQD3f+jmi8gncFsNSqd4FSPEHl9/Y/UEo7drCPmg2zOuIo0lSJ++4mMdQkC6V6vOXz
FodBFxHXKiGcKcmkvYOZzvZg8wjDW1MRzPbgxVeAt2R8XAcKrI+iiig1wgF+cFYiR2e5gxXskKjt
6bSfGwcXR1QDPotKrhqLOtUclA/0vJj6QqAlNTF9SLqhGkpq/fnnLGESYzAxVV++j1Mur4I8t7mi
JgnierQPwLLKqZHy5KEgwA2qYVFoXYtFlnejqDr4bUKXyS0TXIYTK7Se50Yl+yUFyo4ezfXaSWU0
nsw8RO+uBpk4lYVFTcX6XDCPX5VKWwS88G8crV4uB2s+b5hXY1eWWhWe1IaZfk4bQClse38TfvFi
o+2fSaLyNJz6NwhMkfFJcpWE/rzZaxtAkb8hYd4SIpKEZBzU6J6t1rgMkEPfdEqTdB+ccBqGfLzY
YjQTskoCn7u+ruG/3sWiOwGsqugB0yUWiP2eyo0nF+XwK9tT4x3TRg2CJaC/u2ONJQz52aWQrzXU
dQqFNBitKmPuHx08oGKFq5R/4k19j5AwnjQMnv2Ra7jEeQFtHEfUYx9kAOe5vaUJW90+68I6IWT2
4EuJrZAOXIZTJ53ET9KtmtwBCy66d3z+A4XkIfa0f9B1P5KE2uoheW4/S1jRK7K0B9oK2Kb/X54x
bcrd5jHgl1pqmOcpCzS2hJWCs2romrnjtwxiI46Q7zr0YW/4bW+IK6fSl7Q+5lkAZmjecu3pPcTw
/t+56R3lQgUzq9ECs/yxxKuJMyyMbe99aavqoAQpb6GQpcPsbD+nQy9DDnhJeMKzMzKg2PEkYPoP
CjhIIFIbUA4+kNHGW+Y3NDURb+f5EN6FtiBEhCPJ8e4EK6T6q89rxlvG0KrwS90pyjO/tgA6bj/g
zvBKHUaabzEQVr0EGABq6FlflTswAUJLzJzS9Z9B5YUo1pQN2Ga37HwsJfNXR1+or29eVH1J/QVN
F+drdDO6LHbIqE30Za4nSkEzuT6QhjzMNzInoHe76UggaFAPcAgIOY27v4w5OaeaZpW5+grGS99P
I7+QQ0oSHuF4PMdbVRsiQP2vcFCW2jiTIbB62CGmYsVKI6k/qaYgBhOYKq/WUBhYUYiEPCVPiJyM
k7nkpT3T4hQzAzUA6+iHxzJMBplmb4hnE/0h7VVAlfOtH+1xedtTdvAEz8ftp0+2SkYxjj5k2oxD
54/bPPY7rVWLrugLImGLY3yGLmmDupAgYztlFVAl/CbFJnKCFkvfyLOlxNXnfjILoAvBZZ3F2z4c
mOyPcCXBD+OOc38MTUztOJY+5oqz8n9iEcvgnb+k+Ge1ScdBsPtQCWpbqtOemzg5Vk6IIjUz5lN5
xsmOmVjQg2Zc+BJYT4XSXru7iccluFEfqLv2vRsnR590BJXhsF780wNrlaMynclgwP9vbZNrm5NY
XEwP3UGJq4zwepo5CcPCyq2/G9Yh2pOUD4uqbuuBN7eTIP44BaWhdu8s0FSAL+xkdWp805x4LeSi
qERP7d2gyvx7xHk5T58JouJLQhLxIK3LQUZLj8lMo9h0e/VB2LMQ/aypkCr5hOce5sTM7jBiXsXY
yOP8FpUc/8g7HuiQdR1J3K+XNDcdFYPja1VUgt8Galv3/BPGSYMVD+QjA1GED2+GiMUzkTxovbKd
krp7vOjy2q4hufbH3vNiAadL1Nhkl0g9PGhGDuGNFjRGJ7pHtsm8cXRjAcD1Wf7b+5cL1Cipby2k
wSxejEUt+Y7G43OgndfnA18JIvCjFTohG+f93IAKSeedwLK2RnQqhx5bpa+VGv99VfeXRtGv1unF
PyiCPKVxZ8o5NgIUandHKL9fspNTcoifnF3JIg/AI3WjqdAIXPoKm9pt0nXztpJRu5mlVKymp2vs
xRvOEW140eGJoOolz/YI7qOSMONFtYWorBmUZY9DXiwfBLKgUimJDxBsgz8NYrY533aqVkU3v5rM
wXvcVcvku0tW3io6n06R7AmDSmwWqG7aJZvmfp5RmN8Qf+7TDOjnWEYFxMweSQn6RV5bhuilE3Gi
BHRIa8EGFi3Mo2xzZV0C8ZczKhGe80CB2ZcmCmXi3FlwnRvxYgcHDLxY2zHWN0+9Iq03Io5SU6tR
/Rme+d6tzRl79u2nYCHJAUmIXOoSYn5ONqAGsNGK2pTdFhZ6l0UhP5ZQyTdjpe0MNqNgEWBtvrpG
DTYkNubtp92FePH3IV5nxKfAgv7U+YFohjwgALWLUuv30Gba438bsdWtHjKBwb0woyywlo0AMmys
Zoxxj9pQRMCtgbmUVgEK0qqfNncqDDc1buw9B0iUz7PGAnhLtVlmUrYwasBym+5ipjEgeR7nzYbt
RV7Rjwy8q/yBAnP1f1adMJBR0SDAgmMMPc/3hYzb3mTNxVf75PjUnnFEaI/SZROlI1FNBNNm5JZr
haox9T1FQm4Ou65OPlrOJORrcH6Xnoe1P6y4HjpazkIgeY/+Et73VZ+76xPhJM1jayblAJgolVcp
G+PQcG5isKBl4eQSICfqGj7Hr4yX9devPAxo37tqyUZOL9I6c6wwHUcKNgOwA0zAr6Q0myi2psq/
nf+aDX4X4wXSePYM95onnSEM8JgnrxvBNen4EEpyDTvsWo4nAZXWvl7zycOUglRm2b9ZlguikUqQ
qYQgFHLfKv/cc7fUcqv/r4pB4LOMuEs5yH8aGC//7SNLoCFYOjnQhY41hbcIb4gtfAWUBsIfJgkt
rTrXYnH6qICJW7vXfBV5b+xtV5kRneWt/EcgLKSo8Exo/3eN6g0mz0ebCd6X96fWFqwpdbAVmSvI
apwbjqA4P9QuZyDk8tTkPj65kGs9Icy7wsLY9dgu4Q2ux9E2e3LyLtoA0JDEFL752HcFw9ZMXIIJ
QCg6jMRtH8QHRNQBWTj7gzNppseqAlRlpLLaBexXNjcfmb/XA/nI64MbMThd9XUp1umiHPKoVpzD
PtJoBBqRU6FhT6iPZwLFeHk4Hxqh5XAO1FkHkah348iMJYqY9+a8HoVmyodWkKHfFmdLeQKqC3qA
8jw1KYyKJ4gcVXT+FgOAlowQGMxHe/3N+lIdXOj/9ohxUlIMInllN0p/Frx6h+mDGVLYXIrs5IzB
0S5RlmjU6BQ5xGjhAJVYSwhjuO3oeLru3u768pnY0gHkH15qklc7rKVxqMhM0GujurshUcM7ypAW
oyvoKFIx0i3Fl6nxw+tdDPz7dhp7t0ENu0cbxQn8hH8KnDQNplEkB2q0xSxVVXT2bDdLINPAwTmK
45P+J7gFBiZuCaxJSNmHlZ9A+T69KLVhaGYHn72EPAWzaYTBuVM041gVq30Jjc2mavMXKJnzREKy
X0QTJtpDtExt9y48SFqqYOIOrvDiL/MwetL2vEF6nVfiUSrdTrpowZIsMebTDyOcQO1JDFBXgvO8
c4/EP/yTdK3BKgl80+e/eBj3houoNqdH3gEwaje6UUYwkydLe4AXhxjmnuT6A+zxaFA5YO0jJGYR
1pW9NJ9XhPYLoYUoPce0dwqCbtlOBevlKJI+1+OkEIUqlYUjEcI5f0aGkVoCQuCSAQxHjbe99kQH
WJOyqlRncv7508ED2o6dUoEPijZrmBQExvj+rKuK7bG5P48tDnOdVvZi7E/9n2f6xXedzA3NihWA
Um6dlvdvTTLUV3iG5fvAQQ//M7Zy3uRPWQfYETGcfwhA2CppQ8x2BMlDfabfDnFTU2AZP5ZN/48f
upCzAzjPZCbWn3o24aQe+luR5iqeANMKmPEn5lrCqcnKg86IJKjuYpFzQbtXKPnDX9Nip4kc/1S5
AYGeGKKKKM6fK3y6ZPJIL+sHE4T07M/VW9YvQ6wb3MM3By0Vxx+6OomyBABcWVvNr3SzbB307CgH
BN6xG+gh/DnIWU05sPJOl+gW84saXJpwyA5LKyk3qqtO95HTPkyXiYVIg7q1+jOv+p1OL1zk16og
ZG0AqfG6IDZUi3kSTBI+j1oqalmV3oU9NOgUbHPsCjh7VhQc/ZIzUm0A4FUNSMCSOrsOPKWNmMci
DHpVHcfPmSrTypGmWDHUaDGNR2cC41Zn0w95PcJu90B1eaOPU8me+EqS5TkogcxlBDqxEiDS7z29
ITJwIMdEALDIe2da39NhWbmH35/fY2DfMCtnbAlDO7HxdweTW7k+nO1O7z5QKZXJ5IAO8iRjTIve
4Uwq9T7zg0/xrHpfllRQOQ+TMtvF5+lxy4bPOigcoxwO+9DkdjSlVQhvxMp7byTktP51Qfycf+7O
VADjBBpReEqRzZTjTIgZFrKoROfSlaiVZZ9+idOmBIunZGTVJ06ja6z6lSgAOGnA8e4KiOGvWihp
bS8QP7q59E46M3hD8lbNV/HBHm0Ma+nCtFAgHR2UMbyL4LVIgJUe45UfpOv9eiK2l7kNRyiXKfKB
OJCK8b5EIF42vAIUlpg47HBfoHmMPkkKevbdDTvzWnKTbsCrPUzI5GBTmAPuLL3F8UugN7JsUsRR
S9YND5wA+ee5zI+DD1fxmP0aYi01ZfFdhLK27Z+7EmxtkkfP/4Icbplt5mNu5yMgSwrugCOxcpK6
tAAqMH+WcnBF96C7GnKcvCx/VghrWHwDWmbmuVxS98cG7Z7/k1ZVkHbpVFDzEA2l7dhlI8ghTV1E
HZiwTZV7pBTfoQshnXRjW7c+5yLLjwfqckoID7wdGyL+RFjt/hF2AD5VaqneN6AZGf7hh4lo/SdP
5xAZ9wS/WZsjUZHmEdciuurh0edrXV3twelHLaNSizoDUD9jtQ5GIChVSm4XZTXmxJRE4dq9S347
VT3yNX4gRRkD5dAKrxRG8udEvHRjXSDats7yO8PzZNQsEqK+nBLZzuyO+KB9XLIP4flk4Bx6r0e6
wT7Aq+RITYiaq0Ts4SRyjxDRVC5kORtQA6f3SF4QObeQ2sWuhlylXycMFwLsbgCSj5x+q2MsvQTV
EkkJwvMvCKwCDJW3c+A1t9oxu2dKzRE/Zy7s5lkiOnHiZP25UlZ7QwviOzJPolrCO4fUSLt0PUOf
XSa2FVwqKvHLyqcIGxOcfGh7NEI9VmibG6sdwM3cQYc9W/Soe6d+Gp3pl3HqsI2VtYn+EK/CdgCh
Rcd+3RrSOBozmVPlZBNcNLExmK4PGO3blXycusWiB8lk5B/1wcSnC5a0z0f8w0xvhVwCZsijdJzm
vyK7PC0rQrFa8FtQIDfQyIxsEs+EkiTDmyog53LVXFbFhlCLG81mAsU4P6cGyfs1c1K/3beyUmqB
r3nxY34o7U+TI59K3OZDXLBJNBkBeBJ3LM5e9yakpK4KdEyUY5I6c3wlysBW4AxM50uBn6g9vj0e
+xONxhgIY5MZceEHx42TE4XUD0uLBNax5q96QYDSIGpaK7yVp3yjDw1BMDHGk4khiCx80TeaQBaj
kwM5i8Np6Itnr87MS7p56nq5RfcO+JpyrQBMPCMzkkioNgsngefw19V870ASIX8bxYyWiap97siR
F0JuGdiVvYPDLfv04jEe/7Cr/3PNT2GWSfrgr/ZlN6kQQjitNjAR0jQH7lg3QfU0FEzcvZOkPRai
RXkEfFIFdjwwoWnn1SXntg5WIYOvqxLHa01lC3upl0cHiNFtJLYYbh5I+eJwyKTdSUP77E2c5st3
fhT0ZS0LRiGIr6U5oJxVxTgPNmE/kW7IyWRKbRL7JX5RbbdiMetlXTxSHBGxpBDkuaZwjZ54wkzx
uiSA//hpsWyYe0eOGD1GQc3O0dlQZC41Oby+QyMg0OpxGBt3PAK//HaUeuCAyLm4ORa1UqDi1NL7
/Uk/nD3biSoC5TuClxhWej20W5tYvF5XrXRTLMubMR/tbNfwGtbq+sp1pr5DaVWMyEHBdFVXHp7p
GptKJPlKphwQ3CnNbh1ValT2JonFkdAgS5qdsu87XtLHQk3s10Bm8/RP+EByovIsUzcKrNNjAffm
NtWshPYwa9f39TY9sfczp5gdNSER+2Z/nDwVA+8GHCDoxfFU/jsBPsNEYC00ApBh2aynmeVmddo3
SC1jxnVYC4RdJyLmt63dM1SZ3dHq60icLObYoE4dQKU9Iwqqtgp+6klW9gqB4au2TfGbnle4VcdI
BSDnQgt8NJ2Esnv+2vr7Dd2J47csXByZKcNUABomdcj+pTONuabxLpHORC/dURnT190vW76tBfnc
2EVrNQklDIkMZz3CYT75Qblk81ZJpuXtzjZyJMvQ/NLDAIIxkh+EYAGS0/XG+7XxJPDpOSKflYKz
dTvmEmchZ48BJKBLwSz98FcnDlFIS9Jwf7MlSsPLbl+QRmq7tsfkY6Etwhxa9Lz7hAvAJJrMrtG1
B4ghrfBZlMEeHuqOdbes5MBCHqkA0pzMoCAZ+Q2U+pA1hCxWYiBQmLzEAV6DuN3oEUFIekVwUynU
xloGUN3sgXOBByV8dOqqsh6KvI09LImpyQbvg/x0uxTBEWiSfDRjMZAY9paA3z3Tn3BbZ6lYIjue
02AOK9I7tQ7Tcpy+OTaXwyGvxjh7HAssUutI89kegui5x8u6jp+rgxp8i1fmhMj5zZJqHg3oRnX3
U901tJqcXvHHzjhow0G6l4ocmwuZ6S9DWBvnNYZbrqFuYjvAu/uxNBXLfLAXxm2knJjzvSVoSZgv
ryThZFJwB+gdsOILBKgXo2mQCR9PxWkjfkaDvbvUervxte4+hFuma1neG22Bj6aSBAsUapQQk3FB
7iZ5oWynKDe/ZWDI+zvWRfRtTMt2Isf6qDucbBnNo9FhGDPq2xnCInm+8afwpPNDvpKdyJkOMynL
tGexI84MnKVA77YQ5/DZPdFiDGcD9niwNW6h1onF8br8pscyKAslqMH2w4bflN1og8XWQxyVGzid
Up3USiAZWsRZdm9FrPi7VVXAeTZzZGTS68GokSOUQskh/wf89BKSqKsjw1+ku0XVj9sR5sE6FT+s
O/HaCy8dA/ep1pBJrUiEpwcuFL6l5WQ7S+pHpBrgEkTtxXmAMnrWoykI2RFA1x++Xzav9840KicE
zpulRAhNgxIjzkB+ejsXuFJ5XPTYXAEpC8+DCdHVHLWJTzUDiKknoDGu81Qa1iGFjD0hvbDm78u3
KlxW862S+4KALOTtFYNJsCtws5x0TxdaULC/pW7PX524hf2QJfHpjB5j/v7QCZxujVLiIF+3Q2wB
N0RBh1Lzm3BYVcmUKF1qaOLJ+X+qt5kJLxG6SSy0Oh8jtEZkGsg/uHO14xJfyaU+ZmMgRCSneqH2
iT+AHKybZ6RfUROzsVFYa+SnH8qiHPlm/JDJGscaCRGk1t5kFF33c8Rvp9pLL+2jWACdXlwG6hg5
ITtt/ZwNvfi2RCurlhdeVNO4amIRGtlVMnbr24X1lvj6AnulwJ6JD1HVXjn5k6reKGfe+IhAgxDn
H6HVOt/yWXJcSZz6A5a9Qqj+4e0yxlZjiFYj9IDg1mdCkGdrP2G/9SPm42sq1xKITxzp9OLmuvGn
yvUr1Dw9v5HP3ILEklvky90VgucS1SJ4pxVIrJ6DMYM7oOrxyFb9WiXYAharXdlM1NQPUzGPy4iE
lzX03YiI1M29svubRUqR8JULW58kItrVRfGA7ftHdzJROAX01H3lOGLv0ABHfigpRNMN9F2YFIbY
/fWWb7zeM6HyDd6ii3R+hwHGn92vkQA18ZbGOy0sryiQrK6z/kmGU/Jdtr1PsbdJ3TQuFVif125s
kagcAz3ZuLK/56LFn71i38C6+7W5+Js/74+QbJVZv/BaABIGtjgBfI4BVuBYXPt0usuGetVgI4C5
bhOBMm6DApO1I9ElnWIcOSFl26G4X+5lSV/AhXCJjue1DgEsk/7o9+dFHu5ah8Vj8G7G4cRPo4so
BGtXsZvwyIiyNSutWaoTkDNdS9V1Omm3G93TaslHg4MyB087GphWRXiN+9a7wJTwHKLi9inafnpC
MXc//No6AW1UXdZM7Dah5Zkp5uOG4H5kuA471ZBRaM4M2CB5seh8RV79e4nHdLy/r7oZLks+3dfL
Rp6LRSVIDNp30wiDLW9rdMSE/uiGfHFRrKIsccZmt47HNzJtd80zQKMXCd0yVxV7emcppI6+XxgF
LFZbWWw+eiBnLtfdK1F7n7z1Jutb/Wl61GSIls8FS1bwEynxswFdN+MFhcoUyDHC+fWot6/UCC0n
jCbCUCVDyn7s01nBxKpcK48QjOs3ERBPNo151Oqj4GuSfDSsZ7/mtnWDzlvE3eKv0zgi1J2ZVsTg
fU58zXFgKN46lTMgejRO50RtmvZ56ET5W8kk2eRfqIjOp9N9YDeqPuifgJDMVIUT1uswPyN3m1sV
2n7jdXGAyz9pjzwgs6DxRpMSrH1KpqElvBZArXcz5jVVkhdYz04Kh8vdLqi3dYJ1FpwCQ9UPvAb7
NDUe+mItjleB23yIqyZiLKnpASLEY243B/BUyxNuRh5nLIbzcz4DQ30+4oNTmDsUgdjZeEvPpfUB
jkVTrKURIrmexhKk6ymjWL7EKfe+1sF/gemIhw110W6or5CfifgT3xIT3IAN+BZTEamleWc4NHvK
xMGo388gOQUeZV+DxdlhVagtZPeBQR59hQRzAKBhBqojSQTJe273bR5VyEpiZdnqpSYlm5biOGSq
099C7mGNlEciQYnubh/A8vvfI5ArNuEZq6EJqpJKOTussQg7FgHNOv8PmXDyFnClML0XcqRpxHH+
eya4eS44AwnDx0+7X6vwx3ybzjhtUxccE106kkBJd23iG3PHZLUa8A4rRZGJlOv7/r5rRsahYnK+
qVSPQM/BrTAc2vQy+0CPhVqKc6yf0HgFN70svU+VAA0xYi2R0vglequnyqh2zHXxL+JcjjItwYdD
knyrQLXqG8//yzL7OsS2GqqKf6fPur6i3L2wolEDMpme0m0EyZsPJV2VRDk9BpLq5dZMioeNpAlf
LAyzK7lfF+2/BkI23OLK+ooQoUBavX6WuYW/1175af71VSxL9RhpZPM5AMuAxIKChhozmbir+VCx
HkkyTowwh7PABjkr8mkOon+lalzVINL6fhG0DqWd+U9vDkr5xiuwVa8SjZsFlUydL/oLp/m1JmPA
qDcg6lFKx3ka1JGRqTnjOC7ZhOqolLJ0cjyEDF7fWElhT1BxzwFmqa2ctl5fa8OwkP6a+PKJ9SpB
nVi8ghE2c2CGPV+0L6pbX/QIBnAcrZEnw4cXvCBgezpdsk2kz9nPbSka+tUbzXVEmDkcNnE2kpNU
OMz271fIZChASRq/fOZ23A78dofXeVvj1T5jUOJEExhnajbJG1+nxPtGk6aJ8AiU8olKBl1TDbH+
EtTffCrhCW0LxpfQeynSOxU7dymErR40dv7bEH8Y1inku4Ut8N2h2udn4IJSVg+iS4VvVrHwsND1
z43GCIiI16lYxLQgGb27l+aKFhgnTLqGHwIU+k79SAL6itRWBAgjF9RfQbsBUOftBgxBtemy2XP2
Lw3B184IMUEQ87qD1uDBulfb+e5lg7a/qdorPFp1QPYznxl3pLw36wS2exnFq96yYGSU82hLMkiJ
MmegSZrNH8oywQH10V96nfKAWbP+V+OsVtZzhtanbeIUVEwSwiwcDkesbhb+MOxjXRc2FXfwB9+2
ovz+r9soM3KkMH4zli7tRfba8uNSphATQjTNzMRpCPVum/riIVqApMcCYQCYngbSvV5h3H8scrzy
5DShJ5sESaDnu55gHzZ/Z52zzQbzkCaHBl1hA1j8UuiVLd2/NfxLeOVO7Lk9MODf5XZYjo6T8H15
skfQ6j5TVHiS82hwkvZ3UqmvCvc1OjT3azTPAptAs6lztVD9I2QzjC47V/BwdQ2rchun2NZt6W5N
DudxvsseENdw5IwhvDg9IOElu93p8zwVy+MZmhap6Q0t6ZdMwvM7eNogAxix7nULvXAkrp8NOJZr
nJ7keqCEF9mql202Av5E/lg9H8Rzxyb9G1ZIpdqKn3ErfS04ZDp3lkoDp4jBY6r5WJKREhX1xLBd
aerFHPmSSzKrW2LX0ki+OhfpL4YdXyLlo9bzrACXpiJAuiI7I4mJFl7hfVRaAwoYz5XqgY3pPOZ0
Tj4WzY+Qr2BoWU04oNJKy7FTjNS/CtCpTAVXZkEz+J6pNuUWqE4pOFZ3peSrOCXRvnxStW2xyG8/
MF0jp1ugomyRB4UkRoMSfY2gxVZzq6TEAuWTFwlYWkFBDXmP8BfbYxdZNzz0upufrs5LcpmohSw5
eRNgFnfpS7FDzTpbJDxVhB+IHlfA8LmcNNWsM6SXcRTkmmnrjmmtTpAUC5WN1W0y9zKk1c7/+Rol
99/jH0bdzrdymK6sfM7Pmhtp+80Q7TRl5jfKTg/jGxmvSa53mHpIKs2GWqEzipOewW5IZiKIRGqy
y1XwLac0Z/k+KHZX89wlEsB03YhrLz/wl18Sog5Bhd56onN+peDlx+QwVdyvfjGTw6wBCQ3iVsV4
EeON8O/X8NMGFwfMWqkEHPWD51yzV80KoA7FF3IVwsU4scQyYVtlQlb1xJSNelbUYLR6yElQPv6G
DtWjkAKBsjMveSRjOhaZjqDWUphhodRuBOdjLA2Ps+zR9y/xJlaa6wt9Aei2SZUO8wPCPYMxXMcV
Cm3Ut2GonUFTI23d5y9yslfRB3bKqi7qnWXejpk0y2zj8ykxU8uQ2WECjUgy06XRco/nktNKhTxY
BED4KSu/gHWlRTtXzVpSKQcsCpuBdpwdWghcyNDAaLC0j1c5ZTd9w8qoiamraHxETHFFb4ONv/wO
6/qlfzUqsZoAq4v1lTKhKnoQwAtIPADPV8MM0mEtlh8LErkdEC+ZsGdC/fxmeXWbvgrEve5z9wGs
+2s7rg56xqB6XAqnIdxm1FqbfdW+ZUGgw3bN2Gd5/K59hdaS5x0swV4Xy++34MZ3r3Zo8Aq+N8N5
AvytGmM0u1J1sDy6m3RibrBDtLjHF0S9Ym3w33coUUkuDoUgRXS8VbC2mgtmtPMQx+gDXpwCjkM+
dgainj7ekHBR846ytYAjLgaefaGHDZIaetAuVXHxNwOdpXlrkLNG2SD0Nf7cHLFdGoD/HQmf0bjW
Pp+SLuLDGtmTPzs0vS4HNXXQ9yHUQtluAN+DsV2RO3uZ0NC+9gb3VIOwW73L3UDMlPfJdaoZR45O
6JMXLY7IdkmDC1seLZRazvZjR/fYhf+0NljSbTLoGqmxgB9t9kHJeeV+YSQLgj6Z2Gj5/thFBO8F
ntQ2Cgm2oIE7NPWPWJ1FmmW0+LrkypqoINkQwlhYzAkJyIrmKvb+fwRB2xDn1cephCneELdSlhXG
MhYMdotdpQo0rgQpc2yRN2hrFvT3Tana7HidLsV7MUrGYE2Y92q2kWfLeLHCAmUUAJ5zggAZUogM
83wtvJHryRV2yzCtdKVRtCr2fNlURjOD9jIUGcjWOaL5BYMgiVXAPF6vuwPcsf/DBxw5WiijFrdu
2jwRYyNvlffy93tjBkWzJIFON+P4C2Ix8HuoQBpzYbKMMj3+paZaHd6wtNWBRl73ifYYVNzTfvWn
78WmRp1xfjTxNo/4Be8Ri3h7O9dy2B7ThXPNbZQ3PEcx6Uv7Y2hDg9sWwkSQnNnUggCvvY1YsSq/
UmXN+jEzIJSDBuoGim1J76WVi4ojh1wv9AdYjaQuYTufUhPI3Or+/RXkamC0vuj2icNmRF8WU1EM
cdbwGQQcL23pqOKQ2BZy2K06EtiTai2A/TUg9z7ix3PztGMZ6WxUQjvlhbib2+/G6r2I9TYU8ZNs
WTojgftx0d3JORxDW/ukqQGrLuFkhKNepq0sTouuGyl6QGBy3HOCW/wYG6JBTfSDkM0EtqcjsuK+
jhCflfbIGUsT0/Cgq2fSrdgiyU4ZB+BN6Bxz6BQxHFbAwg+C2SymZahFSh2zINmjia6KhaFubgYX
QTDdKsN6+GbhER9dQUsvsG/OsbCDRr04gYGyMgru9gD088hU4tVzLmWWbfS8hyKHLMF/tg6GS5yk
a9d+qPWOtCWT5iXPOqTsRJqmLyubmZ18NLSZrY044Uln6pnRidaanRTHtdlXZ3zWPxOeE4u4XKSM
7wastxDGCAqC+9xG8UDkvBFdQ6b/RqGcZrboqOTg2uvLL73+cLOlcGPe460vo8XcdtaleKWDMNfY
f8otyr95FK8BBCuHEVlIeqbn3Qo+QbWBR9jtwQ/tyx41JFeWXwqZqXELbZmi/jB+Q6S/eE6oiptW
1Jq9QWtwRtZ3d1m8I7nXC+0XIC/GhovSWJ9gWxjuOQF6IA+iy9dWCRSpTWcqOh8kA6nJYf7dY+EX
jAV5vhfW2i1FGAUbkRQFs4Lo8AgW27DqxrE1+aTnGDLw/d/pstIaryKN7XwbhfNQ1nzfoN+xCxBM
5KKNetiuma1JNNruV/wpQLJXHrLULX67xfIU05PNN9dk7WWdmeEWdg6gXGKc3i0gF+vboKztNKvV
/45yzI7Wh5JUseh6ci3BMBSBMFEqAiIW5erradnrhjUdibbftv//bjL8ycEE9sRY1z5OTpwpsDhA
tUQD4z7gfPgUKwQ8MZvs9WU1X91AHHTiw2KMmDCG3AycGRcC7KnIUoitW6B490QxhEVP9BQw/umo
5NCB8TVoKiAtpAqrQhrBCf1s2piZj2F4J3hU4w0KNXgI+qvP9HvYMKm7dou0lgZUR0gB+qHRCw/p
2jvE6ymJOzh9fjhl6kIyXjm4cOHyLBHIwJbFiNFgARtzxy5QUBE6W1GmPfdI2QjReCEXbI6+ZiIc
euN8kqSXX7i1SqnWkEBVw4e1OAcgFiEw2OyJMJcnJwRQTAvjewyeL8FtljFPtPf5hnchrC03/h8+
X7b4MXlXCFZZmg3jgciRfF2PkPaRaGlqql0VZ/cqNr/cthWkxAXvjdNAahxaDEDHp7gqlonjFMly
kYH8M8W1I9oy0xu6lK5jan3EhJvBo6NjA/BhhaKbcIEhZclq1E7TP8MWBX72SeePByByBG/PUWLk
D0a4K9bdPm+MDOZE7B5vUZcrF0n51L/AMLWsNr/JEV4izx+dvi1/mPibygHvS9CzAkBNlxczk6W4
jM1ApsT2SMRGRB5AuT2dn1902gQNnr9yaPrjiZkuxVZ1w+sV3fTQXiC1C28208hB0eZGMlb/29hq
+msxf6Wi4CUXU6w1H8SRiPL3V+iX7c2uiO0VpTNtLwDxMKyuxQoRxZ9+YFKnCsJuV7Xf9sc+oXF9
7pBQA+7zXXuIjgG/mB4i+YL94z6QCDpxVzCjCtM5dlPtq82gifQYQcSokzcD++S9iwThpHFNGFEF
JJH0m17bdSsDqrRoVu0kRdnTeQbog39VVzh06JF2TrPfTnPUpQBkL7rYbqDiVcOuSiEFPM1ivfhg
PKPAxyBMQ8X0OAXL/O50Tnr+wsqKKx7PubRLPPwNuh8A+7KjZCie7WA5sS/hTUBTwJksrdNNJpJg
I3I/Mcm3EiAKb/xt2BWe+7GtXocvxqb1nEG7WiwbEQ11fYq4MuAL3Mnm0F9TNAjuPUnbJUrfICZh
XB2oLz8C2wI1ftN3dZLbxEmAbkCBI/r0Mx1SEQef0k18X0UWThQwpDJcatJhEtCg/qR6x/Lo2QKT
HdhzPJYGWPSRgsQDa6esIgn3jW6qrF0RK+k5G+f/ttOYXib5+UymGBQ0W9G6p0kDnY9HCLT/vztJ
xbceIF9EBd15jpFnG1bKZf59STHnM38lb2CXdTj2WDQT4Q8tGtVogkietypoiJgLM7/Ma02c3iI9
9EEy/QPjZwxoQuTlf8CyGDmE977Kyl3PWUh7J2rGFKxZ45vYDuLw4og/sTukN0eI/sE/xzJWG/bX
X2rlqd5cUmlWVU5Z9q0fi8XnhnS4R6liyBEShwzOhd2/4w5m6T0HQ+rIMcYoDZaRQNez+dZwAZ10
7LpGrGNgvuHOJYwWU2OJYREGsLpsGxeTA08zeTHUz7OSl8AIj+U6ocXiDAelKoO+OnHq4VLwqllJ
bGi+XGscOqVLxzAAp/er7tLQorI2ST3hysxaqpbwMAdDjshoi7F/Et0Hy/MCVlD8Xf8f8STP2DHY
8+0gJwV1Atuy1dxpFwwXezTwDJFq5J5v/kVl6xB339P6hkux7JrGOU24wPKgKyWUfxgF4wK97yPV
XiGVnJsxUgy8DnnaNbxOQQ0LzmsQ0ipa5Op5zkeJBWLPIvgWhRWvFwvvHp/zoCSsyTq1aOEli3lo
wI87Artfy05PbNONanX7ugCJV/RmmaDLSliVNwKdr8L/9sYQRmybjTd+MaxC/ESYa8zy5oRXOyEa
RMuPJvbQyhDLiKygGmD58Y7IGS55KLtzdGfTYndxEz6Y9BlsrKqIl11fGIKsapcd9Y3BdDoJJBoz
DCVzywChMzSMmCjmX5sMvncOZJ8KhdJB21qwOcKZZ394xcBMWX4V/WM1cVQIELbyqPP0aqvdyAHC
QMNmYs23gHtIj1kn7/8K+YpZfUzIIhdH5cGI3zfkjBJXOZIfo0XeWPKTdcqUIeAuZXWAZf6leTZW
DLJm9uAz9bbq4f1V/sFMAFq6wp+6M/Ip2+Y/qjr+xYXlNZc34x2/Y5TLxFrqgSb8QdTUadoqwIcC
GYBaYCp7JpyYoI8Jky28aq41H1WYk6EB3BYJ0EWK8hMmvpeHsVmUl/P+/IFiphNSVZ7r/jlFuIsH
NdDfd7LBtyG3sRnCPe6eY7uyvffnkPltUh0w41Zyfkd2bmzTpvG33npWttswJhTMVWz4UO/0hzgi
WvhllpT8fEro8zGhMDkhGUjHkHt3r10AUoQ4Cvcr7dm/Mk/ZX+Uh2+y6g42ZFdGykSZ2Z7fQSmY4
vkTrh2nDbMSQRvDxE2E2paMZPw38Nne0Oh7roAxFkYF4WrFqW3RYC7yrKAEynLTwDzvHoeSR5Ei+
HL4MMz6Z25ie2SE+Jfaq3lUNuyX0TsHC5azBnVJfiyQkXtO4k3xp254cmm4hghaulzYtf6meYRAd
SC9Yp5nJTE6rPEcihaA57jmsaZMpJyJSf9Xq0EfXEQRSv6XqwGo5UUsLFOtUHoYwsYMj2Yn9zO/Q
cdCdN8Lvs2W8tmfGPMTQ88XsPsLBydwR9mhGhufuyUaZMVfmA/rQCOm3qurwffl35EbrFrUSaQ/v
9luw5XnCZbx/jLN5gulDpsDG5oMstP8wpGCcFB0GQntZ2Ejvtd2a6oh4yN5dM6YsOgFp7m7Onfbm
zUa3O3Vc34vPKMmaAVo53D2hEwRusBUHBuWy9UjQLSlBRzuOEYi4ueWDaXzyhWtzTzyAimbSHFkk
CRaWiAHb8u8EmFB+K22EwijSnWH8/EAQ2EPlTy2lWQJzw8xAf83KyUrc57lWOQJD5ApxTcPmkpBB
KyUr9l/y8cFbRObCBZ2zWhBm7PLCs9CKerbOgRufx+Yx1aurP0YLODI5v/pUGg2657XFVwV7zro1
x2ENzFF09QL7MjTRkOOojW13IFhCfwAmQQvHYijY0lrxikAsKIzBgKNVB6eczUS9JO9pWCkHiKE3
cmnZdW3lCXh9kssysLGnc8ABpN3kk9WfxIdP4pl0vqQ9QhuYWb12Ez/BYmHl0MBJEGSVarrNUxDn
yezTxFwsAv0omuzl7UqR5hmdNcxlz6tMwhhk++oC2UCQgyU3DBIcHXOsC6iGMbMAEUnORTC3PTjm
uMdq4f7D6kX5xDpTxh1i3e5XM3wXcWX8BFDbpAiOTlAh0c41icyJ4NZJNqfizVzJ1CBgx4hQ2nW7
8qXjqC2KbRLkFwOPxcwj4uNW2yQUDL7ZwiLDFTN0bL91mCtPM28fOg4mnTBKeoacnjTdIwUbwR5U
Tc0gB+aa8by4mjHu2hTIz/swLvoHKwnNTwLGRipFM0uDbXb65G65XLqeca5IvBMUc1AO9gsnXcLf
es0ClH9TQCp4QKdb0H4O7qAGyicO9VwB4D2qU/BLJy58l7uOmRudiDlUgPW9OSXZ0dsg7pfswpzp
vm8O6jTWOHRdjWoLKagXm/4p0etM+sAZn5ChWvQBYc3Xy7xQIqN3ii9QgUK/cpXqqCvGZYpLn3WG
pAgTe/PhZtwERksdg32C3eH03tf3shC7F+3glf/HuJqnI1mDXtzVhuRMZW0+FHWZ6+rZGxj5nEm6
npENDcsx3y4cjom7PLYPGyrrZ9b0dJUHKCC454IrVqCFaZfPX0xKcc9KOvFXxc2Z7NFlXXj3KLo7
UMosB/PWdBQI7XNAiIfNWHX+mHpkGuW9VCAlfH2fz5P5EKvXdnMr1mIcTm6ZF7v2RbDylPr/Jjpj
5EBqnZeak0EDdmtqmaY/XR6LB6pBPPeUMu7AYpC2uqRE4pH0sjPsHC993vBqym6Zv1ME3znyQTL5
q+I0zzx8NBTmTCnKj1qFbacyisSLf6OBgZ6SFsZTm+3yQUwiXZ54tJVmxj7SK4Ic1hjszq7O+Pg7
EWWKb9ISaEasToLjY57XQLSYD6P9akK7I/pBjoqtWv30YfYEmwuwVboV+/ycL4rYnpiWZG83o30e
mAy6ZE4SS5FWKxrk+BKm6utNDh/GaI7Std8ya4NbUsHmRr64gXLDHXCY1e0uahOBMgl1k/l+wXr3
stpQpjG8r17v2MtAulqvJmFVlVYpJrk91C6nwabrj8J14zZ/bAUCTN814n53jqDMt/0zx4WW2Z7p
D0mWi/rNDw7BKB7vuGR6V72UM3WTaNN4L+OxqoU6R04HtD0V34ohsedXJPipRDBU72jRhhtFr+nW
r8WprMJsVBG9tzYxKdKBk75uR8vf+Cpfln+jq4lpgZ2PLQlfTvyWh6MD3UmRGMLlKiVRnEJgWhhZ
hRJtshLJZRofRD/a7pg4JV02Qxkz2mSyXi2RFfAjRryh9RtMgGnOr8Y18DaZbHqOJl6ItShYyIW9
KV5DqEZGV0HG0Br6f1KJsz6BpFLvEom8uucnRd2NYbh0nFSEhPxG3Ft6JR9kWLn3PlMOBlRutj8y
uHbOvweUDd1S3t3hJqViVn5P+0VggqzP4X8yDP+3SbWrb1OrooKi317x7ECIad2s3c1ORVFW1sJH
WHzWLkRmtRHaRbO3s3d1oAtSDWgsVsny4johZFfrsTqzbomDewBV0hBhNoCwRMg/9/EcTgZjsbRP
JxD44lKS+BKM47PaTwL/zh3li/4nKTKpPDNyMVt7Z+8waifw3/Fl6FvzRMiUzxDxHPqtuAMr5SFA
WPimBcrsP4WEW2vaxEsJWjpLj4XKnvg6OwKc/108JCOgUVtr2fMlN+1skkiXp5fXFFEqUF1HLQ9s
7ZNdxNOu4pSgVntLOqSCIk8c1anp/9Cqvp9Mc8mIfRIUz21VAcwm5WLUiTw6/PBf7bxIUkuct4yk
AZ7bUYl8W9MoNYheWMIMazWv2XRtmPi1djLnyVmluEraIQNzRXwe3A897nfBxvDdvaz3EIDxE9lM
iMbnF2/5/If6F5zb8At0v/CS5G6PopdGAj0Qxz+n1SNu/FuvdSAxm1BnSCLZR9mKipiaR6ulJWTN
fzy+bzsnqll5YkvGUQegc2GECPLLOj40gniCEfArA4hE7zUwLCXCMeT+QXAoilmRiqynmZ89sQco
QJbqflAp83j+brlwLCffkOaNlxrhOKE6tN9VF36aKqf+381nB9W76fQ+FWkZPs1BEkQqZjuHEDbm
F8N3ZVMOxT3+rWomADeTe0XMUeWtVwtcs5fzj+REyOq6eJMI+zpqnV2YXr08C8A6xpyNVfKmy9Sl
jaFJzPUF3Xa5wE7vDIeUxhTc4pWR1jkAOvtm7wo014MDIMkrnqqcOLSexJ8UPc3xZQbNyz9M2yUh
ZkVZHP63VdcDXm7dr8OFniq7cdVzXXUeUwJw4XktdvJi8nBTdL9HtVMZ8xvzJKythh80XUI0c4rZ
MHRnf6u/OiHZHOW3XnuZniXHC9GZaJLKbEP/kOjcQMGzpb0D7zR8TW5FxQDX2ofA3vFTPn9q5AEz
HUCVnx379AJLuSNh2tKJ4zV60M6naUOkzsS/xRafDhi17e0acZx1a2R4qSBToE4QnETJMxmOv5I4
1HHgtB/1Yi9NfzeYvUpMz+4I2KTisBiJz3ig2hhk4ue1kZ72h4Z9jGlnc1YUYPympljPpJP5He4a
kYXWE1NroHw/Anhjf+4jhbwHUpXhY2+lvEWlILrYgKCdRb84v1xZywdM+JZffAJbeMBY95cJqPO8
zEp1c4x9L2FSPh5bwrIKoPGTOX6Jgwt3cJKepL+vSfziJKQJQuUEUE039OOqY139W//Dx0mk+sk8
fcbDMTeTus3dpXtQee5RCzrctWCYw4YpPUewxgiv78tw9r+1NvsGZ9VyawOgzpZj7qz9Zn6Zrrt5
TC8FnkuID0WkuHcZl7TF1vh+0Me1mE8VNCDTnRnPEtay9n1c6QdSnwqyy4YTTtjtMSsecc5szTw+
zuYM4VndldXLDj14SVbZ2A9CIirPr3sKDxe4WUnWeYCSHp3LE0xFdphCQLohMfN7mcP7V79q3vAR
aoNLbNdurVsr0fc0MlOM8OE692SXkVDe7PDdtc1hzlv/L9ydq1P2R9bhlqYZhA28GqVjTvzZJOiI
zFiO9EhwliBcnx1wQHEZrij0GDSwMkHHbGdFpGPW6ODmg2rhVXd17eqFi0W7xaH6q9UiP3xU7GEj
pLT7QrCPhGpLO+JEmeEVJ1JX17yX7D2endkd1c6jGsVcg33llPOiFiES3oh1i+4iKzLOjZKlvkT3
oYOYROog0s1k9NgS3DIgR5oIV1/NvMaJC/ZHM06Ln7gmuTAd03AFS+MkDybCbIWn7HOnVP8tH063
K2b1bJravE+x260Z/zoFPFnpL3TkWXzb5C4yARS0J2MXJdKxbIgqiOt23An9P8xhVHzVZB+dg3YU
5ao5Mwl5D0Q6l5F6sqR74SNI5pGeNI5hZCRNEK3zVRGZ6l+MB08gSz5Bkvwu9zkOTQ06haz7p5Vi
8l6cZ2zfl1+Cnxcd7/eRDF21ZbYrULxiwmwod6SHSgONGLPZJXWUeUZQQMPveAWfUAMT4kQ3cIKm
dGhy0xoUleGWnzpUbAlTN30yP7Te6T9h7A29R4yI4cdW/WUG200C2HYZ4eUjvrP9QDvm41qxQW0N
jMp1eJAIPHpjIfQFY+1njeeRwbHiFxqatODyXzfhKTXpm7KVwCRbHvxyk0BEtiOmTD3eeUv9tEuC
5Oa0D0I6FbP05RqMIQ1ZxcCNQlWIykx4nnTHrray8fX5nvRZ7+82eAAFIYH+HD7W+bHLogi/Wozd
Znog5BJ3EMQPPYd6WwFhDyewPl1DE0TXFTnkAF5LdoKKoY+IfWinxhf7mNNOQnK2bT96lAsh3Pwp
u9DGnKiPr/KQtTmdK9yZ+qF7/MfSZwrvWO+Ve68QmuIzNlyV+EwJpGSxInL7CwAckafa+HcjbTqN
mMuEjjq3rxTPPoYHL6ZfhcwQU55pkEyfVIHxkGu2QenZppLMeqvUP0W2hk14WfZTqaLYqmV3uUi9
PpQVsGIxsdOkNg8vlkC7L6woMqtn021toLROqZtgEhtL6/GcPVutZX2O+3bYg/5z/Eoad51ixfSD
DMHMqrXbLlHFYBKgp9TXZv91e8OZriAD/RZgxBW8pfTxPZIDbU5IuM1+i24k18UxdbycmbqWvk0z
/4D3GYsb/h0r6Y1hf/fgehCZcheRCUmYqTVBszK5LJrQ1bwUxVlFpF/GDFzYh7Y0Ym/2GOgA2Fu+
Sl6/pn9bpGID8R7vxBugQ4YtWRyDwtsxbUhvwP+A9E4J2Fv2AdaYi1r6J7fVDulsvIXLo7gs4+Xk
pTEnZxN7Az7EQNa6JuFmpcO+lN3OyJApOZXLOXKxNEfSzaKrvaIknwf8I2GI0G1L86igElq9Dyh2
Cl8Fv2EwG4RkPnC2rwuhHD7lPfz0qTRi8SFVbCc76s9iTuwWioDpyCIbaG4dJt5zU/NtqwX/gOOI
GsUeDJEGcfKS0ROVtUj991XWW5w+EcbiBCibSoGPfaKkwlrDG8FzpzOPWgZ8ieVk78ZBqFISVT/P
0snzqVMBh51silTNAs/DGHLBdpWSXqd0TLWSX5l2XFPfHPOnLtxDsMYL3wUirURe2KuAxatfGahb
dhCYGCnBdVuVSN6wQH8hvA36yHi7TXa8GkAJ7YUAcz9+gDSFZ1I5OToCwXplqCYBug9YV147vJti
v9LspOrNf8Nj1y33Wcqamy+i7NKgxLmzeFb0bI+Qz9T4oXHAsJi/yhh2tTwD3uxdx5RUV5k0UfR7
PnOXVqTEZ3GurtxiQQCNSe7XNOmpDqojrnNZ+10ONAwIp//KVFB8NezJVOppfnV0/q83wuis0NOf
tQV9dcQJ3JR1Z0mLNp2mj+5w8u/5bKr2wtwaPoeXlr1J2vDmb5pN2NqHW/bcW/hsad7sQQy+n7Zm
gdcMZh5kynJYEQDzKAotkuIhwssihXRc21MZ/XCf3c0kFEZpI0+ztxftz1ZAaCoFKKMTQnjCanXE
xceJVf+GHcu2ZK8h8DABK7mTAoA/LoOi9e5bAQ6bT26QvacWdJi4XiZXqXa2ZNqeRQwqI8xo70RP
ehYdiaJc9+GU8tHqOx0n+foKz/wzbmxFOXuQNmptGRZPXOrKcHtfwaFM4T0fI96n1wGGjGz7ab71
hk+ysnqehNw0gfbyd3F15Wz8EoSkWXCczZs7SgX3VbJUUamI2atwAGRTwXLZ3hOjdrIjO1Ti1rGv
GfLY0rt0eW9fWVqWykh92nCDule8/ajnfSlmKsZbd2YTlVMffDaqmke4UP+WqtgI61KivREnUY/J
V4AOziqI4m+g+q2ke2hSRzU/8wgYRiRcludb94ih3iwlU6yfzH3njX7PiIUUFeo55ac7+2K7xKbr
itQMHmPoMLkTOA4SMvJKPDZy/aKg7dVm9ULf5X54sTGdYUIWuVjujADsz1GAgWO469f5rHuvq0kQ
ptbD0VVnZwc88Yg+5a2Wy77EBc3a6g17/odU76RwhSpcUE3NvNOvvEiRtskUCxD0XOvTRFUwBGgV
VAdMTPD1d2Zy1GxGUXIoPYA+BCecFCwhdiZxadvrmo6xFjhXvZPZm6lCfTMcZ86Mt0E/U5L4rosr
njoEO6a29cFQojiyso5kffJbRCothhhLsBb345lnDSzR0edGg7uwh/izHRN6HV7f/HXV3YJU7BDU
Yyko9LjmxwfMXZ5MtMpwOEEMflRt2LoMKQNzZ3CRLsFTw8n2blQfxq4xnT0dQxos1QpSolDV1hBW
Uf81AwZwmOb3YFlgCxPxuLm0rtxM7C+JFMKkhXRLB8yv985Qn8ww/xPozhrYmQCAa1qo5sp3Tq1Z
JQzLdOv/XgiW6oX/x0CgBEKDfQw5Vac9AtnsXzUXkZmEi8crf645+izm3WJMPjfFWCg3kFnTryVa
88kZF5xZeAVTk8K3wuG6LZNCul4TiSRek4IC43q4jY6tWKlSkE1OXKVoK/f8vjnhIoIU37UQ9G8T
NBdm/Bh154U8KKsU8nom7S2J8FfHiOVO2YqOXdi9QA7Idul5S89ykX4mTF/R1kt41i2e9vxWgMnh
Onv+xcJVRQr7CYUwczp6J2lQwUVo9gGEchTk/KTAMFieFQPb90cgRI46FNKJ5oLLD5x5lsfie/+S
LZi0N6mt6En61sNzWnAfRNnWBbb14Xlum7aSrleniL8SOCDyorJhbpwwtryxIKTbmvxIgNDj1TU8
a0jbx2J+Tc8H76xDvfU3Jex50P/2CKFGxSx5oCQzgj8ku/fvAHDqL46vbj2AUoZReO7ZVPnJn9uD
lrgcRaDb4R0PfOQ0aGXiKVyb3QsBqays9nI84mV4QsuzIz1BfbS5qPHdYHP3Ob+yCi2bofRP6fYL
4iuV79QEHtW75CFCEcilp6ICNzxVQK2n+j0L2fukLFmh9VeeJgxpoeZYoPeHhves0miOKt7/ll1O
CPEHwbEQZQO9aVP4+LlYSMUSa932nuzwd+sD+IvF5ApKSFXiTVlc0IBp5aY8tD4KV/KM9C8cW/ON
hWJTuWT3t/+AmjFu0PYHZn/+XDGRyFO0nISalIQ/DybFQwtwthfD9TBS/tz7Vt3vknu8LAp3/dcc
O/2125RUT3jc5FtsMa0Xo8XYtuDOoGSFjtQchj+hT+R/6WnxWtw55vlQ8+4uZ0+rvg6p513Yt502
y7AFFuAQPm91QHw5SvvfhP6pbH2rGVwSNKEOzWTiPkC+R/xohMOPGNlMgb3b3bHY9Pk91Ga1Ow4X
f3rZFcCq920eBvw7Vj+hyzgJhMO42eVmH/QCUH4pCfR2binuuIMxjBZTqRgn+J7R8aRBTMhdAf+1
UNp+VxuqGHFPl72bQXSwvGVWPJI0FWi/DPpGFyk3lCAwlmh3PEsF0Zzb2zOfYerLkYfiBeH+MYnn
E3fiL1Azqxqa1zYaShGfgJTVi2LAcAVv0ezvl5LU8FHI2pdLChJ5eembQGXsTKlhwBYILFHUOVOW
hVLqElM/5YUVQASNjFnCzwH+nZHD6AADXM8lSbbY656T2CcoBOx6mcyiBzwg57MoqoZ4u8jxTiiz
OCr9Fra0hUTJoRVGsIo4ugn2J94/5FcjSnFdaXU7BnBqw9PJcj+wO0L52WDMJeyoSdkRct86O/pm
5Z+WlB/FUFA1yGz2F3vMBtkb5euwfr3RShKnwjLee51g+Bs9CdvhjYopyhWoYOOVJ4S6cSzNk27X
s5JyF1FEQf9QaSM25q5yDIH6Vih0K/KM3w7p91kapAAg15x/8rJUdZhwvFyIxsi0bzdRTmkd1yyV
471t240/fYHcGMMEE7ZOSF/vulIOETn0YUHbQT/k/IjNOUJ1fDXGzeU6qj24G+KvzgxIsCsL2XwS
63SUwcSam0ePDHM4Vjk2ynnDlZSGLP18RcxE7jbBXuIMT4N9DgOmz7ngtgj73ThYa5PKjOGdCcAn
QpaQP4A3GKjRu/UHUpAYCzEt//S0iLpQfJRA3fb04meFilJzfrAdEFzg9rqHgmCJItiZw9yw9FMR
XQPOjCAt5VxOSn1X5nwoIaGrjnVCjTEh4Gh7eqALpEXi6logaBssndesq+edAJy2wEaY9cQPQkVx
RgETr1/xProdguhhoYIGrt3YC7Hut2d8KeiBXUlAOlox7lqNMZLM3stx98Grul3SHkVNRl/M8HJ0
gK65S+foL22FEC5zptXJGBFFkLy2brg7UARpCOodT+zn6XHADpjn6x35t8FCNpCGM/H7phWpCGt8
r/01bGvRlJ/wR4IYL48o0eT37YuKgvN1WLtOzrLLF+4bq/wUKULSMMLrNc281trciTn0W44Y5B1N
SM0b8sLwgv04bHVbUnbn7UTD2jRFaQggIBOrT/NawkS4UQ4Ri7CuvXXSvFEKkuv3uymXi7GDGCWD
BVrDwEAo/PIjeyZOKmuFXw0Qpi7C92bc6eSGf0FoKAC65CV+6GTI6UGBCFTGaLmc8aeZY5u8l4gv
rpyOvb1sS5EC+OmVkpQgS8mBqQIZuJIQGDRU6r3v1v5ayRnF8fVqVuhQDxDrmYJOn7wsnX9ICqSk
vn4UBShuoZsXBDuxh70MBiWXV5X6qMfNasll++H9I1XmqayMJwRi8RHT5jQRpX2S158B1pr9AFim
B5mOph4DMDtKi6Oog31LX/bDA0xEY4TxqOYXulHWwM/FxmyIW/RkE8sJSwI5olwixw/ZaxHfCaAP
e9gChsNjvM1rjlvEZjdG8L1SNHU9d1JtNTSQuFxNkglwH/UTuwLzR72gZ1VmWSlrVqUJc2ctNPJf
wmej8DuaTiL6oebgoBE8YoNQo+PBeWkpA0kGQAwHp4wchsI7FfAA4VHVPIPeYzu0hS33GfRGH9uD
OjGC9TV2CCaGmICs1sXJtr8fGQn8StlMDJS8QgrlEAhAMZsD9zzZ59CG4W8KGIzbwD4KWCi1QI8B
bnSBvQsjwYkXnVpDGju6AhAVx6I9S94bnKDrqRFK1sKn+hRGjJnvonzuu2bOgV7lN8OueIdc0mmd
3wXviJH+Yoq/dgBe2zbmYpfvGC/3o14QPz2hvpOwclZ2s0E82FmRqdj9j5g7n8+7wuSceKe2NO/j
vlw7LJZ37HmOLhjmY5DdVEivx3P/5J95pPx+T3qHrMYKjRs2CwLJDl8PLWMcOD7p/nSkrjruRE+f
nDLprqiP1lPY6SG7TdekSCMIpuYRWnyjCN/7enoGGYc0ys4L5c+QVbSxi79xniKCm+H7S7fctjaz
khQoZY5glWukOYX4EdwPzPjU9p5dY5zl5RYYFjvqDS4oAvWOkYwUvsYIEOjHe7pA3jFf8S1P6EEj
T8+6NfxRkcm1lbtWj6AEgaZihChUPa8M6PWGt3J2K9MUXhNrMeRzUBAbeUgMVnz8WJ9Ry1WFnN1t
6toSZlYYH5fWtg53CZI/7tke+yft7bP4PLeYrWdOY5FRkAPA/obEsm214EhrmD+fayIrkuH/a45P
KAp1PXIYTNeq3TNzIh8sQgwWeNoed6GtcPUwepeSWiXHasBcWa9LKqxfr2gYKp2SkDzBAp7enfYD
AdOuwAcChd/BAHgSWgd5FEkeYXyOv+mOi0bjOdKQPpg0naSljfZPHLzRxvGrqKlnBPeSN0WVv4yV
TwGHtWiHmO6H5NkXuTSRfBqPMrXjha+3MBvYXNWJxioaDf6Rb6wRCzzPMXHL/3XJ2lDtEoDqGD/Q
EQGECq+AV063x81zrmTJKs8gpT0zLvIqPLrNKnMw0egIZtUFbZehnvgT7XSaRvzlWmGw7hkB38/r
SQ+bIzIZSP1/c6IMwBQDu2GJkIxwI+9lH6/yvgoK9neT65rXabq0fa7QAhcUmWNcpa1dnrZ/yQ7v
BV71qpTzIvY5Zbt/I99iwZrrE1hfnU3+are362Lg1HvsKQ9nnbdQkEusYBSF6+V0HHCnOaKA6Sew
2C1JRpLho3odv2RuAjWT9IAmpDrHDsfCkHtIkx0oUpcG1cBnDGgLUM5kcyDMFFFUBdGcHG7lG8Tv
c/hjg3YPw6MKB4iNphB/0XzhYI8N/AxDRgUibAxqHX9p09BWS5UHkJFDD+WHkE954xo8t/HB9P/L
mdQjrnDgcBMFWnmwqg/FMjD2fK+WVv1ocUpeKRz/n/w8jRBXqZAyYklNs5aC+GcSZNSCz4v1lCLm
rrjW6baRreBNm6LHLmo2xFYQmb0r1GctSpoAyb/zX1Z7zefdFruodnDE7Lkp/ih1axazHHh3QsOz
nkM2ZRFCX9LJRbe39guF+nmIURrNfZ+MGALIyz0NY7J0we2GJr2NR7GirhPqLhldWiBrmovskOij
+Nnf/CqvWPeucP9xl3fzl8yAt5w/1NykSYHjwoqi0H2XNh1pE+kCYMgrJkbfWLqrluCmvyljgutI
5P2xU7ztHWfKwT5SJBen/flbxjpMMbNXRul90T9Dak+ixrLh1rBlCJeDr8VxgBNfFjlV9/bKS9YV
jzc0aLwOccom28QU9l3zL0h6wK6IfAOZfwPTaFfaz+eSgR9DubNhrFkT3uwklzPlKyhf/mPvZu61
EvKJPApai00zVXJgHQ1Qn0aXVW8bYf2fh7cTSNRWmF5pfWct0J22b1t+LPJE3+943yAv0wQLmu9Y
ke81m3R88EMUPPQkEb3S5tLz2YmSwxQy4/v8pd1tzKpUEkKl6uJCgt5TjkmwFtEJ91yE8NYtN/Fu
TTYP3MzxGd+EKwpU91JemjFs3bWrM3ocC6ORquCKCrjlxjfhL1FxCaB9pBW3tOyKak4DwE/Df12b
hdfex2husQ65K8tSxg0ubM2Xuc7v3Ol50eLauqDkR4sFl2TlcaQ5k5On9B+b2NfFrEoVLwUC4+s5
mj023q6yA2MUCvFc7lz8VGE1DmjabjnFzgukMFrYyQVeM7ZEZPm/L57qVtxCocmB1F5IiNYmgOq7
TaUS8E9oVpgFnF7EI/U0pDW3Egdjdw79nf/yOrfHHAabtKxU+QcvK4102YUchip6RUgo7xp1Jk9X
HKEy1JkuLpZY3NSz/Se9WkeDVyOGiNh1ojRoasIqhcj4qjtCEjse9fZOn+0NDK0jiOqw65F6jmgg
Pfiel72ZjZGvmDggv0kcz/pVZlqsca/MDyIE7fFOCjnx64PJJezxtTbQg9KKnXgXTLZTGXB+wwlR
apaX09+nTRHyZiQ8VTQq8rvwlhCFND5AFvfmUSq7maJE6btFJW/Ec3qO94y+8XZeTJ4s3uvkx5Eu
mNelsIYMZrUykzi6D49oKrRglGfr6V+uhFp8O2kaiofOtbZXHyZBs0IKwFKTPIk5p4dP3iQ7h++P
20e0NQo2PUoDjnN3nIZ81L33m3gGP57SL9UgSIbvCvrOjG8NeJcvnwZdOo8Lny+QTPMHjO/M5OCr
qYEDayCBttEanJJfsTpfc0ETQnVssvnw2gEqC913eKiYh/pOFQM6Eqi62zDkPC5YjtjOndaNTYmz
hV4LHN70Y5oNUTgvefST0lv6eyhx710GOC/q/tr3UOpDVMxpNXdMKSXNg8FzqYbf+zbnqtrCzkOu
V0RCi9+eXDH9A091Wt+vNorHTosqXZZwMojmtEp5tXMyl5bU26DCI4A0sTEMoNDbYq+IseUIXDzo
hEVdt6aSw0gxGlZVdbljED0vQaM37+z1zJZve2JauwFUbPAw/h3X+X5gCQ7p/R3Eh6QV0mk17/+a
miHPtbhpYYTDI+uAT+ODbE/wmbwQJpAsNqA0kvMKZ9EmdEhyhEEfWeq7vBKBfOnISqnUPtGxrR1i
7+AkpRt0qBaIlF80/1IGJ17UUstN2yoKjfJUxOG/jo6i9BiXvUd0NFz6wR/uRjJ6tb7hw6hcxtAZ
E4ee/eWuDlpeYvj1SlLCuc5IWKk4gS7faAfFUBmVFkP+5jnf9VCYFajaIU2SX6y/kOaG29/A8JrR
5dV0nLyVe7aoMo+/u0dWxk07mg/VYTXIzTQUrLNZ5v7aHyOA26UodB/DJa3OjR2LFa0XbLaOr30F
E8DOUEPHgmD+DlhsrfhLhS11ZAzturU1SVrQOVXCM3mjoFfWIeZUSudPhywcb2b4ZNX/A+476vK+
cz8yQAOaay3pWNmCNLcanBG8QOwQfjssycXbHwgRmt9dESlUBTdsdkl8MhQ8QxXKLvwNYavMjVjB
HibYZb9GGK8X92bgjH6I6FIRvGGMCZK6XBkvRyepx+sOiRH5ua+sDwx0sVM8SvzTcMGmiZRFxwCQ
k/az/l9jAxuJdkGqm9luCGaQ18mElWUZYpZSPhAXG4J/SlhfeHa8j5zx4KYNVczKMzxPIV/C59Yy
E0oIzI9XlfYot5HrY87Q0dT1Jkj2NmMDZV6iSqkjPwLsCmo0R8OydB0Dv6z7J87zSBFiTQ1jjwax
EATzMqR4GTdSh+y/Mxgxz0Q2L+lTvO029ORpi0B9p0s4Zg6y8ISdDciWsCm2fKyQw45+bK0lI6l6
M1oG4Lt3VaoJdW/vxajVhbFz34JapzIwVRvTcE9UaUKSSoHpVui3rqdlTeJ0waT+C5IYOVnDyApI
6ot6vF9xoB500ohXY2LwYtkBnCZUttoDvpb9pvLAgbzARVe3o9Quhv8F9TFD8PzsMewK3Gco+dzE
8ZS3gjLmW9GgKlJeelFOqiBvdHpohipA/fwv43cq/EJ79EOhCusxFTtUW8MZl/ZssE7entrP/ZCB
Qqw340fzEynAEn2KyTbozIAoQvQrxJKsVxvz2DHatgKBgAx2iArFNVmIegfjXmevV2onlFMv4X0E
Hr/HqbjGUcow+igzHKSIDnd5V6jpwfokKYaWbjfAFuOjIHhscfSf8I8seIltPNhH8LwNw54YlUVO
u/HPupFAm9bPDsQuGJ+ZP34GFXvG0XmfuP5Bf7leV3R6fKWuSYrKOLa5BDXnIoB49sTJeb8/e0/2
T21/U2paPOlaZRNikD6TdXCjyrIqiCQs1geSD5ciJ4ouzUX2zJJR7VG9Gak848TF35yMPe5Tgk2J
46Js7KKaiEKWAPiyk1TZGOY+CjN1peba+BYXsnZVajxYZke2UxcI6xJ0C2nU/cgmZSLcLBRWURhp
WkT/dTVWfjYAYz6pWnvAn6rdhOupi2suRgn8rLC10aSiB6d4jmwtIAW/kls9j8G5Vzdpro+ApItz
H2Qme5wvHcMkEU0M2TlUBF0Fn+HMMvt/TzNanQjPfFntAC2AXkT5x0GPQfPHV6pHPqAAYPkOooKj
JAF15RQduwEFScWcoBSwThZs4rGC0taVz3JhJhRjh8Yh6Dqvj/7r1gp8XQBa3AeyB++1Qs2bhRnA
qWkJL+X2Naxh8LtBpqM4xxFD7ToyNJ21tmxncOUlDIb8kJVDuVhpizn48bQ+ZYHCCqSl8SdPyr5i
ffQPfiuu+8SOwAEBkm9VHFfLSvbAPIXUgPbzlZy57kghI7cIijiw63xd4j7aiTevKrQ4+qZ+zj8F
LBYOLp5U+EN+hQ7RUO++F70o6HD8caSNKcPcOoqJA72cv4sCrTO9IzWTPV5AMtfmrumutQhfqNC+
SFLdO24hu0b4VNbGz82Nq6pbB4AWeSkm2syxi6oDhEtiKxh6t9wv5xsyRbkDTYqjRNiCUrBQeQA6
gcGj52ywSt1SmFZg6LmbpQypuau/IKZuRNTMGupqyMp7SmuVUlmFwQZaNYRbECtqkJXhd5+7O8V9
XBDmm9lYQIN09iAwtUWVARwfdpdcOR9vccHnkYSYc2F6NlMxxqHYygAgyaDkRRzvN4nTRnYeb0/8
GAUejAOZEo/BDogIC0EKmGZDUEC0Uir0YAajZ8ZN9qH+KNGO/NKwSj6CCSSSgn1DjtXsUf3LlRFi
gRAtXRRjnPBWd9xzwxiNPLt5yCFhBvXHqp412Y3Zrcsre4mRz//xUf5V90ZGhL7++G0xmlefN8bp
YAUpxPCe2zDX/TGzGajCO4qkytK0Inghgxvpsi/KHCR4r5E9UzmXgZc+QBZdQ3rdkNQm0gMRVvTf
PLZVTkz1jNEwDCwGYADa9Kub1UVWv6O1wFeT7dsrZtag1sLj/+bqs7hI1LAUPYFmQ+RqNu3E30uR
VgQAHP5jc8f/ptYt++mAkgPg9O5sEPJDimogBedW4NJJq76bcduotrkbOdS0rDK5bmZFQoUREZTd
xY7Urz0mGw8YU+lkj1nKSV7PppIHpKFMFlUu6tWmT6O5AhD40AmpOCwA6kuSWKxE0O+AQQtjBsNg
J8Uczu7CnYkyVne2laE5TVzAuXRepv1fO9L/8e9XmZ6YIqKZttG8jkzO1/CV9Pr/Ck+5a0WEDY2D
dMsribeZl0fKLlimHcG2f7KmmiOWA8XZmULX3z63EtwuLNEbx0czm521Gh/Vmd404SIH6/9mdhOt
7J91tG/Rszukp6o1QfxB71Qnu4kze+NKhZVkdt/TOFxpqxvHFQgIF+zAH5o4+vs2Y95PiDUiIi0G
GwAJGWpmudBQ8+MYHIHzhvmePXMtpSns9P2VOdb8esU30lY+VzW2TweZOGq9FeGf1Cz125FAAQhX
fcT2SKjx/zSNw+HeymYomh8U11oCiFSfkOTAsggp7roUmOp+7ZXO3N+ZPVA+LIXVe8z8IkeJlBHv
eq8YtBHCHTNQEcu9a13QXgi2dH5+g6u1pwQcNw0oKxgEaLGDFWazmp1LPwhK3iw90yYt0tzGroSY
mRXsfqeXuBfo+1qarAm/4U5tqj60h+olu5odwADDpVBj07W11OK5rvqVeJa/ccTNHCh2KOizB0lU
2GQeHh54BFxZFZ9UApwp+hLu6Vq8ECOw4yexdVB2I9hq1zDNU/ev3OFdluwT61EWpH7iO+0Onwvz
RoDthd8mcS6mBc6/rTChOJ1/mhT355RK95KdaCrbhIEYkdk8yZiFcudUmcwrnxOrPxEasU+CfqRk
9YciCzT7n3AwqvXWC5FZ8y32/Znjvo+d1QBuX5vF2m3z8ZJB96lzoqq2cVM1Y3N9nVMh0yfLeUUu
YZqTKCquncbIDohBOR4oC6i332x9R1o4bI25BhRRuzHq5hLvgnFjoMFrqwjoPjAimq/VAb4Ffp3/
D6xvz6M7HS729XmsFr2mfu8vTgToJE5O9Huj9JVgvwg4Yh9pr3alkarEmGo4rJt2zlYcXDDwChem
zax0lIYLkuEcRRVwCxaGvS31PRGfaHRHhEPeJpUo/MKW6q8qoctOj7kzWzJBinNNwr9Aafi7m/4X
g4crtWnMT06QSM30jO76AgDMvgKUWmOqunrJNr5ryzcZKt847V7xz+81bnLlYs1TE1PNOmAaPQL/
KSD5tRnabKksi8O4zaJEvx2of3XdL4LNHLK8dgdTtHlzIFKmqSv0mi+orAgdR1xNAV3INj8c6QHB
zWo0VyoNKfS02nf81gaLN1v5iIN7wLgStPmX+Nfhe0DUeS2v/gT3HByrz481VtMZGmrW4hhQMpV0
WOISoKaDuxrQ+2r0obUQ72JibZlZPq0a/sECa753lqWjuewyEI/Ze561KHI+snpkZeM0GtEVo7NN
kxPMBh7o3hvj+C3bELdwY64KInPqDPQ4cMu8bhgaE13mVHcnYI1/eUulYq8yM9bZfjYt9QRCxVFt
YSTyYnHdKxG+Y2+f92AppNUp1+g+4SueLHnfYgrHw65PbR0l2lhYPPDKxQ0u9YwYjd1cvJBVoLXg
wQPZhTXHMnEtUHjcqszB2I2Zn4PcC0cDFrxRKsF+8MnB/G2vYCko1lPb8Y7xNZJ01WdiAsxvOFAd
K0BLbEk/W69jce0JgmO52QqTrDZLdsyG7kD8fbSz/AGZPVlWR4ECsDTfNfhYp+KCuj1/yLiMdaWh
NQE2gyczO/YZs3UZEbAT8e/fVdYOjgnMSr0/KGDlcmExSlC6eXoIwf3n6azPbO1MRUqeSDCiwS3E
zaSxSLu7y+MV0m+Ii85e5PYbie6PjB5cyxbxFEnqM/Y4txYs7hGaguC3S0ODYXUPC5QFmsbpu70N
djKLCr7uxAtl/FXHjr1f8uYhj85DY1/DGIGuBW7vw5oGLl0RIQKpujOVt9qFkwwdBsgH4cwVgbhN
Tf1SLl04FJnse8+ZaQPqPv5ooirlUdQI7+whuNONYKfQADWAw95vCbce1svOwX6Adn20iK5hvdCf
pBubOnarklFnt9naFLCWj4bYdtZDGg4fdtNnUhHj0yNijXBsdK2+5n3tdx7+VecpvSPKYrmnRMF+
8YZNsuWLF8ss+2qIcGJ/c9HuCIyGAy7tDjbJQGM+ySZqKjsY1Ihon7uKjxriPPpSsKsjGWK7G+Yw
WhbAStRxwf7L5klBKKlMWB7oZTsTyO3iWfhJKtU9fAOq2mZGkVYgNEzxCLmtFBGRlTZaTMORktGZ
hufZ4wJFzTCTqYzhW280CMkyt2aLpFXWdxWm2qqa+5aWyp3IQvTgaUEXky9jERL5noenKdE650F9
Cgg99jbv2g0J+bjzVl+qP3LbaNGW2Ewn7xpfbvIhDPMEMtH9DKX7/P08Z2nd5Hok2g+uU1cyUd/b
66m1fmh7dO3IAktPZ15IuG/WScPRP8O7Imt9kh4hTp+ni3r0mqxYv/EpyNc7quJi2N/KNTd/ODWE
MmKhoHLwuWVDhIhqHp2HgSujaIKIitM+pfIH3tv/p5kO4knKDKO2Md0/jT94VG6fBsrCRm513La1
zNfkB5Z2JaAnfBp5bBgOe+JO9TjBPP2ODxIWlL9MA0BeZO7JY0FTNri05fSD01CLbT1o3hRDmj3Y
KX27BcCfbukj3DFQQ5ZWSJfvjkp7pMdNG6kjLzOgU8hzoA/cH/f+IKhGqKlRoUNW+6fQ5cbZYdy1
ieJ6rupAtONYlEzcnpkYx4DA4W9QTl2k42s05hFEQQTbkpJ4bWj74D+JguFKpNAasLmHnash0mXm
hyI2uGqeKRJreNJB7nWnrGjI0ApFjd6DuoLYL2H08rvC0aV1golPEQsIlxyKGVFAq3pWICFbQfbU
6XpTd6zBtBe8r6yZ1MRmXClRQwwOM/eSYI4ExpKEP0vv18FhZ8oXOrCnxIvlWPFd/iux/CtSPMO4
svXxaxQZNyhVzILkOFJpQzSFikWlwSRZV2jk19Un6qxD08ngxVLmDXwyKTpAAVcEwXknQAnEsg+L
DI242CvJaOGmWZIKYCvJvy4W0wvnTOAVGdUyPc6sBvwDV6EOpqT750BZZ3GZIIyr5tFEGCa7kqPL
+ydrB0OpBKGNvaEQp9uayGhBeOS6baY8RGvLP2tAfgj4W+FgpVEmuftujGluJd7DKEBHIRY5TnQG
J+YA0cUKaeCJc8RwYWIPhnDpd0dSKcx/UhgHHtccg1k3nRYu0kbqKA8IKcHyhH0P5YMGbTAr9slz
uzJSJvZb4eeM7EiNfMHn4KVM9dNAdEHJ4y/NjwjS8F7OQypkpKHlGkGGtUSIwFP8OM550zM1PluE
AiLdJEpokOP6Y2RmIbdNVxqpO182UFGfJ1Sd2t+YdFsD+dLBxfqJ4hHjw77A3eQ1CbrE2N+r9ZDk
2VKLOLzlkkmrEu9jxN5gPR3nHEtrr6FdV+7GSKENUGlf8c4dN5dyuIsE8vWVQeXvn6k0khfnag2K
db6htQvT7VwALJyV9ByRLoS12apD8dLHd6OUicRN5apmdKY6FYQ0qDlxaCvxvkLNubVNnQEIpIGw
vRCeT0DROZx0Zq8vRpxo/2VLd3cTbZqPHIPEcL4epON35CTqs+IoRe6LL+b6s5ToRuK/GQc5s+oX
MHF/CAmEIpC7bUJkN5q1Oh1rPKRxdTCBZOkVsgsRvQv9dKx96K9ZXsKRzci0+9MNLOoEuSxr/nrk
/TjF7Vy4zhdhW0XhbTapYslQ7nBSc61NYx0GzEANqTH/uBrhE94YxKBTr+TTbCVqNyKzFuYeWuUv
5ESQ3YPg38StlcA118+RoVWbxOaValNbG70zXT8clpdxV9PitP5OLg/H6yigeqehfdsS+SU9zEtz
SG5exv5KBqK/+zxMD3Ofocyf1tckuMvDIrvzF4cZZ0rmILlaRmBk180NaupXbs3i12nY0Qv0Vd8c
2+kNJwwwOTXnP9ogE/opNhIEPOdikLtO3sDiXgKojh+44XDhRRVVogQq24XAlhJpPwNNQaALjLw4
0OuHd1wyNpCXP6s+7QMfmKESG/8f2D/uVAHAglMcaqtjMP0z110VqzWegkNyjmM5diTqJsCHoHfG
Yi+DaG6lS39S9HKwT9ut4ezVlxHXiO8R0P7lUG4fw2zRZ2bIle+XgSylU0yWI/Zj+OmFuAfySVzR
oZH/oXKJbzORtL1EX0+39O3prQDhT5ABetzsMOtL47N56ob4RAvWc8hIyoQu9SGqTl7Aq3MRL1p1
sS4j00lxxMyc6KxXi+TxyFAWaPjzopTGPLZypplMUV0/nPclMRpLUO+s7IRipUln9uiQHwbe8iEf
KEPJBOElwqKG/fO40Fc66L/dKNOSqW90FjoZI6kCyszo+rBceH/slKhd2pnPvIL552kNRVWE0Mpm
uCuvGwgnalheFZSSj2kLpcRpmmbufA7NbyzDVnYjA2QVjOjD5d+HX/+LGnn87WqjTH8V4xArg/Lm
BLSHLOUkvvC1btTBuLxFJ9KehtF/yxZZSlxs6rnBn0AGtrK08JWV7n2pgCr+4syV0D6N44/S8ak0
QF6Tu8baTdTXKgsCMYNEceyxYuATctmQy4MaDNnR8Y1UDmrM15MMRxAf3j9kT7q2hCnUjiq/V9LE
IvcFkn2Pch4QLbOsrf86687zTIYYr6EWX03QQ5BO5/PCVfT2t7agdPH8pgisS5b3m/1+dMjJrAxF
hyvjRwkGAee/P0MQP2QnNO3sqbtVDbiOWVZmmktyPaHD+vsVOU3mCUbMCfO03ZgJ6nUdPhaZ+nww
V3jdkRgea44fUkwBGwzfqUWyKc/U3Dz35ciDZwKOn0vBBbzLI298iEBTBFcPX7DMbI8Vvtt8JUCT
CIEPhE/uKCQqJWgY3wB7hW2EUpB79ztU2QgxwAzdC7BblxbwJQ5CAFTybxZiZFdh22dz7TD6egd7
Cbka8gF8YaLQNK8ON8LO5dzZ1QndXA57sUC5VF1AJ/SOE0DN7K8Yjilwa2REZZYh4STrisga5o5Z
YuQ31+13ooTGRcqmGfIvaa/EB/zyrCxJw+I1/GMXsiVunRA5nq5MOUhvudNn0BOo6r776i8ZBI62
9X0oMmeKBpSalfXbxZ/iaxFiTYjQcIdcEYujqhbdt+ifeW1CwewPMQ6KXlIAjDCc1yP6p/Yst9T/
mqPTyhejVQWb8+QMO9yT7gaHO4VxMbXgbmRnLGOwx51XsuDsddFXnJ+Gdg1r51TdPk14ZLCLzSZC
7N4KelOwKqoNzAFx0Gmu1Lw9bsITQS06wGk4mdKXImgql125PvXS/h1Dm+pg+u/6bGrtMfl+uQe6
8ddjs6EoZjG1WzdavnK4Tg3Uuza1+G+qckFYW7ASomUjHTkTbCwg/Cu1lEqdmJDkUKhIwikMUdQt
U8rsGfq3CLEHsR3qz+6St1Er4o8jzlXr2gYfMtTV/iES3SJYW01O/MCJO6xOmm27MsPBeWZZMlvq
1RnpXtV195IemY9zoGC/ACU0tJpcFD+gYtWFG8yAzzdtTQ9dl2rPlGG4KuyApGEOixf/p4DNpzxQ
GekgZ/kX9RAt1O+Trj0LYfstWmuvXjXaTyuQJCfsutC+RfwnS8pODRuE1ViPR1YcU/YVv45a750n
zYLV5W0su5aBnUjBZyEoT9n98fZPnv1qlWhTKKfeyNaLaVyWDDiPk5oRSvp6walmD+5CRD+4X7re
hPZbDCx8nyDe31SSlVPt149ese8sYZ6lpoyxgA1Ym3A7htOdduk6ehjKp89POvibqXi4I2bFc08q
lU17MxRGwTpbz8fPfzHYpnfMR8UQP4Y59G0E13vuaYPN9beQ6AKoKc+RhiXASt8YRQsISRW+EnKx
svit+mcZZgtYe8hlVYiUpCfv6Ma1xCAvi4lB95eRIvrnLQyv3qNGpuJicncN8yeih1Bt6xL56QLp
nZIwcFsAyYNj3dvMaaBYlakN5APseTLqvcoswBCk2+hH4KpqMUgZdVCEgGbEGUELS7e7rcmdRs+s
tbOf2pKwYL7wAtjeS9HR5vKgKRC/q/6O92Oc+9jCNPUdlg/h7xw/tfHeZm2V7M5TXajfXU7hXO3o
qilVlyhjoM6RmrFb0Qj4tV28FPQbklnbyHkxp/of7oG74TBafvC7YNYGsP/I9rw76lSsKe6htbUc
z0pNAvHXW43j8skGa1Da3F71DDkgUGDXkQhEihspxhrI4EOGVJ5zCmqc+LqNHG/rGiOpD5LFBAEo
qY331bz8tpM8f9PP+RiYYbgwBq8Quc0ML1MNtLmzpN1TyqpFzsXqWIhHFihzK/byOSAWKlA2Z7Mc
ZIF15rc4EGbqrqBzK+o4GPLvx7Z7bW8WSdkHbsEwev7Zw6040i2I6U4Z8dZgoAUkUUMZGjYUImiN
02bOPDaCi5x6SZSq0V2EBdiAja5tZ/Sko79TK/icVFlbV/Kf42T9M05JsDTtzXNKBrbIbCUEAXp7
YWhLS5eRdR3wxqwOUIny8jZa/xd0okCq91fex464KgFwdPKF19jw49pf2eRsfhAApBtF4AkrhOfO
EWeeOF1IKDq+Um9iHtREdzxS+YJD5QfogjWpLM3v/rko/fR4SU9LOyqkP1OR2CwW6MOpJzjX0ZUa
5ldearx1Cz6C6dHWaZCNLFyKnbWz4LTMr48ofsA/f9Chep+OKGhq0BDYpiPQt51QTmexDBpG4Qq4
C+Sm1gaDDobmbcuK11HgAU4PfxRxhp8yWGSwKj2lkGX7tzVAtjraqgFvWzmR2YCTp3yk1l4qSjxT
u8AfQdRJJuHVQ3CDHQLWEKdEs0bzCUEMM89vkfYhPuNKqj3CsatOFjnpkxHiy43B0XJTzMgW5Pex
ZSbi0/akuzSMhmjWNVfT8OtNTXuONHXRMw/1YJjcQ9VAY+ms7HMUX7D7l8zAGs7FadTwdRaHecKH
rjDrmnFlyg3FAzFOqBpAr8i90SDAVy5VHwrT3Z8Lcu0nB6lQxoXeDlkGl9C0596eWg+N4415VBu6
qhWDidGNLSQvsXbN5ofPETYlbn85Pod37d0AdHZ+P/G5jGWE8SXpaaj3nzgEGSKutqpiYjR2bjyU
YQwwWb3QRsVK1rdLm8y64j16ELc10oMLDQieoPdsExbtGCdSjsRs1ufmSbUCxUUpd3EF3raMU363
HY/7FfloENFSC9mr0cYuWe/ez7Xe7+9fi6+3aV+1Cwzuou14yUmwgfJWt6SAjCnH1sjmlJHW8+Jk
HPKmDDLSpnSpKUXIQH/SFlRRfQMK+tlhDcjMWxo7WSWleCXqLZ6ypQaJuOGfYz5eYBd/kNreRFSl
34oxOmu78Xwkfk6ENrDwLDcRJfoC6pq5qpV+SlUhyaNWPIguxifBFBkLb7uqodDm1/U+5zGOHiyl
7OtHjhSJ+fxaIXLe50UO5qkFLFOUMcwU0uXgpMgzQ/PViRMLtc8sYHBLl8pPjqtWdMogBx3A3W9w
Qgl5jk2JHcYeS4DFdw+7GK/Zm9XY/N8TNTIskOUJp5PIM9AI2/P4CfqD8+RbbCuG7C/j69xvuhy0
QIot+ibKI/J8zYxOpHogJ6JLXOqYiJj8EjenJRQc1FPAfWbOmnVQHsXY51US3tkFPgP+dIoLuLv3
TzAHw9S2zLgdiBNdMrUkVmfBxOTYz/gGFO3lQGTgScohq9d89GcUg5bW+XyBBAFxrtXuGSD4PHVS
AFaTBn9WB5NStU5uSlYKOaMiNTsbUVOhIUxTQrxqO/PqWG1gzmJSxa+guJs8/oidCJT/W3TZerS7
EwGchCSGjLrOSytUVCNdRCnB/S6fk/p8cnSd+IYG9rD2uEzTZ/xFpJcAmtQM1ylognSwPE3eFm12
Rf4ZvOyWafYjuzAAUwoGS1GGvKjqnDxahI5VxwhFjIQmm1CcOvYjQGZsF20AkwMg8d9+YBJRblz0
CMHrQS2V++qzfDiNyLz2wVsPWKe8cQe/yZBnpDWsTxiZTr+gHCvKohGKFfMs5zP7OzslerWrEx7d
gNsC+MT3A48lTHkrJ6yzd6/9CrbBJQbCrw1TB8vrsPdvOwaMB6HmAYH+zEnZI/o0dWtktMac/5Om
CUAq/YVY0w7CexHFZmZuMR+F4LRYYg1mFQ9f8Og7de320pRAmybAzUmTziBaHYdfLlCcqI+FAOTo
A5h3VRudrf5E7wvDJyJ4yh2We9wwEhdEULCxCo1Yb8GNUGn4If6/OMToUEFJJ3PSYerkmpJhuC5Y
JH5m6S5Lc8VqizYaPiFyRc8OiC2sEK8a4niTYiJL6APSzoyBm1sc+GVbLYZQxVdW2+hE3s22e+PL
xSypSsIMV/62jkHtYyeThJuwRQ8nH7LFCcmRiwZrfhumEod80LCueI3FgQeRGTOUx8gfuNd38dny
CSjdrUywsrdmtK7yT4Sxu/dQi60cMkQAJBGFUfepBnNQ4YacHsjR+GflVshthkJVASdtQ0jcJH7L
6JBPaJexu6FbLFm6ORvCStX1JMFuR5ilUnz8hUdTmTD9wxi5WMPVIEjVAqVvAVCWXoBdsMZNUoHf
WZmPn3zGfrf797a/QYdLcUq5hsmbYTYmU7ikVu2bNMBbh7Etw8FGacNbTJ5cH4khBF+26pWD7Owk
QIIWvXjeKpWgNlYT3l/rt0eUbnIK7K91L64a26gKwGkRj+ot5pQgesT7eN+/RDtOIXxtGcWTrsRb
v3z1j0aFmVBiZw8BJN9FxINgTzd/+e7YH++9tbrYCF6Hh6y6e2CfTlGRXXg9ej6oiQKr9C6p7QBt
xrjBcFpkllPtGFG6e+kx0NvJAX0WqhijXL0KSaMflSzE8k7nMxR6EW7oqVgnJ8HnT/2XlXyZP8X2
CoP4gI+9fZ/EcYJU1kQiOH7bhVkz3g06ZyVQ1/aQDWpcnwiJ/TSFgKX0EQuIG6VWq68iuQDDdLu+
1cunfx8k8/WTZa3Hlh/poyvsoAJnn6ahDk3mkx6X6aCQut3FLrcnayDMuNSHJ4IP0MRXZxZ5Ai3R
WYNeLmcy2pYxCLL3fIIp/4l2cKuNdJVjavFjpNe/JdhA+uB5VqsI5bmh9oYhb5bEfNkus3u7rtB5
pWCvfKdc33dVijARNV4k0kyLXoGVP4yWBZe0ZKJgye+6mDarr4KIpHA19SpbvvIRQ2vjzmTsVxZ7
O1XxWI8SP7tko2oTHLVtGXfLl0j4zG5ew+cF4bV8cthTexDpTZ+zy2jh9TcqCpiT4UXvSZ4Vpur1
hri5MMot23MGnu+1kBWzmM/IPNYsEJpQVJOLq8UHm3ciMn3oboIkm2g4DPly3mZ4jOBMiKwYOyQY
wxZ7ar4ttc8vjhUwFPjmtdjJdksjkd/6rBsp8cAlSZO9AdIPhFA707XOGP6VKD57Akc/DCncMlEt
WduIvE50RSWJ6qMCdOGARmITJPyrMr7hzYpQKY9f1nh2juuK9j20neaIJjvIxUupDTWVn2GYxMyI
L6Qzm/x5WtCKkl05IR3deUVICO8P9YzvZE+paxISbzgnJcz51l41ZlpdfDRshTB0fSOE9CR2YeOe
Uv6dYuayxi8oMj2Kzp7cWC0fC9u1h1B8K3eiyc8O2z7M2OWvkzsxGxUdoallhggCFu1fLAPXs33U
ygRovJQ2wsUZjY95EXUYV7ooSoJftqkuAIhubLv7zJQQQKoBcZksQY2TFoIWOzin9xiwJ3kYxPxS
iYPuvfOba7z+8NTwsqkhp/CdX/Newz0CAripcfPsNLccWXyFX3vviLVFXiJyLk3Yg8+xsLHtvi9a
c4Ti11BDgVDWTzFyGfDHdrxgVlcBDdQejXK+lG5XTgeqB+ZR4G1BOsHfR5pcfdIbcAovLphvFEvs
QEYli+uy4hoSaSXg0/fttIr4JF30AL8g2aezWg2Kd9VRZqlcjVDFpYHN+TxhNp1Hsoo5x/mFebSB
BR8fMIkR3Hn0/vFvUm3p8hXXSD5NM8W2lb7wr6r/dXgeTj3aZ3DLaxY08TVxubgoYyAoy67MrUT9
3FlD/SjFaGevqgsXo89H6eiWy4NvxC2o3oz4xKNPPeiisOs4f5MVB4bttig54t/9xiAO/7sVrRc9
v2upknr0qZqq6owxsHS3OP0zkaRF4RZ2P8MYn5iH4Wj7ujOvB/jZ1qNAwyxVfmJ7qEzPpZrwg7eU
a+Ui+COZSrJFz3uTXWwXR0BACMlembGeWHFTfwXfex4dweCpjpaPzMndKmrxP9U10Zsbm260ap5k
VoeppI/72+mRbONe16kTfx7abl12vC4J17vYjKYAgIVWNh8L+AtRwkXEVlg531ucPkgnFmbHv1p0
Soj6ncWB/6PJIxN7bVH7mj/cf9W7CZCVYtCHb9hocCifDMs8EjuiiMyBNbEFOdiI23MFbSUw+xJF
4mjodvfAulcZJYIDJXbHv5Ep5N116donmI45ZEHK1wbdYOOPePPjiN5XD/nX4bY9CQC3HHR7rpoR
ZddSKyDQNrMUNalGl3OUfyD2PT/ugUVLYPA6sXTXgRyNxxYsptWxDSSY94Si9FuZvXVF5hf4H8/b
X3yorff6181QkWA05z2RL+730FQDEys8zkO6oTBhmyCsWbKkZUIdTNK4yQhFon9I3pt8o+YMoKYd
b1Os7CSPdK6hgjtEnK+HO/0TY+N4zsEbcosWtiujVm8zC4qz8scfaxvbhHLxQYVLACxoP1PcETqY
gJ21FmS49zANHM3DoGgP6jGvAOv4Bm/yUx5fFdKBCMrMPV3y3u+rLBkJA6xxWFRid9o0+8nDtCC0
4j9fdoRBJLyNLRBdni054dl6EFpB8HNN88/uSCEtqfPBp9GuEp6Tv7fKoVWPVU/T5NhznGvkjlPv
A83W+mA4YTQM0olsScjvsc/759j0q8qomtq6mMhnhmv2iY1hMd/Iysx67daRr3Tfc2yZCcEKoQ5q
NlMCxE3WH4vPxi8syvGCHr1pUEiVIzLFHGtdTG4g5DthA+IdTfWBG7X91KCHC0ds966EjWBKDDdV
1KQzWYA5NATru/5OGjnU1ESPxiCNfc23ho747vhwmAM4Czug9SQmilz6yrED1dmJgwV+bNobpXo0
VijUoZCahEa93EvcEfrEZl2mWqPa+NMidXVAQrDmdqSZnG562Bb5ddHABqtA8yPQVvMP1QsP48DS
ct3LM0iPphUag5FPwpRkVS8O/dG1JMs8cWNwle2Be39J2Hbukl5IIKN1QZi4WoZOgNfPVQfzhuO4
qD3D60rECDpSiwFB8xrmLDQ1BmVNpVSOfFVA1z3oBPkuigWHfeKA4YcUljuPstb9T75oD4DJfKqs
TWLe/UNvUcFyRriQSLWC0s1ye5DBXCqyogFO84t8/MwpKtIKuaQmeXmy7gPMpJ+LOJl2KI5ge54t
VLJ/Z7ppckvfylNjuqta4SoV52IqtyINg0hjlkciL+PVFm26wkeXTeVUQmdlnTuhAiBWIPcFLdqs
AtKRrml8y9uA/JfsgMhcUUB9q/LY3GkK/UnjBLiSPAgbSkm1ap0LG0iUt5qTuATgB+ocWutDXh/4
+5SmLTsRzjtXFjGROVb21YkiWbeJNLHw8yLOtPhp0xz7YN8r1bWjje+lFdFYeBPtl2XM/5BB4GKi
7jZuPc0GoQIu+8HdPeKUFdzt9dtP2xujOoSztsedmq0VXurci9IEIyQR7olUrDJE7sBM6fZKKf0t
03BZwW7gutt0cVA86pP9PcypzdtDcHrCpcZY30PGRhLQ1Mc+ej6AR2R7Kb39BIsi+75et2LPv0rL
upi1jjCHS5CzfXjgCC/3t5aX6kpt4CvWiem1EtrKa5Yk1v5NICP7kXYrlcrZxe5AFSYuqYuDyJ7E
n7OJDvPEGu5WgRx8mXQcBHH5ALOio0tnpBBVLNTTeMjbLYVscVEL7lckoGbnQcpAGAaswd2ZS2O/
0KZpqxPmJCZsTbH3/uKaYtEca0SWXdaCD131BnlMUGYrr02voX/jeqzDKZEdpKJgjUiF5IAOGnfT
UrdlpMRyb41gL/Lfw7FoumY72xKIa8g3as+LPSQtCe3R6Iza+oTAaIA/7V/EcRLauBXW5Y/5UPr8
N9wjsw2BY1rIHyHD6Qs7GoFneJqjwhJRiO/FLmwLExlGd02eu5uaMxaYi6L0ArMelZEiEc9CG43H
XTMlmED1JCXRckyL53UZq8pXZSuaAFL5lDllAIcgnScBFTmV6Z8WfIGPu0crRLrGpddWalkzQMX4
mw/D3Mt8pFCpya/D2MyNPNfrOV72tS27TlM3JMIbEonA6I5V/lqUH2JY4yQhhAGgAW3vMDIwConT
R5oS3QKB3+6P5RR2iAs9Tij+8TQChfxRQKqae4b0XKUIRxzlenXSKL8P262zvZ8+ftc0GCeqF+YF
3i4ezo64So7oBqMB1S8anYQW7X6GcYj6Nv/yd58w1WGGycNym2IMnDAAivwisil+GRZ4DRlJxmL2
XzwdgIa9eV+gSNmC24q5InBLDyZfQMf7yhzjpl+uVlFnbSWCDMEZURVTJps396V9m67woRtitGSh
aRUUaAxpxLKO730bPrWP18bCnR+ve4+wNk6mkxqT/z5C21C+TpzOGR9q2TEJWwTebASSUKxESWrn
7zP2GRMj/nnZ4+a43Ay3wWF+uNK8RJ9ralSPxlrICu5s42dtfvYhBIhFTsodYy0GWHLp03epy17E
T20f0WAIFGXZVkkNSdIdQ6Tk1e/R0/217sVnPEIgDprsrOde2z12EE2U1Nwcf1pmkPwFFWKNfX3N
kJ+42N7X9PHn+//SPkKL123t9+4oPgQz5CC953NwyLUXyY7R+zkUrCx6Cs4WGzVLNsrdgT2+HODU
UaojUJENhsbVaFjjp3BxPP0iBCqC5769D10/lkK0Bx7uTEHx62XNqa0e6gqLi/33PRF2dgQYDE2E
Au10bGwSMO711zxcsRyI37VwMcaODHtklzK2psGFycjNdGxZSgYIzeR9KCX7cQT/kmuLDyzAkTkn
0WFkmHvFPcu6A3Qzrl4cDuwuxT2vyIZDptw/HKA5rrhsL+Sp2BT/9iKL4lxOZQ84TJFE1XPPuWUo
iNkf0XTX6suknIwL2y3mqfI23UDnsU1DuTRygC8/ohaiQZ2HPQlEOffBozsCmM9S5SbRGVl0o8mP
hjlB0JS4Pt3fB4wIbPC9WmCKb12f9vugEgwvLMk+6hZ2FNQe1Oq0C9H7KEecO2XRHlAYLqncKtTi
BbbC0/tX91/FtQZPgKF41JTSS6MfdPLJBr9k8qPCo7m7wdR+PGmTPrmk0CfMWTUNdznUaL7ya8GJ
v2duVUEwshEjfMCclDPopjPp7J+Ap6Bhy+FPeOq49Ff7Ln3mKh6l1WdtoqF9Ytw8XvfdMkE8jg7Z
dDX6kIra+cYGVXu45eJ8r1OzMS9+9YNhPdgtrxCO6T+hx+smWBxixIt8R1ckRk9iq9HtIxC8NJqg
/NWt8PH9DihpuEwAbmLIM/dqv+a+x41rZLjza+UyaMKVBFNDcqUW2kzgm2K02wrvcftqnbgTs28P
8uh0TXabzb25HgOzr7+qJrXzbxI+CN/VLD9lyrzs5Kvg/UUYB3C+98VVO/S+PhH8YCDxaoiFZAHW
M054TgcvPY+D4vHOW2UGn4S81gkplGwLzSYBW2Vy7SYXZwd4YG/tpmAG6UrPfHx/JvaXhG0XDOji
U5BC2SSHdCelo/7cLwqDO9owAAVp5Ed5KK7crK88PO8O4S8BQfM0CmpOjZGUL4jiAzLzkgYh2uzw
oFMpAzIO8u/ZBMAxoE5oMJGqcBftD9TdsccTyuryEGopoJLq6W5H0dpE5p7UX41WFyawJf1RkxuO
bbjzlJ6tSTVP/hzLiMLhyNT9+0dwhODAobtTHifePZZZMQsCDYUmdiJ5UdoHKWrvNbDFJHMcXodp
6XIkN94d7Ig2N2iyEJR1oOlYUA1uF8xLBm/zfuS10klPZARwLAwQeTH10Kh+ut5/UHpgTRrrePFJ
fVjeyYrWmM0eJQ8pwllj4HoSNyE+vqTELOpZvjm0WdWt9YH6i980Nyo/iiOa3PupS5+rNsgeLD01
8MdlZgD0jC1HLeQUAg5o16+MxGB6gZWk+fZlTxw/cZ8VIq33tZy8ggNBBgkUXCdFzLYQvJxH7TQq
/rIZaE7ZASsd+fQB6EglOthT3uZWw9ylUTfEuyzIXqRruTHSnIVOOU37PDW4qzDbpD5x3RBV+PT8
MM2WnsNJnmexRcBvzsPqMwpzb6jxALD4AcdP7hkmREo5IL4SG7dHqWNemcuFyeQKb99O5x6qxvyu
warCrJjqNXqs9qz9OMhh7eK3yN5rYY350CqqePU7bgvEfoiH5zctnBcvZxqa76mN9DVWBfJBDL6M
DeZBZzyQo/t5dMmUumDxqNs6TI444bl4ZVJuYa5t9MUDgqEZZ1oH6FBgXS1jTLexkyo2zTLWhwCn
w6glzRxiO21Jfz8wThGfXrYkAfTkkHhu9RWS28pa5xvsYe8e2Hmnd7mDFMZ4eFRvbfFqf2ycqj8L
xMkSZHuXuLcPneHrpd68Opz+jjKmhNRU913hu+hoNlOVUhcKZd1HkAfnFbExHO96T5bsA0YD4ill
9r72q8fu3gPpvvuFDtJgmZDiAawcuW3WTFq5ioTBg/Jf1W7M6AbmO/OvfIcQ8kZgU14KdMTXwE2o
aeWChbRDmSk5hLr5hcybNN3KOWDP1jROd/ySGlMegt7e8mtULR2NKEeHNPGIjEFLUcQUgU/8pizu
KVFigDQHuGVNnrLnRCETajeYua6lJLyY+eFJrvFRrXPM4SkuY7skUYo9izkjIDYnwDBr5zz/6Y9g
JbmuZVLCdQV7TeBRJ1UpJEeHIMx4fgOKh6JFokR/nHph3AC3oKvojjB18unc8GVYiexBkzaktYLh
QwhHyrijJV39+wQCzGfaorUHDEspPaMOJLM4JNoLO5P1T69hWWYnpJaqGY0iv0Rcno6PRSTcJlXL
Qh2ioiRvESi9GLK95tWF1UxwZujNkkkdPJ1uSze9+lOMNAfMXl5MwOMFUkxhejrpe18UHKaffvZC
Vi+HXk2YTmqtvwfEIZ4a98Na7oGFbOJJzKd9n1VQZ+J9lTNeSIHqoHwNlIYninwJvaL13AU6Joh0
7n/3RBncOsxcsWUsyEBHZzN7M3dU8vpj4tQKjf+jRwxjwyWiFn4iglRF1Q0EIT0TgqpaIZUl9Hkc
D2V7TPiKlr9LH1SjTSTvUkcfdBEVHdaLLSXiOxNVr/JX7/DYcdDXN94WGP87F5Oe07YSsvy4Od+U
fAqcPx9LvRHCwEEFGaTRExVMWgxoYS9oVYLrpfQnIitNTz5wpabagdZYPjswE8m75+DX3uMGFf1g
vL+V0g6+A4crNMIwoZlHA6NgqZzNSKvLMROrFCEjv8g0CAhvn9MZ1bQb9QAdK6elhHh9jS/dzn54
egg29yRWb55wrjZJPGKo5nApg/jC+cVMJO0bKC9LfzrjG45GI+0wJTpW+lR+ZxYSwQZOeUxZCX2L
qNEwsOZdLgUF5/63HBue+3ylzrr/Gb0N6aKqv9YYDdIkoOIU3eu14oXDrE7ee8IACfdqn0H60C1B
jHZSECHuMGeSi0ecVWU8GBA8qWL+CE8aQ5etFUTaQX5zUea/juJh3upmHZaVo133vfkz5EPqPsWe
Xfi7wE7g8FQhPOhtre88ZwJBksM9MBOdkdTV5mN01tabHrZyndeQqfHwg551JFKSQXjgQYQDCKML
Hmd2TdfENkOi9Mf8rMboBxcyRH/jQePopkDaCPBnfCl5h/rcZMYHJe8Ag3+UwF+r8StC/JXwLBNg
8X3VnK+yKF7QHZTUuESqqnwdZjJgo1oy+WUpuXVGsR6EGB4bsWgemCnl+G05iOM11sfYSb5PaKxm
h/yaKrfbt2XW3Mexq+axUmjmeqW+6t7rWb2/thJRKtkVXXvm6hQY3GcmtAIYqzl9mtPQ6V3CcL6x
LobL+saWJeb6OlW+15yrcEKiMkX5PxY9u9FPM1dsKGardIbtwRik84eMaq7LVYbKB/LG0ORqHMEW
LBsSWKPnRGRarphftv6hniNJCmKDmv/GSYb5QdO+I6aKmSSkiRvMDB1+Wgt+Kk55nMie6kMwKAx+
/HVR5okgFK1T2g3dAyRTKCEAKgS1460K/GMM7RqFoS/+Yp56IKtz80smKeNjM14zehCOzetOvYL0
B6igs053m4Jf7qL03DmE8aq4mti+DHH6iXbqemT6qYHr6CqqIa+zIHam3sImVXjIqWEZebLiNnnl
ORDNX2XU6Son/S1Pkcs3nByndqJva7kNhStsk5lRXFTJPbw6ceXvt9sTsWY+ZMS8YMYAah1ab5f6
d+peLYdRgpquy018PTwQDBGBbqY5glGtLCLBtWrCzbpKlllc1zdbvl5VTi8xVNUi9pKIZvRhtjs8
jvaehGYW4TZL2Lh9eMChRMRkiw/hKWKM+TiIaFT1pL9QsvnzKAGwMC97GBg+waBZdG+xEMQ/wqwE
qYN4Dac6naheIGfqCK4adFknWTKo3peU26FyBAdrqc2uA2Wi1X6YKbjqhvhdn98AP2KlJhBA4dmB
vN585Guk6z2uaMo4GYywkfe/xSUqN5AAQto6/jA6a95V69Lnrlqggr1vq9J3lLX0QSSrtnKZIRPx
ykXpEa9HxanqtDOpaOWLxhoTRo8zHW6JAkT35x5eLo9lqRw/dx/ASMCxZl99cmiP9ZPYyUJaEcA1
3e1jdaSKhWH7Ge4kZFhKHKhn+FVR5tW8GJfmmRfsIPDBptdEvCo1Xa34SU3ERPEqD67ORQYDIQdX
foOMbfo4sEzJYvzX856jzK+5thFDSUq3+INcTpZKmeYQOgaHuWXz+mPiAhlLnPYPwMQK+XimBNUI
Awc4sYJYmlgknyplBbWtPj8+T7eAwHveniBq6HJ/goskWcW4mvHLffoCnYacssOpzPvGJ0QQhsVg
iFd62Xfwmob2SXMzcguyx6gis1K8pZM0Q0is9sHlapEj5ebHgUKBkr3fbaKJg9ACIh/boY8I4fj5
lvNiFtAa8pNd0Ru0ybmw5AJibJdMZTpwM4/RHaXbKxGsK9KHT0YvsHZp2UlX7ZmWpheuiN8jMpNu
aHMh5+yAZWCS4ds0hrZfLMdv15XT+ERVXvzDm4iEk4xGfB/D0yKUqrDvt4ixTGhq4nMyGrJ6fsxr
jqWvK8ivZwgEgmGFQWoUiwcSdEwNcBN2gz/ncDeT8oiLCI4HnNQkRj2Vq+0qWkNDkjizZbGRaMsm
z8YqExPECqkYPnHluUpCMeJOeBV/KZLWOVOj80Fs5BqRdur5o//pK/L7retbh1dIiB5h+mXg9xLF
Wdux4FHhlFqNUGU8or1UbzIdEIG3NaNOFEelIfk6GjXUqnH2DafNP90VeXS+cvya6ftpPDra3sBf
R5NKS6EnGxQ3akeL+h//vpXvHnEJpBJAYgyXwJInjKUJP+4T2QqYUMev5rZEn8ozdpuFmX0sOqn6
ZOoWx2MiVpF3Ddh2WDlkiGvDnvodggk30qF0IHoJg5wURcruioI2veJiisoCaI7NnG2fFcUiIOA/
NKc8K6VY4rsWiksTa4DyCzXBSXuuacLxAdcQK4FOakxRNT7jL3fsJ+aQhGjcOnHjchTQwtExDDb8
xwGg0AooUwHI++aATU78AB3fcI/9NAduZprf8CH1fKg0nsD7MHy6b0iQgJtJHM/fW5ZXNEW2r5Oo
DY6EA0K4ca7ktPhbPZCdX9amxrfcZZAXhL08Lb5dHas29UU7CR3DDVHg8sq7uU6ESx28dtL1AZNF
CFBsW49JOnQhn4KNWiAueSUDu66KLHILX5VuJi3KJ1rTiJXE9D+4wZoEexRlW3JcaJnuI8mlRlrD
YlDfqiyDoeezx5UECxt/74KBHOMyQpqu3aXtpOsY3m9Z6pVPQsrw3hoOhO7phvf8s08ypD/S4pxX
8DJG1LbDAs/RsN+C8Qya8JI4bOsLDx5o7sPZVCOBZ0RcY5zizH7eBCDoKiYcMgOee+VQFxYNElF7
W8I7dLSTplMPqkC2+9PgaYbXJ+gx/lGnQZnDMVh3u0/hTi2/t4QnCpcNSwEetOnKsaOHCLYX+38G
tW17q0sWJ0YrPl73ZMok591jnes+e7nQe/g/Bw5zLSAz7Rauh40wmAfK3obY38VrYgNNSZzrz/sA
oZZm3lBvyZhxxSif+QggDx2zZq0RB07I5G+d2NWIzCmczQebQbk4cunzLR9lFDkLmUUim/WdE4+X
AV03JMmXgREgWebJllDVvzhCZHi8/HhqqdmNYagLDDTBB009IMPgtp+7ogIjRjF1mzDf2wY1Z0DK
pw2d44cHz5DwxDKeCEn2dePnuPF/0Io0xU8r0ycYIX57vBA/Rm4ltdpl0ytUrngW+GTy263ZJLVl
+0fg7sOZemrLYhYtYmK9iOHyiY5amcPVX8vA4d/jq2QLL4fmdvNOAvw/P664IOfWzIHnYFc0SaFZ
D1SHJ85n4a7k9plbZAx4b/lpO4y/UHPKW04Rz8U4nhzJSPcE7YFVK2PzGpz+h9kepLVzCku7I4qX
/sDJUvWjObvsUrnXneUKNGZZIR4t0ZWo3+ReToOo4bfUX+VhFq3nlzJ6IpYXgfIAio99KhdkWAQ3
6U19hM08m5xl6YANIQjspLikmET3ncqZSo8yRzLf3kMIYNAgKgHVsgYA32hhX4rofgY77JicH695
yaM0TsDdorOvLNtSGsha+dxdQZFS3j5NRh2e39ElnNyO+AotayvZvtNNDXHU5UfQhiVEhkRGf7sb
h/gmvwJg40ynNrWxfwIGvl23OLoLSbwiQ4kT9ACrIQ4GYJDGXgdB52PJpw3Np7Aj09KRzWVML5ph
AMeeNxaqP5YdYyrA2D4djVnmllXd+XZuBR7T7IDtEIrfbD6pkN3RtIdIVJNLDCkjVXOCLt8Zj2Gy
fM9boDDCQ5nKYBVdqY0gygR9IA9D9ALlbFAAPNGGXWPZ5OL7t0BNmE5GLakH0ZO7Fq66+mg6D4QS
IxfoRVQvuJ3ySmMtz/LIhwMSaFFwU/mS6WsFI7Liy1FD7vEGqWGq5KSXRy4jorEZ1Ng+MNSvi7Nt
acqzP0RcDssYwr8pkknoDgaaMdznfVRZaHGq94JjdpbaTOKPgRTYOcY5VAj4/lRy1zM2bsHDZCo8
/eQdYk1NX5R5tNwPmgYrfM87JU+iq9vKQdXnzbtBVLnvahiN63plYv0jxF3ORhx0TgYwpoh6OtAE
xe7hpZfeM48axN4VWwqbT731k2zmfXKrPrSrSZN8+1uspe8Fcyll5W5EWS93QV57w7JCzc0hl8Ok
nOReeMB1s7dO6ixcY76Hc7DoPDtPP+nlHsdffqygFd/64oNGIiEeYIbMsNvDxwsvs/C8EfdyLsRj
Shr0ZTMSGxO2UMCSv2kqaX31pkMToYXuoV+Rz3E49Prx9aMbnAA1n82f/Apu+9PkJUSAsNZgg6s3
AqN5OD1+yQqyMdc6M/+s5HGgb7puGjx5Y6VIvCMxAq6+DvuVcLVW6wVoyp/kvZf3SLYUZfmooAJ6
5sV92M0I6CQITmvDj/sX9RYC7fOdrvcAIzmqMvYE+zxO++6lckvwk6PZco/HIgvII7RaqAj4BSGd
FrO//V6bxZ2FUZfeMPUXcqtFnrrzeOsFdB4dWAdCjM0ktTjIDI1OfiV3Jt4/JCyWOc+lrTqAPgBP
ldsKrCcuWEFd/BdfUeeTXp89mrrqhpmlcRK5vPzZqPIH5CbFzNP7OQvkzd2HS4Ngx6qC8agw0vkX
I8ASncNbvauVC0/BngYUghkRmahLxJqaKSB16YTbRkP2rd1ovSve8UPZGPDimRq/YBFRk63qYyuv
8pcuOekif01TvourHD+HmYeDEmqaODS7pPlp1DjiGWOeTKHSMgVIPYqaGRVXIZIBeM3dGxkqZW+9
BC75teEO6rk+jnsgKV8FIKuK2oD4ZfZeP3V7rpr7aHoSy6wctCVnwew3YRVvwPd2UL9dN8H+qUrs
DnehQBClM9ojCWwP1yqc8pJHsJKz8i5tCX6Z/Xh6uTVpXQ2M46VpiNpxONJAIhzeDcEtiON/+W/Q
ChwZO8gxTQ0FHIgDOWXSKRbZSRos4mHuHuftthNw+z5Uogi/PIECDqHouqrA7+Qd45WIkvJ7mBL+
noyBEykLDPbCmlR5lzAD5MtdNIWPeg3acS1f8ApVd2kA9e0Ttv1ZTFocGz+Jo4vGGjZ47y78teSS
PGdoYgAeerUFyD69Qf6tTis7I+VhVoWyFPh6/lNrYwnl6DHAReOwCgDiiehHyM9U6Z3rc9pyelnm
cTOccnlMZg06it7n+4lS6TNlme2r6cRpc4XSilVlMt+XFk4Z/PMmdyyMmSo9s1CkdF83i2BQsHzz
BIfT3lpmFP3TJ2c6wWVTttI9hj6ikz3T5XESBox+AiAI8pRJRpVSiXt2fF9ByvLjH7oHPzbFuCJN
yaJnPsspfxUrpj4jgj9G+Jg4EJf0Z/pr7Z18r/vn0WocsfJtlcehnHPtjjI4lFgUwRVJYLi0ITXy
VCJhyuS9q5Os8RPe7QAZCXtyHHsjqFuF5GguvN38vUOsdZF5a8VYMAqPiC4S/QDssZpOzRDikSD6
LSvXjdkb6WOHnMa6qqUZHnz2Q3rN0n5xdi7NHHeQbwSVMUpwY02eCYhrWE1ELlksXeIpsgeWTwT3
fjvWncrtUvae/R4f3CraSAQY/4uoZN8rXp1ahRCeQl7Gk3hq8vO6SIug+VHzcPlEGc3qoHDXxLBn
G2SB3aDz16iR9i2sCbIWR77yNa0fbaHIemb/dPecrue9c/QLQYXgnIT7nwYzNr6dBS/hcnMo0uFk
XibEa2AGUJkVVJQDvFa8MrxkCNgzo7W7OR50Fu3+Mp/AruDhZZvaF1YKwwYv1rhkdluNBhJD8i9i
qO0RVLleuMxStZEVr4XxS05YbTtAWqDNkSxZ0z2/SUCmN195A54SiJjEj57oDNJqljdcsIRzCPk/
qlLkX3DEiNqYCY9Wl59zyFopda1M8+SS4iR+JhU3mk6eeHl3Z4NppFF64B7HFwbwPNcrnesK8S/a
oRmeb6pOHJC1gW9be7dOC4fwUkTakZQoAx+oTM9Fsr6/AX/qBAxDR6Fzm04udmeub7JifoofJmlf
Fg71jQhjShE3aeQox7sEKEIX4or7U7FhZB2e92l6pds/u5kiarKubg4BGybpPPSoIh0nMdcvvSMt
SYEWkQzuZ5vhqk8Jj3fKgY1CI+OgswQhudqDmCwTVcJsDhs9VMLqnRK+Xspirv19fHutcwDDu4bs
oyRt/6iE9jLK4ujg2eA/llJjQ2q1zujgit4VotPBoIXhY/kiC9RubsiplfXsR1y7a34NTuKOFYMA
FC3SwwqYrGadsWmctTsUtGt/Fdp5U+JqEYticmEl/6svGBJh+fhZavvuu64Ht+81BT/OdB3FEnL6
EEhlujWinbeUWPR454FA5OTrulCMIyBgXhZVrvOTQ141fmZPlnpw6G0cdroAMc9vdnqzEjoyDKo5
udI3MoTA2+6u5kpBLqJtci43uu7BiJJfRxH1IdzO0I4h4wpBoFBuVpQnqFIrVYdJj3B8eA3E3Zeh
gHJ4BhSRxgOGPYhyVO5tvGPyJUhy1fwthVosiAAIlM0ZLsCm2IugZO9uY2n+an1CUCh72Z3E+8Tu
jXkpJba6xW56L/HdVBotULG9GZhKsFwn6A0yphldFx9vDlJh5P3f8Ee7x78hm1L9z4ce3rI8neIU
5xE9RAuUGdGnSs7RBfS6H61/70NdVSMmzOtXZq9xEpJf8ALk9gm8IzhbcRAw+3QNO34w/twt4zjs
LByhX23YajuTd/ZiQLEK89M5Z0k2S7VuMtVfFYp4Z7ENbJ6IcTNSpSKZeZXtLTHtuMuY7q6bS0ip
WJ+D2drGZTO5uR7iErfvU9W9xGTFZM8DE3pyfK9lKS3QbKu4NOpbkX0sl93TJ847UYDXunB61xMl
TK7tUqvG1fGL/RmKu8iXg/Y37MeiDj+VJ5UPxgiPqfD0h/bUklxsY2/0DHX3y5YcmzES1sW5VGPr
LnKcIRPARMtBZQVG7ChcDiZh4Dq7AMxTjrJGcgDTpf57bnDpq/HQKs+rgDe80EwPWktyqrWRUyUm
FL8KfxUlOO8pDV3TyghDAXvPPzi1Qd+byCd+0oqcnlWlGyMAnZ/49gOgpylnjbMxy6ZWYdi3Rwbx
dwcGf1I7IvoPVsUjjTOep3aX0DunomtrwjIkOSWvuPi1iKC0PZlYV7NSKgkAadj+sMn/JR05hlFA
zegJRiCGin8qY+U2lcFFmNUsrh0AD15hsZPy4tXT0S7TAoK6D11P1ZkvKxgrSXxRybxE9yRk5wY7
fNHioA7FET/GgmDLQMPWzl6IV7bZzlOsoTYzc+xWRXus1bQWfNIU4iJCR7msSgpaMysyqUKiSzsq
ddLU68NQZiCcbhDsy5Pv2qOUixjy51z8z7zlzPapa+7WkjPKbe3q6I5vEJ/TA1CZGTaY41r7RJ3L
rWST+OWbSYmNCLRZwlLnv9RIRtEJqBEDYW1Z6I+31AsNPGIpDNMtDkhyK8ATVm1DGQuczRWCAJev
NJ2qgmKHnUltUksodThq3OUU7b+KH7i/ij/sAByBEMOSMu6tlmjokygT6p3j0nitPI1i34TZmQCY
nJvQmhAzx9zQIJjL0AGUZj0+ek4whLKzq1QnQvRnzGcm4g7qEBptIclbXrWwVEfl1poS+huMpSnT
ozIrp4vCUYTXubVVwpvCgW41Ak6YENjxlPj/4UyIwFpo/C7TPf2dwj4jxENuz0naw8t/fMqIy6s/
vBR+u4m3wU0xVG0GisQuXzYr+sAZtle0hBaL305pX/pjsv/FhyFaN/GV5yiUnBsAVbsQWz8ujVYR
b6S1o2nsuBAx7Js9vq6s12M/hzHMo/lQtPRryKxBMpWH46GTdl8rjCFrNGQdRu3dRMc9PfF7IYnF
j7NYSsYFuF01akl0I3FN1xhW1Od2E1RoG2uv5EVxCPQMGK5wKaGq1XfhVvHRC3CStb/e6myXRMne
JKKkTAzm/Bx8WGSP8UecL8kHK8amdJbFtm04bhXp0DqcNPyuKy88E7iCnkSXr6rzTRWI8tXtSWSi
CoporZ/Z9iQ74dsMt6REDbrQ9NW2jJBiCutspNVJOJajkyNsFP1vJWKbPGG9J8vZ6DPVFm7r1nVf
rBqYkB3s+cs9jktgxhHtwxq0ZumCNFhdcnbIBfIsnFIx2zuWGkUAUDOPBMvdel7FqW+mJpfpu4Gq
8ScbXDOxrPqMTnDX+hBdH/mNEuZGIHgf30G3Pkn+JAuuLS/peGH8rKAGn939xlV+wG+X1IvzdAyU
9HzgGB8c/1l1wvdp8SyHT5aJ+TQ3T34jmQoe7exYTufhQUqAGvPgovqLHJSjWLnbfmeWT78E7rOU
2RFssxEig/m2KXKv8Cq97jm2RypccbyZkuVJC2PP/sLvthVMFS2H+4fZFmAMI0sTiTeRQjfmUH2Y
nyt/nW6JQ0OuQrxVAr9jr1uEhmC5vrFiqKualoXKtq7Z9RuHInKjCLKLuP7HUv+7NWOEF4XQ2cw6
HtABG1ni/ej5qSogGx4oS5GRZgEYTGLkAdK7wTpErLMoabscXfK3uDGLqDL9ZwXQewny0PlfrMjO
oEjur4eWfbR7abVoQigIAebOctQyrS/ok+5EZlvtQf6cXXI45mQ7+GAjS9AiG5zkpOUT76d+iZwx
hSq+ol9e5BG8xlS1ea3OULgle8eExLuU8PwMpdQtU74O6hO4JohzNz7aoTgtyEpUtlDDc5W2xBp6
dL7JI15fuEMNOExRiJdnhv42wYblcjDgQI/X7/7QIioJFsLz0dYM4c/OuLS1OOdZZoiSdkfv7/0k
71BrxLLxanP1V6YR47etdqSBrBgQF988T5UOlH6irQwSB0wbV30VuRTXBjdfXdBf0qI3jK9E73ad
YxJCAC+VBRYkErfVQLiaIgoqNdJ0nqrCfR1H5VyfHYgz+cjwZK9m1P9bXr27CPB4qb1wF6c4+/5z
MixIAdH2xqBSsKXQqbPnZtUADxW8zrkPThvKmfkfwtkh83ytPObBBtwYpm1eeRbOz3RkO5FTn74B
oWnevT6nVZCIpFQTOkMoGuT5mXtqSFrBReC9W8wLOUNtHFl17Aa+P+4yGeP7zCSnSmKacz2PNPV9
FXQirU0ZZSqUbYsp7PFWMep+VwXRDL2OGnRpn11ZI0rHnYE0FhTzCoaiCx4GJqi+vR2TgRQdcAmW
MDNiXSaXrFngl4zKd8O6N3kntv3uYWyeYjIep61N4k3exqeALcQ03n6ysByRFloKc1AWbZ7+EwD2
P4/+m05ay8wsadxCuQBWGF4He83xqyxmS0F23ORxuhLjUkS323/v8fa2TmVp+Z2O5LZXhiklXSC9
Z75x+Ap9ApYdm+ruSoYgFeiDSRrlAtlcyb8BWWR9tS3p+8PBF2m4JWjVZywu/8c1IeUssrV2vNuN
0sdkR6WJPAydV5nHrC3xppYzXIPj6WA6yeHHPNYibrrem0G4yc/YxyAtDA6m4Xb5mZ3KjR4NtIog
TI7BSgvEAK6EVQuwlkG1ItW69fKV/SqJ6/MTplyzgJovfisdF30vYMeUlAvXOzVP9jAqaPm/w3Qj
AQxLPfUK9aVd89G2pZUfN6d31L5GhtXRefjNy0oLfcih2FC4NMkykkZglBAw9ie0ItsH2uS0mltD
7JfBmnBPI2l+iHGhqEMgaV98VyjKc6qMQEsMj1+3vUPu4ReUl3KWd/M6Rc0NxqqXVlwDgB16PxiU
bjJqh05wEuEAYwiR8G4aeKcvBtNmIevGACWoVprPNYmlc4Xbhx5AC1Rak7NEbfhnfutjTiNxMQvC
aAaY1pL2ajD7PL5+SZCRv9uQGxROrBzDPDajYABOKe424h0m5ICzlWWmQCclDq9pyiuXpZioPXnb
A9O4A7pzvorXlkr2pY34ShALunvcgLxMw/aTMfr7ZLDNldQTrDazoru7dp2EsUFEdFAinRim+Ie/
edTzoSTs0VesAoKjF4zMaykFADu79bRdBaRxrW5mdsPnVmPUIuwRHIBI/I3BmP/Id6sjRQ4e9yzk
yAGC0esUXhLOTqT1E2zmy/siIwASxbC4mfgV9lC9ARUnoHT1SoD9vT3cojuQoP4HRAZhuAfRE9V1
40cMWV+0DwXrZmRT4L8rcMY0ljLEa81Idk3shLY9hajVAZm+GUqrlz70BAfmUVApGlByaXzs/TAi
cPv1eusCqztUYpMPgYpTqxF8JCr+MmaIIqtE+jMevj7r45C60C5rM7xAnFAa6VCG2BTz8jr3GFXn
lxCo+kJo/1SYxqGXVxQlEMRAYrC63+DljW38Ous4FDwzWwWAj9jANqvUY7ZSVjjSRMuXnsP3Cmhp
Zj9yN4IS1eJyTBT715HzGDbAGMVEMqkYJnMIZh2c5C3x/OvEbD9kEr62TGPLkGI6PGa1OXuDMOqw
LTJ5JVZvU2JhJIngzrSCEVQlrcSAPfc1MFqcSVYsweireqw+jAyTCsvxWsPz3ZdNwDUODpKAwnYv
GfhGx6TYA1utFxb2A+he64S7YesdIo73ShfuJ36ICdwF3r350ThL2yqBCsMkGy6+lrXrQ4mbjALS
MQbJCunDyBTOxLAtThsO735hnX2/xZBGlidXkdocR23ZvU1s9SM383hi/CRAx0CrLAmlBthqbZtB
+pW8J1YuXCHtt3RTaGpuqYC0zs7x4zoZVmolNSM/4/fCLE4xCiyzFDTrQjewdhht1PoHrJjzF5WP
Qmzu/NHParTFUDj93dUttgObPKM4e+FTn/NBrjVUtnBuFd2Ykrdcnxecsym5isZQ5twcQYzFENV2
24oYJJHCO/iHLPl/+tAK15bihcHhLZRP8dVH38teq22XC+B5vgEknNjDtXt6RMrVxX0/rifjPfo/
uI48j8QYp1NEBIGPJPCFu3vV6y0C121QeQ52iGo+hyCvsf/belzL87Rc1WiXj4bRcqV0zu+KwEO9
I09LivDb961xnjTFjRFr0fhKfxXJU1pQLQ3FLv7Tn2vBei9XeGegnXmfaRBjmDBLIAqgxg333uU8
peKflhsAPbCOYtkAe9nw/dlDf0Fw2Fmu3CLCSIgqqVQUv75qM3puXG8Se6VBEHiT8nefsuaw3n1W
9fdj1vFhYTZ6WNJM0o713CgUuT+41ITRe49Q7JL2aIBmquQL3jYvB4OwEYMX77F+8m527s5P8cIy
b/7uaZcab9D6ZZHYGulPVZl3LBXxVinYEOZ1GQHb9LNazd098XnLGazABsaELqBEhhjz5dt0LdbF
o+wknC9pk+tiiLjXvPxNYmynrCRQiAPXob/63E4jDiZx7n4syZZ+dNAVl1FyLY+owx1YB8+/5NJJ
9C3s47gKO/BwVJub4BcGn39w99kDq3Y1motk+68fc95X84VXD2Uub+DMmEYTbb5V0Xx/gi/0o7NS
/dBQH07Xni4FqJyeSkUhqjRMHPVM2gz/7ClZf/+aROr3Z2fpUzB11vRCaeelmKoqjhAEUxXfgr5F
MV4BPiJxcE+olLZkVGeYVmNiIwEnc0fE8eCYm7CSlmmoC8MQ8JneQwyw4RmSnCwb4hCw8uCdevem
F3eechKI0Qk0gGBfuaus8BnJBQgAezqA26+XTcPrxyITz/KsfO0YP60EIIMBKEbuRrKbElOhXKb/
4+3DPDNLXPonjYSshaZ0XuP6aXHrobNDLahE7jFGWsZZslXXlTUSkGeLUMvpbNhM+FKeVEJiYxR1
tepkNxBCsbZxUoQOJcHKgP03dxC2aUpVD69Gi7V0aJSWfHuHXLk39/pPyPqT7SkWR/8sgQ0qqHhk
KN3H09rHCBFmrmTVwdir1lTVSSY9Cws7PIXYp9caQgaiFKC/wxy07ChEzeA9h64slvNJU3o31Ksq
rT8zyEDX6W3dnbidZd1S8lZvFbsHMHGoHtZlIJh13pMvPsZCJaJT1QTVzfgCiuuwt2CW/d8HWdXw
gd1ZE2yZ7n4bszcB0U2ibmhLoarJCmJQSjj0kQrcrebGuJ44GpFfQSyDYtFzZqM5+vLAQBOFV9Az
5rksl0BbrFfPTEP9wEI0OowEd/N7JGdZ681xzoIGelXGPBESwNd+Nnbb2fLj03dH7HAJRDaZVJBs
w2U6dBvXoFtnUHdQhN0c0qrvFA7xP0ZvgiSzAaqwvrXuV1NgwGktsQrYOWzofR0V8L9FQIUKnzS0
qKwzH2afxjBILATF1tPIS6YUV8VzpWsQOHWwCnZ3euvWxt/ogQoyP8jzoUv0gRIShlH6/Ws4qHQ+
iA1bCM+JrGfbKvzXuxJ/x0neRh3UPfC6rpFLzZsUYq7bPMjrOYUQp10ubQ9p0ctI8/+pcqh+9lSM
O3Bfnudb5ywqz8nhrgw2Jj0ceVAXLX2M8HsmleSu3+s4uoPwW0pW/jpVa0X3nkJIOCv9oUh3mUaX
z81Vy9Re87bHhHdGoEFk68Uqpo4xjnP6BYHlXvK0dhmBUEFZ/wSBMOZhgzj26Dzu41rYKLXCmCj+
wdOnQ6g9qDPef4axz4SFJhArSrB58Ep7e9oYCYCPVHTu+OWzdvOYlpZufTOQaOXAEVd9NKZsZJ9G
B3F6YGXgpsSYYnYIJsxb+kxlOp+9OGG/6ehTPXPmIArG6+ProRnmduQho2DqJJv3v3zvwSm8w82G
1Lj8hFPFgC9WMowyeMtcwJMCnJynPs51Acq2o3kFHVezxnMKP4EoCy1uCb/Lm5nOvSQvxhjpzq8D
DNZP0AScCRuMTaMyXN0sFPRVrtfaqCqnklhaU/2F27dBcWYAxEP4CUbropTRudjw2SmulNpLOIIK
cRNHOCpUFvq7mRVNyXNmaGfD/Tcm5uPPV61tWTFennHLqi6LbHrvAIW1/AGEF6hPs781co7f9UHB
nx0sxIifyCTSO1cIevdTglLdFUsAihF6JkMFi5LKVCenU7P8tnX58otRIEgZfsbz8n6jRXSHbPeL
qrSyrfE+aJJckG09XTjo5CmIovS9kduFH8d43FfmI0qetSh+72ibF6xWacPOWtYmZgrRWnripRJG
63M8RQy2W1GbwhXqmI9HjgYa4ZGOmmDAFf+89SZbgDL7+lI0yvdrl/dNTHHAoUxlmk7Uo/YmNp1F
rZTVSDqz6rGQjAabHJSpGvjD9f6+QuBab7JQ8Kpl8a2+lnkfm67ZW1VV5Eu+QT/2xAY9X+S2c5rD
kLO9QbSHOKr18jRYqoVSc2M6Us1coUB8awGrlpCeYQIP6ARDKbu8tjQhZjb0lk6Ss8rqaarYFJlJ
qSX52FAwCd2k0iVFsXugQO3+2+m6gQgZDuvKReAKEAkgwKY6Gn9W4nB/vHnpRB8DtILChhMtaSwR
pqilIzm5rAQ2Lakozztj2JNwkSCUXFA+WMZNi73xlckZ06dipEnpPXLVOBfdVrdjOorqfld2dAEh
d11igex42XJOcZ6gyyha2h4/959U9uoqaPxyQE5MwiKXYmy1BgClV9TVC78FLz/59+enK0Ei6ZSm
cmgSchdCcn4pXymEHdMH32MNMLiEvGHOWnmnbWlhT4hRpKql7KSTHcP64yZPvnwlByfP+rDkJicK
5vuoP4h4VsCmDTv/0o/phRNzsyx/5yLQbfu0joXbJJazQoe78E8uRhiDrU9JfWBezL2xXDYv+bXi
5qh1ebmQ8QO1vr+Z+orsvTnFm+dWRfkQ3Duuw+3+icHNmdczo2GfonXw1wGQojobW/j9orDDJBJY
/6g4mFGnpUxkf1HWC38g/zPNdUZRnS26mR1BpFIuM+S/ffSRmdHv42aMCivHYWd5r4tbpJE31anb
Kb5Li9LccQlanbzShv5o71YodughA2hIGwy9U1J6FvTaOH1KE2mWWiq/iyyK1KV2ls1PXxDxTJAV
vKoy3nTFjsAzB6PV7U4GKp74A3E6RkhzsymZ82dCZRuYEuhD6Ta4dNIE8AkbyfVxPZ9qBJlaEtEE
XeF7OS4Kj1dkI8o5OpcNGQwAaPTPJWhdBc76bhOOEANksASaStfLVUMvoLwYV96Dz1lwZZxY0mol
PIYWLN+msivFsI1JwMkN9Ig5kS8ZRo6hZSBmzkp84KkrOPi4Ael+h9VxI7Jl+Wsxg//XssbYwG2/
gQk3uiFUmFYvSn+Ku34zmDNxoLWeKzI2etTl00BV7CBNHDYbu7ualjzdsh6XRRgbE8jBJI+2WGyD
y1XYtyzg+dFJrFcvu1YpERq+CDH/0dac86A5O/5Q5M3Fz1mgGiDcZPp/1888jdatIVoiDYfjAs9K
1kSBKmA2T8N9/1q915mJUS8QvYRbL2jkSlFxyzWAZCR+Roc9NRSlcctxbXXkTGi0iMmQms2jQNWc
AVs5m3fBk+aDLEigzYXeL5sgXeWhAM6jS8nKQFe452y6EfTtPUH3/FXJJFJHg4Uj16wE/S87KqjI
dHdsgwEKqzwNLR1/aqIweRYdMr7KVqhEAibnVod78Ewl4NQSeRiQiTXewv4KIOqGR1qngIbUf6Dr
Q5ZB29RUmHDzLgQKs3s/ML67GRUOhsDdP7AN9yod8yLDjt63rbjsgpswceuOpoPxLAhD0ZShQHmA
ECukvVntr8oWo7Os/V0vsdjBAsDTC/IxTuxUJEBU+3uw4ucpSSHbuLNvR9HihNHKPut4M3IQVB4d
bIRP8hD1iH4xhfFGfLR2CA8kp7WUlWzZQyCArWS2XifOl6XSOxr06HcKtGrsKCZx6c5ZslwHQZmL
fXD4zfLrjyzwWwps+3qktBcQ6wov8uiV/FgUnjNP7KnifU0GomJEUdIxWdKYPJIQXZS3PezHlHWU
3PFdpsOPUqibR4mwc5y0LJUVLC3bx8YyzKK5LMfHMfl97i1K24vGSjY6VVDiHm91l17kFoSQi2my
2SmBUIcjyruDaVUpVdCjiB1Kbxmu/eTX5z6uYg15A5ApCb2Gdrm3t/KSCr7dW/lr9eE8R2lsm4A8
rrkPUbgyOj6hEn0eB+X4EF39nfG6ZBz9YltJ89uoFRjQCpM18vQ6SLYODJ7KLOJXz86JZkGZbZMN
UsllmW+ve5/uWPeCSSeoR+ODsnXke0x1+TezmnAst8pjCkSMFSo+ElIqDik9PDoDSsn7MSOGsB9G
wYpG8cEe5fWD2z84zgOhW544fYS8fFp2ussH7fuYZp/ukzpJoMPtxpSKesvV3k23kTYuUC/6Hw0w
AZ3yAr+puYt+No1+saijgsn70PXa6jeVLu9VOFxNw9MjjFMlVu9/Fr0cYuGkBtPA3yFSC8Pz+yeP
/8ZD/7kpYljUjC8zvUtEsYsIKOaX3WkZ1Yj3ojnIXq6XBxfj2nYSiAEgOIieXyfcV3nth9esLg8X
VrXl+JfT03+J272kgB6Xf/NngsIA7+O7zcyR5gVs7twOtSFVVxNQrgROjJcV4pMslbDMAFVkXQR2
BLR92nR8tMB0vHdJ0HOlqUvngyMzEKfLTqw/IqOyL+94VhIogGqxr+p22uMulbA5yPYrDjKwy4QK
R8vksJPGQPUsUXK2Lr1VYYE7Yk8+kyInkDzS63hVuZtvsTNSWyA77gfY8phzatVPSFE0OKiyci/+
bAZLnAqQBjRJQ+1RXwBzbv5Y2+3pTXYdQQ5rJOad/PcY1G4D2Wt7iU3lRugSGuAVN3Bc3D0fv5io
oZbVokC+UNP0i5wh4nBiQY1OXxkyTO8In7cQEMZYhno3PLksmg938ROxjKNsjvPKpCTmup+a65FC
lp9JWImjp3ojdm4isWLOwheHSQKQhjN4D5ntmSKbRY/otkUYaMACdU7V3D9FULxlgsuU+q9y6i05
EopYgPSYDcYG3kNJEPBJ+L5ds9rwshPuDYrYJyExHOEEB7Xy2uJiZiKM5z03Zcb24xSErEBNTqBa
r5oFB/Dy+9TjxWbmLFZeENQLL+N+AQJg13BXA8Cz5eeVAPVu1ml4RPbZ13XJqANjfxunCC8FMDYx
L9ldS0DQy9m1UAdkB2ZM1FhOgbcNtuzoKWLUacnvQ/xWDeiP8y0qJX/yV/4nhO0NQUNEKOsWdpWU
y/No0AaDu+Qgv9uwf+OXgO54DG2fWJcGQ/4++lwMO6n+w1pYka/z5+QW1A/v2xpxTJZ3Ty2et7+e
vY6hUuujuSJc6v6Cybf1qhbMdccctCc42H4aGruC8Ogea4gO+erSgi5IIkhzOPGIzQMGKOLo1fIN
yVWgaO/LYmAqk69xBKGKx4cV6snidiXgT/R4yAQFvcA6n/I1C/PsUJ0/ZIBQk6gIeUSmeFS04jag
wBFJaP3WCWChxRT8AzruLfxYApw/6q9QOlzxCAM/dKeQlAHf76pI26ADYP6NhLdT0zfIpY7+J4BY
nSL19kL1icyOVuAH0P7MWI/GY8+2WNPejkinrknUkGoVJbJdP5r7UvJqH0ollOau8WLPmT4mhKSD
cdobNLyPZIJzpyrxo70FfEo4ZfSgwBW1C4z2NRQSf3gDNHecMKFTZ2Cwa4flm0ltDqTBw5gXzrlf
pw9dhAZSnSIOQGjXdTH/qw4R0XLaUbz+Bx3Vn15lyZxabbCzHYApbBxiZH3RkkblOkuPN8eimStG
N2qzqFo4Tnm4AMR4tFRu2MykCqfE3ioOXAoUKGTH9OyUiV1Lsvf9pl+GcnLvr3MUQhlDJBTUeqr2
T93ziWk/OkjIpONeA9z32b6eMAO8SVbockR9bUrnP2tpe7AP6nQaBSilrZYOQejc3Kj9L5CjdxU2
G6YRh3dtBW9C/SPeDdhPRR8t8trOcsqsTD6xQgX0xcmNqQFRB7xQE/ZACIFZyvG3aCBmi5Hrc91i
o8+HLR+WbB2cuFnd+26+M/eIJO7mPo3E/tc5EAdBUPyBOatbd5z29uiZlnvKSfl2/dBwoTlzweAf
1aKBiKNWRPIEhelfK+Oeenyx+4s81CJ0zr4Lxpvj6MVodQq2IjEPC/BnM7jbFrsYi8Otur6gQW8q
wgcYwmgCbs/k74jLsU7+TaZJ094Vie4HXp4+DNz5craBiOLuJK5/PuUgFr+MCsgp2oxriE3OuozJ
VQVQAzZZ8Z45FhEksMPrzsSzS32etKZWj902hX5je8QfwoQQF2iOk1zMvUCWHupo2kXkMHYu7xhf
XEwH4RwpV6rnRuUaXys69cJ/B/aLSR4K0xfEEA3HPiVUlRilzHkRDWzUes8VfmPyFUnlrCDun0dG
2d9HjV7iGmhvxVYCyJ/9RI6YQRGIhHTM3Fa9ODubJdKOv3ewxRRNBkiqtF81tJG8TSDIZJWuWS98
d4AnYhsGNmiDEvB6Z5xL/ZOKWO5QtQUVsHcg9UNWNy9hTv65a71azbIyxQ/3Y8tZKCuHC4xboVM/
SfUtNu/N8cXzma51Trslwjl2BmROa9OLLLcjRKTB1IisQfeVvmtMT9HjIEnRZXjME4HSHmop6XUv
uIUHtkncYvehQn8UmeHSlwb0GEc48Wc8lH6MCFTAx7hRi4UCHYsG887e7Uft7KGh5UM5RZ1aXlj6
OpJIPpxFltLH/WbYb3wk8BOQwlkPhLWfANVcjNXTeY7Eb0g5Z1BNZK985cBSwEx02qoH8uL4Zdxf
zXYZ7RWuRiYx3R67kjt+23opVMPstFO0TaU0P228o7UMMdXXsd2exnAbTFAdlOklcO8C3lnUhCtu
kdSrn3BCcPZDwXWa9R9qmvwD9GEgDJFnTZJakFIhzDOo7IBXpxsUXI2qqtBioGzj/eO/20AiSiYG
NYJoUHBEQMihJs0iVaOO1n4qn00HLZ3U3MieTd3aV0ku0o0PkFetjft4oK9kW+i+16okLQQfjLbp
mHxE4vQVGdJxzvJt2393I2K3mJu3Gx6CBCZ4Lka2U7Zv27W5zuo3rAP9nlq6BrBhR1b4+aDJqLku
ps0WlTgtX2wIg0DpCfIbeJijNjmra1FGc7MX/+GWcXTWU/2SZf/xtPJAYC66PiLvvReCbXMpdDBi
uQutziOQ7nyZiCdkwLViSKby+7KfI+THIxzHmiv4qDeuy9KMPqkfVLBgEWQi7QRPP7PsSOyxHUCU
RRw+AYDSjVMZwtFQQZ6XUd7SWmIRU84wsQdhPWhs+QYoY8ULuDlyopC4c+2wXzqmfjSzlEZmU6up
n8AYDS38t7pAJbI5QH5JM2HDibKepI5inDwZ0RYLQxWJ9qTHEIFlHlRDi5zMLAw8GsdNrv4NNk4Y
cQGXFiEKuz084t1w+cuCXqOFvIwup6UoC78Vq4GqBVwC36Xf+rMeQV3nMRvC4PgZ6iy/JtE11six
MeebcclbHWy9nZY7NosvSvpLZ9WqxrJiA/mlmT3h31TAiKnq4A3r5kgYCqHR692A09PhQD9hWg/f
VONiFPcYtvdUCzrzg0ckXdgpmwP9Cw6iEhHJgoDj/d369cY5KHodBPqnNINzfWO8Jc9vLaoEt/aH
lmbbvWufrwrav1b0WsfdPspiCEzykAW8M0ZFIHSA7mnIxCI663g2yE8FZfpjiGy2P7XaJVVifbKk
Hl+Cy2rN7vZ9+JJsT9I3ToKGrKxmPL7VJXhDaykHnu/ZqO2eZZcNff1swQEvGwDHa5oVAU3z9kuL
W6UysTUV/BBB0xMOs+h/iIR8hbpwuDu/PBcLU1Mkr/YEnNukQcslRIXlHfWDXv9jNpQOwqVB/0ie
L1MFh3Qc8s069Gx6RZlwGmtsIXy4/kcZ6w3Rthb2mla2YRjqmaCTVpWBi3o5siANKk6WlUjRtZYn
/qdf8KinMGKNSNl2t5lbydM1RQ03d960rJyAP1wiBfmjFK33Zfs/JcbTJwoJwMbX/mx3NbTFrlHe
JPNe54D4AxC1Trof+I3wRpHxT5Uh81eFMiTixxj7eoaUMs8z/e3NvIHL8TV7uL5t8Dzom87t79CE
eBEDvGKDelq1+8JPUV+gfdxvaq7FySclnKgdSD8MpnTYBhTIcW6TfbY49ioHVOY3dA9IdaRVrwtl
yvjv8ftmvWmTSg6KwveZjb8BoBnjZr9Rg3D+X30ocUmpiLxEqms7ZfBVasqLXjQv4LtJhuFGHD8k
d5eJJgbL7c2to3ZKaI104bjp4Pnv4d8W/RLOaUVJfwUiG2qL9p0CoUDYWKjt5KQNeUdd7476PdDz
WxkKY7WeKqG1E1zWfwH+E7RQtRSPjqTQaXEKBry4Ri8zDHPFZ+wXA1XbyIyTeT8nNjob2dv19P1c
fzcRwomXaJLeoT0XM/4GvlJvtsY8sXf6UIXmmzlVSFQwy0HxBm2qxEeSJE5GKBF36VzTfSFsr+aD
zn5/aveb6Q+UDt0diz0bL/mwhvybH1cVZHu7ig9ue2DbNP21Rmo+EsECId0qUG7Mgj6MRsDs0QAZ
4WOlkU8kxSKHGxk/UOpvBGo3UNxQyqCw1xaIZGZpu43aLHnqRe2/ZmqwAV0q1VijX5dgOIwgYDuC
o1woKpBkgosgoY+bUm9KPwOXgfzYLGKepywAr366N+SibwTjs9RdyO2olh5uGeSsO16c4/fqMhB7
uDOsmew/UWsdwf7mXTUAg8rRlpiGp5fZqQ2/gmLXivqQ+81ri7+8FOLIIMv5EM0Nvrl4DXk9XvvZ
hWAAK5mpRUMJEhMJVLpdcC+rfGteblulpplpKJQpOQLmlaKBJNeYFniKbY6gCCRILAqAtccL1A5c
GKCNFBiJo80u43FhRxcLEbh513oH9ggfXaoYwg0+m5uFCIrTp5mTeFB6MqmOyPw7Hh36Eb78HB8M
r3ilxbN5O7AWNl7dCF2UnVRGFfwkznhNzmzLQUTcFOU54yjXMxHEgF19rmzZtOy8ZZL41O7u0jbt
2+FAvcTGMgdK7f7anKYv0MxchY5qYwxUmjd4da2U2Zx842MscLIatDcWFktz5z2csRjnKvErBef1
HqPi1d9VUaYsUynR9K/rfssVVOwOq0oJj8IpnPXImFUAzLUBhwWSTJJdcES7Kue+b1k61uFxPJtR
kjU4m1F0aB+J0XSmjMwQ7zAwqKEJZfedS9d7ubouFVG/YeqeqCcV700Dp8E78SSAXmIwKAqPzxGs
VQ+G84Ymqyqs82OFUvKBvYwSQ4d+p8tCy5ZMphJqT0lfqxu1kAqv2dK/Pe+ojSY7MvJUOactkUmM
8GNnAbdK4RXSGmCJq/nEMHzbtAiBBQIRue297XfGetW0yPgHvRuYuxhaq7+f0EfhIOgrU8H9FlSU
FdqkuKU0FIXnQgEMY54P9vX8K2NtYuXzCMbdK/M0gKavAIVWwvbe89XuA/uZweBWaRb4Uy5mZtZB
FyQekDtpuvmnq2RlRK8FXY+S+pq1Y8DshMFZH0/4jIJILAqemfJHTnctsQkDH0nmP/0zmC5zSyq0
sgtr2Q9GqBYFCEOGJMje4Aq5JdhdVrhhCSbq0K0GS5s6eTw0eHCFdjVG6Y4Z6mBnXpHI34G7tRE/
Yt4dtd3xOTBxfmWTWC4SzcivHRQGyVVGYhOYYTjKSp4YEMkZ74Y1jL5u16cb/wgMhmSBMsjiiPjC
N8WYsxxhFc1ozV+NImr3pkc/ydHSaWWJs77+U8TiiNIFxH19ZP+2p9iKioTxnYmgA5doNGdpgAaE
FpXoVV6Vfy6S18hIDQW8xlxDha05AQPEvgxbaQu98D0FJ3Pro3ZhpzOYTmDF3ypDlB5XyLqeXW27
gpmC79rX+WuAWuwIR+Hd1P0zg0wF9ZRrE6llQCsDQmnArQre/xm8HTGU4/Mz/nR3NfTIxh/oYg96
a4/VLQF74Gp6/BS8dHeQdHhE34qTQQvq1BlysyBdaSsHfUMZNZjXra0pXVpDh5omZlhTlKssEbXh
rqdQR7XDTxI0RdqlAVDu8D4kd8E0tuWmkiy2Jp7IRPtHLBQJnOLedgQJIT706hs26uOn5CPPI32M
pOa2pxEH6/b5lrYdrVE3mFboMyRS+hdRRCmtv4TblC52hTM5PuR/Z5QHzxCT/9+14hIAD0+KW+Zj
Gn+Vri6Og+bE3bm7doDCuxiETjRq2gnUAtKKAtKZOeLLxHS1vwlkFZF1xni3LfSaO8Iits4oJD6V
XE3m08UVBylGmE9YZf39cD/i8+uHGTvqljjyzWwvqVkxRmG2Exv3gMFBNQspdWadsfB7ip5vpFXh
e3igkpj1umOPL3KoFX/I0hdDDcUAl7MI0YG+E2UUmID/efEaXVhKL61kl+Xm8V8A09xe/fJtMVqs
qy3hU1k5KZq3paIAkgI/SbVGJBM6V4YXZ+5Uyn2oMm87iOdEYNmIwgvFnYI8z6IHpWbCntZRU2ve
gLIoHekkNaIoDtPXmOkZbJjobROpjH8n18JOCzhXUPDwHtAS6DVZAXNQA/R0LojMi2nPR7qSdCDJ
93OR2Qs5YHbk4gpVI6TNORsYE7Mt0KT2UrPmboABMgj+5KEGDXVPLotoRlYfXw5jsmaPSWExtL7m
73aSsPVFxoRX5mKXp91bAFCuWCeB08G8RmPpthAwk+59kWoW6ce0bWLarwB4WGAcCnZzPu9ujlz8
SgKPUkPsHFJMwBm4a+OZNQGksEDXKkoSJmcElX6u/EyKWt945OcA3sckYwWazh9aX58jGQfDR8OD
qDKM+hMvC3isFVifaOpzCnJ2VQavKc5T0DaapwJGrieoL2TgxH5b49DdZBOsKEl1jitTiZEq0jUV
EQE/jXBdYwVJurn7zvAmTxBrhK8sztzAmic8dzIO4sYSlz0JFXWRRTVmJPbxrQe6UjwDIWXxvORD
A1dsLjbunyLOJRw9TiHxoo5pWfRIKeebtzQ6na/PrMYVemgLEpkFHkfYlThLuIMIAfBzck8NqS6I
Iba1qx/ANm+jCubzmRccMrJ/opBWwZ1Ms0AzjB4OFD2BHWXYZhsEO2rk0SQ3N4CEWlAAavtC6Mxg
I2DxXUoeYmJLoy7MFKF2TWxrfoNbruqrMSKZzB7tSMLVcB4MSp9ySk3Vtko3F0lDEwi76KQ2SGHg
MoM4ZJ1LbUzVsGYbz6yYFP8BRq9jc8B7HalQHBIJ2XnxreMM0A8EsYd/KgQ6dDn0Hjy3fq1ATQ2C
vbvQJ/oK+Ehf5ELC0M4DOmspZrlQYtZyvvdZHk3wkEgdotUq3SvMV5rMLB1wqFxVg1G5sGFmzgQZ
lJQBVLdQI87vTlHUCN9u4pP+ufD8JJW5qVFnSzODzp/6OCksKUN8n3EiYe8zWZQvkrk/kO8TB58a
PNIz+ZwBekzSpPBbXXS8ZWMtrKW+4i1DGUJrHAnaqLHsUqFCoiYXfBBnVcP5KeIYxukBVoTpn+Rg
ZzXn+Jfhc6y8a2YuuPHny22SdTbXzys5FkU25KFSk80/Rzj3WIA4iGLeWKZDtRGmtpPo67gvnOvL
qSp1nULhBSZ6rXzhfJg1faKf1N3pLnsyyoirvF0EzL+2Yg2hFn9Knn2nzyzsUy3WGRDCk/1wmBRn
QYCiehZh+l2S9g3d+vqu4EKnt3/ZybFjPmtFKH4uD6OMbDYVgDkRFDCtD/YSFrKrumP7O6bI3xEa
/2ZE8fyRGforZ6b1Abp1+8bKA3U/RhBUr7UYj7KTPQwNN5FY/KZL7jusKDjgeKq2rJChZ6AuiEJz
kFdPOm0CkpqWnXNJgHAy5A4Xoj4qv9lYyYFciW0IACs4YayHC3B56eY6m7qHiFoSJgaQJOV6Wf1m
acd+KJtJKTKePXggMNaqf5MxiILi/fCBuH7HJIm2b5C91LyDGqaSjI6CjPKNBXN9k764SzoxRc3Z
C7THraNqPagcAiXTi3sZAoIDvNVNkj/eI8B3OiBXuHUM46IyjabcA9cvA5FyFvRKwTIe5rl4bl6q
d1G/qDuaraa/RD2dYmiTQHZ3s+VvCC9SXjKI9wA4K4YoOLnwDNRd8wF1vvNMuuTV+PGtDiDtahGo
cckSXNxpQkkDaQ1lf9Q6ecXXtlYhUsbVY2On8TQumYYSMsmaHZ3tXg+AtCc/fjyzcM0EaQXTsGUW
D6DRYWHljHGIfe4LoSWumeto+JOhVyRfF1qYQfnmTthXfai1uVnTbLTaWpgwGiyrWR0CFTbm5qVf
XETQDPYxX3uFg1mOvUMPsF/ujcqyFp4au5mlL/qIXWfqIpJiHo4lz7hXdn58OeTF29dBmzxrCPmN
Wek1LmWc911AxzSB+GgPfC52P75mWP7RFVaHKlvfDodzllOM3yDe4rDN2scFCZckL4VW5TXwCF82
MVW8Prn+hKO17bk5McNWeqe6DLDF5PgmLZp144pLWExiJneHhFWh7v0ZSpMv6TxmvlQQkboBjHET
bPYn2CxTmtUg5ebYU/N3d0VXIs3roEdnPvXBqwzBxXXloEfAddg7vpuUjdlYcpCI+3WfQQuPXmTB
vP09GHDANmqsBg8mgVZ7cm60TfhKu7eG1F5T/Ykdxy89RXDr3NlOqvhJFVmV2f2yI/lIKhzN13CT
4lJRby+8rWDEnKtRtuyO49vtc3h6N9gAjzCFH9F9fBSDZPA7pEfmTI6W3/bQOJOKl2Q0xocKjuZ4
F4Z6eGyDXv86IDt20fQCTU5fYCQn2PdnQMKxT/smU62u6R3WdbkNMwnGGSxKVQdNACNwOAmhA38k
WYdAxJ7MuODacFlH87O6u5lbmUkMA1mLM3dOiwZeHYiSdhxHdmBVuFQ5eNzfzaDNKnaPfAV1np7K
LFORFDugYrnvnrNqO8JCoRMr38RcfB7A+W16hqxMmVDATiLHqpnU2VpMZz1YIfbDGLn6cfDpxq27
sbbt8hPkg208PUZp/maQVBV+esEwSlCLCNTlYvtiCLabwjnw6eZYkdpD4oxnAEE3d4tfEKUoW70X
0JDc9e3CmJjW9v0PhLeYUUKgtN+47qSYU1qmhAZIdqYlsOedu1DBaNZtsLwPj0yHsTBo4uKS9sn7
APn7N+3HX+caXhT/sLNjdF+/WVIF/p/8sX+4UJmAfATnXuGzri2n9XuMAhxvz0rxSDmR2IqhdXkv
iWzyXHvNc6M1AqN2ngsPsDbWI6vAOQqGVlrEZp2OzlPVQ/KUoM2uZxV6VcGnI798BnYx3NChzdzl
ygyZn8vhrSKO8+Db3eDDXsECkMahT2PrOTToe3buUD0YnsbH7it7HpDBdtV8G7kE+z9bBNhsM3gv
ymKNmberV3Fo5yAqzs1cee6Z7YEe5YcG6Yhkbr0R0pxuYX5oyVgErwaA9uTwA2EKFo4CxSmzcwS9
Md2QRPhuyJ/SnDS/ltIj9mV6a13xnKss4rIeBaBmmBO7mBXnFjNIDFeCyALNQhNTUueRTi2afAe0
y9eSIrt/IakxyPGXUV7zYHI4J3sorRmtMC5C2+Y9hxDO95EIyGitY1oMxK6/HQapVWmxFveCbuNN
PEZImSgJCDgY30lizTPnTd5IpOO+n+ySzyjM76QqIvgLkKG76VZ8zenTXiSC8/N4+LijwrTS2Cy7
LuADegdgRq2uyLdU4+REXWrE9A5LmPIfKfPQlmXpLBNUDcU3dR1Xj+iB+qmuVD2NY+ZfJnBwDEW+
tZXH+X7i7CoIaueE5+o1CqjCl05S1XXJQjbJVnj9e4v/AXxc82h70z2+APEb+rSvFKa3nvbXWeHT
m05C9+CFEXEGsccipmgisrzidgLKBuGTPT05WLZsNYr3HcR2NZmQsA1zgPggTl8YUnGEOCuZ5VWW
8oRJ0rnUPD3GbBy30EGDiX7WBV6LDjFUeapQbwNTTNtSYZ9Nb0I527f7fGtXO18iKy2GzX2ObMEK
sEoNgm+mDkPTl9EQ+fp/+vuKVxSQFtSgMD6Bqak9573yATKGxxE2fTyOaJINTye9C/qtyIReSo1H
kljQaZxPeTQFii3aytqwiKpee0XXj0XKCE6sdc+QVT/RVxx7C7uUzMGF1G6vEnKRb0QBsWT7YUmh
mgBAR1yHrwwFpWsKB44pSM0GL+catDOXgRdgA30ZrIPeox9XLfHCQ9QDXX1WQzoSdWCEM6qWfiyG
RYN6PWQG/PPppqJwI9dZGtN0KFGI0+/PoVIrxxNk4q44pNRWP98X1ewVbmdyAnPF3GC+7Iu79/SP
xXXele3dxhRx0eUWU+Ic9GiRfXFau8hPEShGV37YvTvoi/DXusURSaL+PN1RpNujlb5ZvCCcyi9k
7vKEvz+XOGvEt6h8oVUQJYz3BGxHpI5cAM5WqYLKXuaUCgDpgrLrNkd43jyuXykt9zup+M45tKMk
tK20EwL9BoO5uaccqsQDzYAiqo+TN1SvdL1mH7FlDXSHZuzPe8LckNZCoENonIpmdFWGSUrEXeDL
RxFPUrHDv5hUI7d4XyPmTrqeGfyaBjCcWTw/FCuSiXKWERCviynyitJYct6HzJbvYDFmO71yGPM1
W72yjLIzUek8OncGMZXYzI5pYRNrhAjLBkWTSKnGAgNfF8c8b2wy3oE3xzjb8ZamYc/5fyaSC4KH
MJnKQ5Mgf+xN2m7xksajm2eMqSlnzuvidquhlOROjmgZbVHqyl9SOU3xRc0HxDXGTZDCwuusuBPZ
du4grneLuRbs4mnI6Vtqk618pNgFcBGd9cJtrjZradhRD29na9i8U07bNzs2y74gtGsUEeHtNC20
xDagpYXpj8CoX1Ym3oNhnzRjkEhZsCHRfZ36ZPjwfcQ7Pyd4VBw5GxMMTi3tCza9IGTv3C/Tok7x
3k6JPK4/+STEVz51DHlIV2m5bfNbVSCvEqrrxadKBufcfVdSQHIqwkCVdgF6yNVkZ4A4XZvsPeJX
OBIr5sJU932V75LrqNNUHSOtFamtLS8IOFD6kDc7omZYNGJc1JEkIrYZ+92gV3uTr7OHuxpJiOim
Uh/Tm/CQtuYzMz9fioYZ4IA7QicG+Dk7kRDMqGVJB+rGeAM+bqxTqC8DoV0UScC5htBj3l2gQi8k
xRweth/iEuZigwBikGFp/WGGIDhB+9i54zDBKFpbvrzWGj5dB/IdVm5Tbii6Kmstv5PUSnI7Ic6D
yB9x+dRPkIkQUXhUuW/HH8C7D+Q4Zy8BhfdomCgQNlr/LWfXrS7pIelmaUEAX1L7jU0X6Z8tQZMR
51w2+Rjzbj2V8DIYfTbhzWQy1qmWW5gFrhRPrCgjdokhow2JaNnZ3/zGhzG4g5uh9tnMrL909vIj
Fg3a/jewSwHjhfhuNjXI2NO2ZjVByrZ+M1OOzjkHwNyz2vcvWGZTk5S9xQBU80jSP2jK8kx7njf9
oqtZECZF6H8lcGwTNZZ6HKt0jfQJSWw8ARtfD5MAwIIUtJujQp6Q5iiuSPHaNY4MBik+Eyktshry
ED5qp7sOM2F4VsudWaKEiJ3UFg+M63k5mGRM82s4Pfeedi8gO0+xJZIigL3NgOo7iZ0ca1kILSdV
BSvF2okslwJ7qcBtTxqEygvItlD8KwGZ5EwaLQP+N+dxLqddXrHgfNiUV88rSQ9zaQljurS8Aa+3
8EPEq6VzwH17Uw5mRvr00vZClCzDvTd8F5RCO89dbidcdt8fVfD7yY9Ft5WqH2vQbp0sbED3i5dq
lsFp/ePAFWCydOMnZ9IwKhYRVZ1Bbt+Sx+LqU0q6QWRAUZD1Pcutc5RwSTk2AbomrLQUPKUjGC+2
rvo6JkUejZxw/yPTBVokekTRmVpik2sKgAiJl9n4ZaPyC8Txt1j0pg8vxRnKMEutpfzDk21OQbGr
PqpmH3M9yno6t35ZpNCsKWy8mPZg6+tyAWGVN2NrgAa8Hcd0amEHBQUPdpy+nPqXulKS0Diw6vPo
5KOpLZeUVVQcFzwDUcHIckk1CfufL71zd3yHRFGcLjmR5mrS27AKVBPAU5ITxEwgUgHZ2AZtKC/o
9156qaIR6CpCWdiKmES/uA9ocEqrfD+SG4LaPR3Bm1J8VuVaBRDkSthewhJDvHVI2QOdHojkcfHJ
JD8HorfLdB+eAGgA5BEP2oFoP1sspSoz4hi67kUKscXIaRQelnwAJI61cdE602zLoCmAJZJsafc/
vqHurXIE9uJxFjHSaOCh7DwwaC8CIhzNw20pxoqSa9Z4aemaqxnd++ElstTddZQhXLIiWISp6ntB
Y16+tCl3gtqssq7LkYAOUXSqn3n4uYDcOXLKV+Q7es5e4QBqZ35Z3ET18pidKy/OJnR3ti0PCfFD
xVZkZU9QHJDHqCKiDLYiU5GbT9PM38LPBdECllwU2Xk2pca3SqU6Y6x52KFQNw9RelsX/NftJXNN
6Gz/QJ/vA+caMYkBkLnhJzrmsFhgO3H5LIz6NesfIJ8vDiPlenkWXAo1mfY3gnaILwK26MP+idPB
isgCzwGhST75Ja8NgvV7P3y753Ll5egxy2X/iIhKpCnXy6BXA2aL4DDuMPuluWEQVDy6Cb6deR8A
g97XbDTQhE8xvA58id6GkPwxGvAlR7RUIhPRb0X/2xMEmaUPjyNVEyY3gZLxun14RyhLZwLtH8DU
Ll39XK9TBEabL5iOc0bVfKS2k19XT2i4U26h7l+pJzj85Ti7WKHEWWSECdMcS3OaZPC5rBqbGYhJ
1/XnY43DTaD2a4OfLvFAGBrA85n8BYgDmqF/S8Lf0Vcqj39uoj4cSJ7R85Pf3X2Ch1A7QSnHcyND
W/MRBxf4C7zvozJC8U2q9cT4jeH442LKxvVHV1wupADgxavt+BWV5Qxo3etWh3G8dSIlsdsvOVpi
rmYxAShOF3JAyRp+MZGqI7PWj1v4hdyavWES+wWrdCTo/e+4AuBTe4OFAeq6JuAYz3b9J/fqMlaL
0MtHjIu4t2QR6E0MGzaFbtDO+RAcbStudW5CcoHs/u3y5nrpUCz/9ZeNZVslc1NSGUncpaAha5Y5
N6C1+WFHgxBsIQKmAHug+kEMgJjbpM/EYJyTt+UP2IOGRg4B73ICcBVNZUc3XkO6DotziyiSi2hH
cRxL6KGgXpcJ+V8xp26hpqQOUZ9V/ZkeoYVEr3TSG4PZhEWgV8r8BQwnmYdQNrzj+rJ70UfF1K1b
jXDfjbZkPazW/lqTvfQ3lFMvIxhpg9EQqXFPUriGPDc+TvrDQp5hIS2d9nqs9A4jheA/C08fB8fy
omKIdwYJZaJ1KW3NXijhNO5IcivJBY6543bMz3rZGjSwuycaegaXoFT4XTQrpAx/FfP9V1H7aM6r
SZmkCt8dckWWoipET5CJZC4NOapv806DqCNLSirMfzB96aTWhi/aXJLVz3W2ROZ7nsC8lFVLrO9M
OFfymtAzMGL0kyX+UgOapm8DaXHvQcrKF2IIvt6TVjEMtzHEYTsaypyC50q8w62ldaaPWSrdo8//
tDKb7XDXP91Uw1LgBFPHf5piaWXC1Xs0KGfS3qGRkl9WuKcJ7i45y0obJXQYARCOkQwhwj53tldo
I64ZM5MAC1/r1pVeKiyKvS6NURCT4LdZsxSF2qIAp6oXM1KYOzlv+kMng4+ZUkR9WiIEln4+eaVZ
cBgMQakQFX/tcmlSHKYKoOy5BUakryVBnRWfs44iQxluqPGtL889mljceSn9dl5oE92MzCQKg8Nt
S8jVY54ko6nRox3ptHS+tX99e0evxaU9EyrQ5gD0Uyzg7yTaHTO4EDgESqRP7obgN4jTs6RMxHtR
JEaAJ7301UtrhlFVXoVQahMMu9pT4+ZkMrxbNKr7iq8oHCecVeTheZOvTBtgH5SajCjmc/Pnsemy
RUeYKV7Uh3YmfMICCg6gXp2eQm+OW345x0efcG7gVVSo2LpmHxOCBY4kKl/4TryEIMeQKTG/c99w
cmflMtPdIrZpmW/h9m5+/CXYJPWAt8NnF/1OQ7bbKWCa862gxx5txy6eV8QHWX3fa1FqufOULkfD
5SPCVRfltUOJou8dltgDwH/kahWqytLGMVdsRyb5/dFrqm/VI8OpP0PHhHIwTlrVjZBUIptvboJF
2hi9yl2oyaBG/Jl83YsgFV2ZcNqpl+6lea5QDRSsywXZFfeCgQWxLvjApcCfkW/Yzf8RWugIXwF8
+n029miH69dittKKcGCWTIGgDPtWbhUsSYikJIGJGvK9bPuh0/U7Q86WbNuBqZfwxtgRe2dl8VA8
AZO9S/8tCadcryqzIl4HJzFwS8Svgxtu8lLBJkX8t+/u6FtSVwPEun4SK+OC8cscFK90S9Xc3aPe
9n94zzbyvYDA01SSnL4yyXxl7RTfmWOINm1nNNbu9qtGhfpyZrRtcQrs0yr35+IaFXOSHT5B56ZB
Kul2Niw2Km4ghtbMF9EV/43Qe0DP+2DMp4KaheUH1fj6e/bus3IcEMJfVSYeezDdjHaAeYk4JKFW
AwKIAPl4v+OGevrk5BEj2+0+9PWKqNebGHvn2vn1esyXN3rBVQWwwsZIsLHTHzfc10XXa90qVLFe
ffZBnD0nCl5fPFozjHxTIVJYgnOyig2067DfKfSpiW2NTPlgOn3k6RUF29E/Kfji5haoJ4bI3fG2
O+xJUmzhKiwcI3+q+Pluyi914rWdhmPHoIyDSJS9CrGgsmUCPdbp+3Gz+tAg7vW1GYsn8nyIeX21
cpnsWCwL0Kzg9+g4zRYj8fLViB8hHh3MMcGOM57MPmyYirF47aOR+9Gv+fPbV4EWx81k6HQFV7rO
3Ex+M/6I8vsICJY54HOFtmN6pznWX0rQ14GhNKzUCohIclxw6ApFZ57AluBe8YGfRDlVFLjmnf0A
Ej7+z1rF3IriM74ZTIkWxzQEGMNlsogZe5QUhuI/yQPCUcfYRHr9U4Xy1j93caVtlM00I+/x6t3f
FjjcfSs2uNhIgUSQimzbO6VGeld64bw2Anv2ibHcf4dGY7xBVOsFG5c77XCezYQcTnNbreqAMngR
2oPYOrtCTZaoMd5snFPMvlZ46i1ln+GyQjU08sBE7gHw+fnWTjfzo2EZBR9YiX+m5egqG2Q9UE4Y
OB2iFe7IxxolNgBfCaddDsCJhpKVSorJaCUezc9QJB55h0A6jg41wwM63OyEWCqVK0u1/ghXd0Qb
rk7h+afmlyumKy8XyZsVWy5e6Jd2PsvmInjvChE4eSVcaGxgTg25oSF5+b23i0cb5Q2kiKAYjvno
P7/hLs/wR+sp8OJwDK+1QhmtmX/zBWIPcdZthS47xs5Sw8Iy7QTWVPA4ABX6J6hlHwh6riW6HDuj
e/fI++xpVXcR1/ZdQ9ahgUfv2QO7uboUwKCW0SjXdCAbZcBXcByuXidNdtIIVxzocIA4Pum3Owrc
OcHfeRn+QlQ8lBy+JISJjU/69e2kSpvAX/a1BDZ1hvh0iYR/PSVnqUX4di0YbhvqPFwAIk9jcdrz
zMIWD5PlbdZK/qVSbLVX2oIY/7EIeTYRVfk8Z/+hJT2TwxWyyQiajEjeKky2ape7qVcOAsHyMZ41
UG9y/noGo1am7FC5VZYz1D1fF39StG3mqDyoTmZ09u4KUJr0MPQn1FMx5yrRydhgN73uExmDjI2w
AnqwfX9ZBUKyOFs4IhvIP9K8snONCUj8IOQRtahkp9zHwA5iHCk8AhxlRZBH2KrVu9r1c4os5uu0
VPnqtjLmHoO0kNJWVQMpaJtU1T/M9AnnZ/m7PTpvnP9CLFjbHXlXytC5uJPqzxanTzV5DoxADqFz
N19fY8ct0wnPJedFQzVEC3JIs9MIEinROAFqtpEYKRofSt5olHSYKqQRwcGeVQG4zBdnOeNjgXHV
wKMwORu7mAiI0w/ynA8RCBVf/KJcvJA5VfdZrK9bYNF2VFs2GhM81HgK6rFFaLhG7TunPHCy1vPD
dRaHSviBpkzGhKCqSyQIzInDPK4JIVUGSgK2pPDP6rsrxAn6jwKdO7Gr+I+OkjGoDqwuaCzCSlJb
3wSbb92bnEDC4OTDYevDFTnRwqDm4Ton9WqYwWqYHnnxzwKsRIb2/q6ZEtnYqHtojQ7egiHX0rV3
jPLtOgI/upQ9aRCLwfbBhX/uXQWYFmJGMozxDLNXPgOdOU6qR3+9hFPnbxXK3B/SvBX3+TiQrW+1
Dai2eRnTDqQ6MDooUSbe+ycR/Von42lvrTLepdw3hj2/vL8Y6C3PqYkw21DL1E4QYmCf7uX7/cNA
5wuUj2Qn/a4LQUITYtphtlnj2xwSxf0D26PoDB3V3KxCVzLmD6v+Whse4gyl1/BCSqJ+qHJkO2u8
d+oa3PsTF0xlpl6kxnuR4Yp+pEL0AM3Q13xmdytLFtBxC7VbK3kMqqUZPzJCZEPn3zBtw5fIlbn1
1/eYF3GvfX781wbQt0mOoDipUwZu5gCJ7LM7eeWxEOOGiNY9yrMT6ffwM++71xdYcmDYSWtl0wkg
+xnYfHzb1ygVFS2HE8Q2GA8NjMWqs1aGFrENUIfHglugX/0BSwIIJjYeexGnVceDcuuT8WNVdr1t
VQ5IwKHC4r6kAd6VmyBnlMKAawHYocxUUDTIXx0TyybEh1X3Lj5ywK5vmoHfduOBFMqj7QpVu02f
qxEdZI+CF7p8rpog4bvXUMonnxzHZP1HSm221k/aeMLCrX7Uv4Pl6/TyGSuKz10KIhhHJsNyCDQx
aan6r76wUFXUUlfvGTq4r51eCQ1XVDZDQYgaSwujOP2BBgFI69YKlrihLfczh+EEmlzCk1EynjDM
YFTz6BLh3C3TW31oBhqni9PKM1jgShF16tXxfEUAclU5dcJ+zyZO1Q+GlovRj1pdgdHLn1NnzrpB
Zz5PqW9rvQYeMBYFcRwLCo5XCTBdKGhb5a+vwbpPqcHGJgkji8pNl0wsO4qQx7zhAZUdBJ5LDg7R
smj4A0a6Yji7EYGVUyG58DNweFcvD7EHuDJ7fId3uY2t5q/sPhLW7fLCPAXsE/Q6J9ZXxKKRLRkS
xpEeCwkJfRXRHhFXDsOcavdu/xBFWKoy4p8LTJ/3773SgBZFBgOTHsMNvsQ7BMXEj/ZWc3qPMNCB
SoQ1lGtrI3WHaP2leilCsgGdINTikiOPjgNbtyRheYlJZ+3ubzykTaotueW3gONq2iq9Z5wOztwn
snexDMBGKD7VpghDQGygYhyoEgV05sN5vGXd8VfPxi3r8/bdvn1k2LVSTpU0GVI0l+eFcRPY5qA9
FEgk9GcFPSJrF29cJr/gcAQMjvK20uaRfGRLlNC1TainurLp6xwMYW46I+mqb47fZGBsG+4cfX9v
y3ce1mXD6f48n+06AB4lIemV0OmgyPWx/1QNdECcVBg3unUMOw+HpASrjkf0khsZGPm/QxTGmVB1
GA23jgICB8qTToGb8GP1QidTowv0jFlmuCShwoBH0S36sDFFQXbveDCzK8iGq+UTWhQOwKRIIQjJ
7Ej4Fu2XO1N5qATbKUkWfLzZ5ZTpaWSWCjV8O5ha8TObyMsj+zswNgXOyCkt7sFYUIdqIvVIxIxe
+hiKekROqVc5c6qwMJOdl/tjEZgwSdB81W4IYeLx62cm3BZ0xskDS+ftEkgSE8rvxZO/GRdTJUi2
CwM6ISpN1lsUJD+Qq42wsFO0AJPsQ2GSbt/StnTlLMpIxfBTlR/m00KhbxfgzjYGr15lHVXUXhlP
m4yyKGnOIV8K3sQgux8n4pQqqZZpjU65F3gYOGbW0nmSCvWUB2TzdBvZ5hfMu0xYk2HkdpUcYFT2
agdHDGFJ9Ao316XO5TkJb82zlJkxEDK//QW/fWzht68cAKaN9pow9rmy3B8fklDrKShl1ccbCp8X
0xYafl92k/tMk2kAnhWylkC/+t6z0SaGACmA9kt9cOTpc3VAve5xU4TQ2oviUpSVgiLhd4YPxV7Q
QlglyUppsoeSnL5A8y1q+eqR25emyvOhjuWh+mjQqoIbiXHnG/RUl3Ds0qCXggacTOoDVlSIfgHL
xT91QhwrMdwrzh0IXmXrqHP/w8KKKXcmEFttE8UWiaFZI6Na+y+Y3ztrWMBud84nv9e8an1KUvbw
lJunhVcxNnlzXlArUdJpB+ER40tyFQsBcKimDp6ZG7KCNPeayDKszsqYnJEsEi9GhHCk00QCQQ1c
EN/5YHJZNt6eniRJlxR9XQYgWywYY7U7symcRCQy1dr4DuziBA7K1TSergGNanKE83QWm4WRITuj
ER1/oAnITN7B+/7gSggotkw01vZyIJsoT5Vmvb07OnmnfGqvDwAaoDdffqw31YySyAYOABR5A83u
nJu2ARkdrJlXWgGSqfA0e3xUo2y/GXE/dMvD5MKPs8NO2ARspefwFDNn4pd4KBTisIb2CWhZFWtr
7Nhzrw+p+0er88M5Y9Lr0W3004hCvulQMV0My7ym/w59/b7HTRkW9dLQnLLSBPEd/7R4j7ZK8rmm
GInoPJ6W3neqmsGMyAy7iU0dU3i8jmXWi7wDcU6t04A1yJ1AyK9UJypDL70GH85fARY4PuG15UID
Xzrexca38XkaGCBmYaqdO9KoEFzrgoMrUDn4mzfimDwEQ49bdyXqRMferITCLODKTSffSRkd7wa8
Mn5jSS73V3gYUh2k1guKisvJt/tyycrybt75Lc/tjBYRDS4Iv11an3M0e3WCuzgocP+uK2vocG1D
4CSPSmY1g7kvsIyKoX7zi0OAfvir1AYW1xfNRnuRR8DqVAYiEJnD7WH3s3z/aGmmRcmyff6376vT
9KkdwduBzKLmsxq4RzJMLA4YTSFsn6L3R5pb6C1xoqsk4UPC6vxpL9obwLFttPoQbhYVDsOGXXb4
1z8PYbhLgPe4QHEPR0ozDm9kBRXVPYppQGHlnb8YLMiU6dIynFK5a0X9KWeVwf34hgcParmCrfN1
v3MnUkB0rnFf2CnSPToDje0DX7pMUJWuoAIJbveweVJXafjuMq+5BXWOI1G/3Roxtkg4cqrnFbnF
gpWUdQZqXeuJHURCW0lgjvqNUY13rW4r6TsFDZor3o7+qgEC0o/RP4wkdvbCbsFDfPjbGjJdKdfB
uOTb4rw7irQDEqxoCawU1cxn7WwEdlPlGkK63y7Y8nGEUBu0P3xUB3cf3oCQy+ie3To09TsYB6HN
0EvitpUw4TlQy/tKOeXKhoyWow6e4ZjJXaBJND37GJfOxkvPwP/1BD0O3WKIDUvn/bcr9yEPl612
rQKatxi49a/H4SuO8obald+TUJ1YfANUlTIkIX0UtrDXxv9VBZj/atlaTFEWzCRtUKxDdiZZuwPX
gCTbPwxgQ2/2Um64z7GAulOtgMCTpcn8sGUs8U495r6KNpyf/FXXvbQx7xdqXmoQdVcRMapoU+ec
tpxyqS+GXHg9NIB65ocPPdYzncDlpWTSBzRqIvYz9Opaxw+35N6Zgm0hJCUTMyLgpDjJI9oiW4tx
oTZDtw7a9a57yX4lbM6ExLQdV7o4qKkj0/8GiDma6tjEJjoKUkSCXnTKdXuBwDssV7OpI9jfcVmM
sjtrtURVlSPGcN84Yrxwxox6LbrHzff4XOE/Pbh56UYganoUK8PIb4RcY8PLEu4LUiG8t1HaMBVm
goWryqh57oxvqJkjoKOJp6ilEZV18A6u8+b8B32L3shspTz0Mw2GD2BCHWZ9ubHFTIbraYa9iv1t
PqRn8Qx7B003+LeUMQLymn9AO8Jdj0fHs1OjfqCYME93mP/gJMPOkaEI2tYc/8hLV7vN0LHxa6Ga
hrlkqvxYVfGKF7riw2EYmysslct0JfeimesgihwVLHtpZg1so0RmUYO90jeTpzwlT5FmL0XYWIVg
DL58CQuugbdp9ybRi2ZLRIXBSYiiAlZY6YTjlN3IhYHJDRYcw/nmPWR0FGPlyWzdPwoWH5Se1XrS
tvcltSVxj/vSXZ+csgH4wT+hKZNokWTYwpVohhcA9cYpvZvBoIgJ4cE1FdmPLKkMs3I1AyH3ieW+
MPe74PJVWxRFpVX243aWiHQmj3lQE9nxMTunYs+sDwCvF0oOhqfRSafey1B4ZX2Z5llI38KK5q8X
VqSErAzQTN50J0HJzv6AHy2pbjVfl0S8VzrFryYjrk7BkWx9GX1NPrT/gy3vfSin1iSm2bXLob0O
vYY91r8u0aX1cCuA2BhecRmScBkvr5y3n3ZDDjrHE72B50UlYOCn0+pZBSg9AYZy+lYVNy8b/53p
V4ThhnaQT2gHHkl3amRQrE7f1CWPQUp3Sv4kqRE4Il6mri7chQ6XlZXrjfo8jr801R0Dc0oTiHOX
Rs7KxI5fp/nYCz2G4AIlhKl7ShSZI3RGb062KBQoOvbkEErKLHWFcnAaDxc/Npum9wAjxQS9YNGV
/rgdKTsYYFog/mZejlwntj8xwQJ22WJquyEqhNvmt404WRK+3MpFJQv2zybtm0AYvud0sjhs6j69
soF2KO5ksVZF8QSJGfJs49vsr8Okq5Kb5J00ZXAobvAZao70v+z5LkZBzdUQ/j7oRPOsRgkG9Scd
vkkfzgyGBELNf+pn8VeTEbqMXkgkMwG8xMso7QLA6Tw8b4WK8EvV83CeSC01h/lVHUSHkrkdlu4o
JEguGfo0AtFxxS/MdDxK5TEf3+gLdfUwezV5m/6Ln2XceIdCiReWPqowA7JlkVU0YOUHNh4Om7Gh
4SOUXy2TCpvkN/pib0h6UBkhV7G6gbX5a/T2avI3t3qEuNtj55iaw4R0Cj8jIQi78gNaD0iCPfoB
J13zVEb/MQBdoRdvQ5pqoR6/gHoC9jF/Ddskm8asFxhQHd9WV83kRbLzAzfIWRDTP6vXKNZgI5DQ
daTNl6yNNLlIHQoMv8/CU7Re7MJfPhHeMDe7lTXzo69PYaF3Ovbbxmj+05/MRaDsUoS3SCPL8IYw
z14U74KRmgL0Syt0GGQmghgqznSUtqRb007jQq/22btEZhy6X+lLU8dELAKwryxVG65vJEYtdlup
OaR7WJLGlkFtSEGaCwHCMa9Sy9NKA3EgcFxVFaWkkon2HGvi70pzH9JynYqXMD9cM98q72hcKFQ3
EPAqUPv+Z3swAIpDNAK6LBwVaoMlIIaN4ET4wC89Mz4VruFtH+xhBRDX7f7qLfYEzvrUgF7pct7K
S6vq3uBnolVAFfzHvOuusCRFZ1F2K08KGLoMuMXcGIf/NFtA9g226m7BGbe5pAvTPUr4RuDdJJp0
gNRGSlgJFGmWduqu0sRAu70/y84o009zTNwrQw5oSbaeIFZVvAE1kk/hCM3JcNOLyUQxB3duE2yR
+keEGavojtdfT4eACgPo7rjNHiODovQdZl2NeldVk+WE8j5dkwq8X3g9MwnNuyVgAo1A0MQ71tw/
qw24zptC10vViOEslrGwfW9jlE9Ct+iPrhzPGGzHUUgW1hrtJxRKoTvcyaINdbnCchkbdfLNO+Rj
ubu7q7WA+HTGXK00+s8SjYOga7RE/uttLQPkSZtqyYLjzlJNLAUMHKRh5xodOXieCGU8KPennztL
RvOe5DwLNnjiSRsnNBZlbRJRGd2ZkdRy3j8njZbqOb+4nCUvQN25Rl405rgV+H/59cG1NlmCym4r
FtjktnXDjMgZQFp/+hNKEI6G3IgNhJzqTI45B+M459xGMgHyHIDQp2M+xlJrKyGQk2ElBKmXM4fY
5TTnfHgMY6Fe3AABYgq5PiLuDWaxzL02z/oTeTeJ+7SYvHjxFb6t52pf3i30Ax/nWLpymWrcP8US
6u7e0TgRnwMPK9EvoWEFkCcl7wdikTtk+7vGuzY+qXQ9Row78CaROc0iYU2h4YQGStpD0LScb6sE
oWBbw7wcgscyyRzPtTnXzU746JqfPywE9AyHw1TMCk8l1XDLmDGqQAqJV7+0rwqjaS4CljjPXJDe
Qzr/1fbP+BCrwV4TSHYUD4J8EXbjJLDQTLmBr0Qjqpa57YlDq5IUAb19QahqLuPxF/9dyXBLYsIr
C1Eokeo9Moj6S7hs+t4ChwsYmAPeae6mjCJOFkf5z9uC37wKey2k7I3KHqYv6B02RXX3U7qUxbT8
3zokhNHep9CMhrEXp4nvPJnhKoAA4cplRwPesvnvD40aYrw9XqZ9fIbBgFvpcDWDZW0iW6oTm6zQ
VUtiDSQwNkxlWVPyRBTsNCp52b7wLF4P/hdRhturjoRRwydD/OxBX4F00OVR0LV0+Pd+cMkkgZP9
1Jp11T1jGiy+iTp2XITpTYmGA2G1tGPkEGHu/XGEaJjnEUL+qvm6wxZVDL4TO/KZcJIcXbCZLM41
T8sUEeMmqCsUffr80NlQrGZB9QH5zGpaE9vT2UJCZ9WYshmkQmN5S3yPHE3eXW2L/gXtzCpblMnp
fvhKUG8XRPQiVJMZ1yQATGI1r5tPkc5n2xfZP1aBUngHvF1VtkTjcD5Dhy/uR1Bl8YkEtp9NQpAp
I9jfmszSnsQaQcmAFX/Hx8/+lek3P8rmO0rOcHb+AhwuFhynZTbNc+LvyTc8g/XfPd5BZrUQEdHq
X4Ma4xc+s873Voql0Yy5kIldjuqzjK3IeyMWYsTU9842vrDB506htrzjyAjR+pKNSWJbM02wFERc
HIgnMx49uoorSnGNxXRA1FKQBbIJTsiHN0MNdIYK4sZczGbxo42ISfg5UQSarsflhL4x7c1NjsPe
pSwPo58NJ0/4l01d5yCj8BFcAH3BqGi1HIIAV3fY+RKfLN3bVKt2LvlGDBNncJTt5p2KeFQHzcaO
t57krE01obozI48NhgyjBznBKHrZzt3n/TATpYRV1IIeDVeY4LJeiDDCuR4nnrtp0kyFFO6M6H8q
HJ+pa20yV5Zukf44Mp1VAP1baR1kviiqqf37tnnoaEnyecxluy9YgGcwjdiYQ2ARDQALcrjpppHP
dBCeX92rTo7kWNwg4elVZ6AV4gmqFIywoUuqEsL9VcEe26vm6YZn4PPaNwxN1pl/YuCoWeo8jMxf
9dWD9vq0GGSUhW/6Kmp92/1AlZriFccbiVScP+vdVaw0bsXk5yiZw1cWLO6ZTmhhE/OLySKe6so+
r0AgC47M9IdPJUNYhBBnRR2Cp4MGbJLboi0X13Qm9f0uS73y2i5NlQt6DLSf4PwDgmqWbqHfbTr8
5bJZnPRbLZ063rN8ra8Kg8q1VOV9TLM12QkSZbTQTZvw8JqWyV0rbsgLPxwVqsFHXKjY3TFZeSjd
7p7OuxdPzdJLcU23EqrmdM/EotghigOlEe7lvoHald1glR+iNeL+GjaQVyTFaGI5h5xsUmKKLxSH
Sf58VUfRThdYH89Z5HJ36ccIas0TkGYSEUY6Q25RE46q3/DhM/HJCKOKcVWzki9VJ9gt2ojipTDC
bx5Jy/Loz7BooUyb7QkOMOq0GZ90zQIvE39bMyb5sfhQGcjLa2YxGnyVtuiRS+hQE4pEC5s3dfsV
WqYH0RUrdSSpY46a1O61N1y5Bm+5JzBsM0VSbTP3QFj7KZS2Gb+eMNF8Mwmz/rY9+x1nwVdaLMKl
xX8ki7Wi/2VEwseC97RwpfVAUcUb736X5YNo1Gl1aq1q9Tn7v9MXgvelJzEDg2UsJilOCt055WO0
KxLw98WVC6OZ9k6Lctd4WdM7QN1OO8sMgeCRYqtzq+Fk+nkJdFJmtcEfXLFfES10WPWG1fr3HPni
SDgI/yh9bSiL3T5cIdvJ0aqQsf90FsDP6E89G4N90ZkpSwm1ehL5aztMMzusbyfUHGfBRTbQGkQw
6Wy0KjclHsezEcghA5eo8Ms0yV4eMI8ilBjognMHo4VsavsYgFkomzA90PRg/RvXxGgYdXWBMbNW
0aD5WqLUvsWTWROpJpybDc3mPpTXz3nbRPr9Wr9bypc6gyM/3EaH0Svfu0Xl05DTsbVck9yfdZx1
BLmjUv7HW4lC9Kebizrg01ZtCXlZKO+VKlkxaomY5ctNhxCE7SZ9kNNI9VvJBur2T5qR8+BynZh8
/OmEMTqcBH8V64GXAHMufwKT6BQX6hn2r2N49Oiw0YJte96Q6Eq5ZY/mzdZ8e3LzZeVlfziiWKXJ
Hdadg8bubI00k7ZyItrG4AACWjOMMSHSK1jnfxru/gPzjxopxP4iVI9olf/c725GfsGkfJjogrW9
BVgyiTto9ypHsfN2j/WC8CM3U+uFjQBIdq09PLOq60Mvq1UZfknimOtt/VR5L4T8sWsHOe7MK3aE
PfnrCzESun7medxkdkJ7kXsXRxmqpgiR3U6zus92pc1bs4FgBoL83ZWhRz8fIW6bUTuqBwiAUn9J
X1EBYRWRTk5fCjK+LbYw50DH5xGfWAfOVwIC4jRCIJHvxYOJ9uOVeUo58V5FUrvPNmI9tSurQoGy
fCv0eo2D5ov0VqoQsd3ZXRX/M8OwglPK1PPuQ3gbKjCyELlOyuaAfLoyEoSvt2fMBNjpv1OvOyLL
w+2KGeUWSBSF6aPb7j13t8TSlVng5tfPcLQZVI1KjqcrJALvp2yOfaQse2HignAZRURuYwUCIGO+
eH8rP7n4zWSuX0PsXPxWFbK7VRFIMqjjMiAAAF4CTWA4mFNgoo2QQ12mkafDs0qv6T+e0ZQ0PhAI
qb7JalYNfx8p0ATb8my/sPNmTXYnxohwV9Qy+ktsDKQgP9Zfh3wPjm8p3mNladXEzb3szwCGZuB0
prGK7WuIry37fWWhdTR0RdtFnoGbMwat0/nXpQVHS3uBYs1vMVN+kHXBu77TYIKCDH8jffiEw2F0
DImd1AHJN8z7zBNXkAwbu8oiEoIdpN4NDeY5+Gj9MDQSD6plN9j7A337nq9IZanKuX9qZeudBg2+
W6KZGO3prhusQa+FxEhK7CRjznH/yv+TkD87BjJDxuRMePXdyYmaVvXOILdtdCVEl+IjJn+EFm67
7gu0pfYCwQKqy0VQHa1nDQWBAbAgUvS0ulmrtAd46ZVJ91n+rUxGx4qdoR/LkeAi2yroJmWwWlrM
Yj2vXXXxdz8aURvGoyX9aOI+nVuh2FtokJPiWTI7WYQkRKin4SNNRDBAoximTvF2ljVRhAKKDTJt
4bjpcTPt+w1KYBddFqWEMLO4zGeAFXsRZ6RZh2K5wdOmYH28/GiFJ3A9PRmUatm0+wOrA+/OUBlG
5mZp1/SSMxyb3FxmfB/BiE41MBhNBNy37wBQZDjW3d2/2pKE3Vd2Gc7X7Gov8hpGTSCqa2DgqyTi
IQxVXdu17RwCfZiyo0rvxe0ptDmXE99MeT2p8aP6mkztBLQtMw26XE1FsRF0Ud+n9F1bKGnpv2dw
vbKtU5fe2BA3hOhJiiV6j8KFBaViFCJJkEBTWcC8x2Dl0MfNcy2Pyf9n/X2R2ab4t/mU0ShPz/5z
7RSGdNREYzlYJ7rKr8aDbcs9DAuXbtgkkDGlKw0HIIjIZLqqlm/o0spbn//3zr3YdepChpkUuWbd
eBZZf1+di5psW7ZubpFwG132sWLwDOISt+DOV8p3y2wHnCezqoQu3lJpCr1MVMoL6nCBydObuhq7
4PU7giUHXU1/Eji+Zv146yzLW2TA2QjAcxQSALZ1ywB9ThabWMEWee/JalHJFKaeQF1fmV5DJt1t
6CFIQ27qELRJK2+Lnqk32IFCrVxfT4+wZ7WnMSfeKJUEoEa1CWH7Ik2L92hqNRP8cbPFUk3WfCDe
bK14DzjnOg+0cAmp+sNL3RY1d0PP6OXQ0QHnADFnuaPhsPYsVAhMZ84Meg5VAWwFtyU3ayQDPljX
DsBwgnW8fE41yOz+Vrrti8rkdXWKn3A8H0Vsb/YeiHOGuksX4mNW1utMYI6uniIZUaTeML2geFd8
jiUktRId9J0qqGR05/rxX2XD/VkU1GdxOxwni/pNXpioDbBv8iGp0W/rHhRrcpD2q+/5yp9OxfJf
Kt2TpIx0kK5GydDmTni5bHqvGj54tfw7InvK4HEdWiHiaFZy+L+s1+ACI/0vGp9yuWFjlVhYPQ8e
DcYwOc39XxoRZmhS/dtAD7NQQ5JO7oRMBpKxG5MzUbTD+/knB/t7Y6SlqJXc4xhZ8YdeoGXUrmr3
9IV7/GPKGGfA/W4bWjcAeCkunHid5MKJ5hoHIKozsg7pJzSXCwygPe/9ZJpktPJwbxF6M8lYiARb
3h3IsO5YdwPaAIOlXQj1vTWRQwyhhruK8PzF+JMc+Q59syE4ku7OLdZZTGyE9W9Qb3nEwoak9jYB
aTSpMPhti4B+Mbjhg/ZDAbwy02dLc1C5N/WhaLrvxoOLqPDh8KaDPjq9UYe0ihefMARmvOU+cMJ5
ewuog0Mt60Xb/ag6LCmzQvCiXYY9I1DF++IE+w2dbftloVMq6c15j2Kyhy2HywhP0Ww6b4OHWzOb
V00G3jidTmwKMfmNKNmz81o8Wjvt1LaVu6+1EhSireOgwicXCz+TQFGAJNo+wKDqtF2SjYiYte8c
43KhAonXhTCoJUCo7sbCghGr2dLRcEi3GwJ67LAVdPYDMq6b0ZVsbPv6y7Ql0pIIlCrXHcV7OK86
mBRCEo4MopGeGLbmbhOlfggp9ofqztBYRG81Qjr4ge0dAbNZwIWHH+KteKpV7WQbua3LgysJ13A0
a5CRP9jJ0qf767zo2swjxhIZnVO5iriwBlJDXVKiU8jGfscB69tJ/lSfozrfGEPokOrYGRd8W0pc
PFpXOzvLj7db/M21z5GVxsOpfedFjGA5SDAw5Hcp/N+EIbbspuO9pEIlbVeG0/6Li3ZgG5XnCxLn
W4LRv3sksMn4nDt2GTRK3lVPBpFf4gOUeBIYjUNTMsRc7DPTFBxx0ub8LI4hS7yQWeVLNKvu2+Rw
4CZBtfUCRhXhtEIt8z6YoRnNTEcz3jA1OvHK7E7rKNwVwr3GuLLQJmb+ycLOMuwtvsVItG9ZpU2m
HT0TMbzjsgEE8DvkRo0yxO5NNCUeAP2r/fDFYOax6KMqkuAufssvaLFo2EfcQ7Qrn2skCCtQtVAa
2/vSyBNr0FJrwEida/kt9GeITov0GN/f02CRqgVSmai0U7euKt6pjRML/iEvQG8iJ85D3DrAQo5u
g2CA04wIsGw7Lm3wk30pkzC/nvPK05BP4R7+iBJV666eLc3hkfLsYR/MsMjyPFnedvPr9Se+bqEI
duocCZ0usvkXKsepDD5i7byGDJvyixslbVX7h3dJ/wdEhymacX3H2I4asJ2I/oNIhzXPNhWSsXxl
QS1FmvkAl38c7mn67syrmdcMkovqgXk3M8uvzL1pBuqvJZY1VnqOZH7pSu+Ok0ViPb1aZRV5vWWv
uJuVkcQURXKHsBmiYjYtN1F7DRIaozWdxi2lN16LIIbZHV0anPmFuQ1m4RYhvVjcFX9HKJM9VVli
P7ml+3eVTWx/wrjdSE9kPeJJ+UO3hxF5tREwouLvrRLBq9cTGTYHXawdL3FPdHVEQdGXgLqzaAQY
1tAemKpP9YHjwbds5if9n/cqnqnEn4LoYF8ZQG0IDHB5AjsYgDhgCtu13f2LvgELClvTa6YhaBrR
Ko/NlYgcCFIyVJRqTbwXDi1JuGgHpMlrRe00VccGwFbhEwfFToxwodAjzLhvnU14xy6r4fCKiz1M
S4f26nEy/NwX5radXY+1ziZacZxAOwaMzvrIKTM7WINWRZ6BRXd+S9nD6GdkGElCJQbGWAneA0YM
rJlE787xjY1sf61l12FEphrBi7RSom0DiORT37CIRbfJYYCmxFRqiV2E0bU6FOF5ZCEUTXzJmTXz
7FXSFHaMeSrUKtOqqvzZB659VpS6RyAz+pi/1FD9qP8mEw7N6R+M5fCUQxJCd0AxTuuEwEHI1bh2
cThIjMMlBP0DiLlKUcPTm84rd+HSdLq8G/cEsTrZEP7e67fEAx1f6y9ro2X+DO2unEwPav7vswie
xPzbr11X3ZZby3QHRX+7hUtl5dY/3jW4WR7CiUy4xNK2VWbjW2SFOLFdbUO3i4LDzdqSile4D4df
jloobvSk7a1QzKmx0UOy3Eisb35gduXXrg3iqXs8ArVzI2DLa7Pd4k4nyypIvf5sz7HU5X7kc+ms
4nUkPIcULUN36hSG9xvIg2EahFWHRMJHOjPTNiFKaGhtrsNcdPzGNeRYBsgyRwbJ8RfReFO8zr00
OeNQGbUK28DqG2igMCqTDInYBczE1fCVGr2msFlM42ySk20/CwIMlrEClVN1E3LTD/v+x1l4hbj7
VdvBOB2GI7FdsU+/J+2QGcpEbNNoXGJTgpYzcvbKjo4ApvHn3TxI1KCP+nUPfh4RMDupX4zZyzM0
4/ZpVcEwf44xMzl0LxcARMueYdFc20B6Mp1YD7dAH3rftuSbhqlFqk5iRxxaCQRBZkhydsSdhsUh
rXeUdYsgrsqG4b1dLGybU3eZYuvDR8lJdhwBrVoHv8Fammi0JnCosu/6IvfCvhEowQmcLgC8oe7D
ML20ZHR48blnjihg4HRDhPHo6iS/1oyHwuY31hp6vH1WMumyV1arUJCI5JDYtSdw3k7YHGQPi1QP
AsVOBhHFwuk4iWxTuRDgn9bS/JxTSqbI26f0IawSUe90ENgYsgLsZLhzq7nEdiZMs9XLdbS3mmqr
Q2yX5tYh0zHWZVqIHeFFlnk1XHq86PKXa5nHjWkVchrmg2Vkk7AQpjyX6Mn5FXYrSSzm9kf31EfA
CxWOvD7lDooh3TVh8GWN3OgkMwn+yWUbvllcM8ZcLmOJZ9ujoEO0CqMErkdbfsAHuC8Frh+D/TgG
WIsFC8Evr6C0Mm4rOsTyOgNTIoytg7SVMtmoAxTObUDHpsn51WmXsQwy54oJfIQ6WKadtKoackr8
M56MfpeulzQIwFdNaXWypCAhFbpLhQW2J8DGRjgDE/6AcqtA83DFypMU4RSIXxAcAfWvb+DPLvpC
0WCSROCzODATxgv2t25aKzVB+0EbhXX7kZlP6XQsxF9I61Nwm0A/zti0BGG+tTsZ4JUqSIP2BNWi
ywreAhPckLKKqJUmSdR7/7G25/cqJ6EMA2bhhuFazZH43kiPAw1BdklDL3WycKWY0VB24tv3RZKT
MTNrHcpd1pCxmvTUHhLsooajlT2EhClx8bRBsFAWxCNO9GxsgTsnrvThcjnI1/20TV3+loJADfFn
9XkB7BglWoh6EYbm3Fi93dapygjPAm1Oj0J845EvzkI/mNTIHH4BrolzrXgB5ZVGUvlwbxRnzfQf
i4KwdEQJ4Og1DMVOwX37XZBd2smAHCZwVae+r3kqH9usq+mHrJ29PhW7pboEzVpwXUt/+EoSjfS9
ES4IoRFPp9UCZFj+vAHYXO4edN8KHbcbkUwxp+Lbj7U2ZRv1SNc9HBjvMNal1gmJLqAVs4+jWImT
PDRRLoTnF6AyoHb8NwoPOuMf8LUi/TuaUGBNbT0OKZRexAkIGLt66dnG29I6lixV6yirPILp5450
QA7duzSXP2+XFNRYljaqctx3uR4Ol9KxhrGutWehe+0MgWKiUtV4yjF48AgH3xc4IQsReLXdo6wb
+KMG64vUdLOCG0wQnzYccr6WG5XpL8Fkyc62T48CX03P6XRDr4sDrrHaDpnwckR6c2/sNZOmVR/o
2NCUTovcP3KBuA8o1lNwstw+77bnldWvSLY/nj8stS4zHI3hkgNUluVXxsHOHS3Xxf9MAJdGG5pc
1CK1UpHyXlGoPVKaaU+5xGiBwaVBIohBszHf8gqTe2ry7cIVx4pqX6PbEr0f19TktD7WBnjCre0j
IE9PH++3Qh7FdRduwiXjwFvp53n3TclSYXDWHTzNlqCDwqvXVAdqGg9pBlaTLD6VjzCue80a4JEk
r2dHo+10S7EJ6k9Mpx6LBGkZ/VfoxgG7ZC09pons+xW5NOAG0c995aK+76+4IqRxSo/k+0C1Jklw
uuPY31n9Uo8wwAQPrgasXKryXNziPS8cpXtHYw/ZyZOlF/+27a9gcaBHG21eTTPUpJKSGzNuOlXw
nXB0qi6BvWv2bP6s727O/u641KKcseI+m7g3j1oZnKjLAhRVkO0OovzDRBXHwl+xM/pV+xs3AJmj
h8DTsSYk1xdXcaEDDb5ik8zY0xjF7R6j0urGsAxabJM6suMWJlUvgB6tiaFXU8iEl9j4Iq45GpRD
WKB56KpkYPX036SECjyEgLdbLCSZ0j6At+o1gjg9QkxTXavb0ALLKOKZ97vS/MbDXKTaq2pSg2JM
E2j0mBD/VE1pQneg9Qrk12P+XKk1KT5slxDpoqghC9mheXP+KBRCIRAh5zkkp5darMyUt/byielP
4GWfMhPGMhKWShMi797njR6aBari+/eLzxkVMBoGRlqCfqd6F819mb+6pck16P1JtMF4AdJLsrAH
U6Q56Q4II7JsS58N8vhV1JnROiWSvmnpLumXMBWlBlatLG5V2XwfsRWn/hiefgJy3lxlzpGBT9RN
kV+UdOYR5PQ90fsGuPu16GjX59YjN0se3UyTUZjdR2B2TwXIgmqy0W4tp8LhOMMF76HYYr6pOSxK
Z/yr+OPuVwwvnjpzJqMrBprHrJgVqlFT8dqGKaN5oWMXLqwunz6THHOMMM43/kpvhUdBbfvtaN+m
aohV3xCh2p8nrTI/WN1uzvJSsKVRJSYnUPOxwL6RsDRot3X8Hvv+nBjgWKKa2ZaYU2oww3BKd01g
uqsXvhEtGYuyuotBA1y4z7ex1UaD3j96pO70ObKW1rLQWd+ezxW3MzYEGT1wS13WmwglFPg95sWL
M1W0uLoEn9vQ/v96AuKTEE5nb3D8QfliU8WRKY85bRwXWUtJNuX1lbjD3rzXtlN0i0PrpHiSQ3q1
8UEzrihdHIJ6q/04vjqlu09mNq9o7ZCp4aTi1YiMExQZr7ltEfMa0NSyLYOEQYZitXBVaqiJicfA
xkOBxMwreUsCGsj8sbcg59O53/DuL0RzP+HANqTJ7tnM3kCGWApkydiviQQAuO77UBC1isd3lFgj
HdPfUkzA6gjq17hNY9QrMQspdAU8SoXvhTBVY51FideifDFlj+vaxHxcc7ZhT0xgs+Pktg+Cc0ah
oxnaN6uEZJjA04cJamfYE6RfCcuIUSanK9zbixKTBraQSQ+SuS46+GWC1ROGa4TFg0XyuSr6JtOR
caGRA/JtKP2n7rnRNWyxpTLcYVKtAtbA/NHnmwZKuBY3aBrEBv1x0qU+ENIpLqacOywYDSTOSAG5
TM282Ac184Iw3FkbHS4oDgCYN1P1B0XHgOKdeNWDSEnnJitJkicYzS1PJxOasYNBuYFt+gZ2nkyD
Xpyc/vaTLcZmQbrr0tC+aXDzJYDtAcdtG0kiNs+iSgokHPPgF8NtGn2kYgipwMbJbotyqgn730kL
Zv6nBJNPM95Iso+4roKoT5etYOC7RV31JxWDWTF/jwZ+fqFfjnmgc6D7jNXMPYsS0fyjDvELPaHW
HMxfScpskUAsoeHUsRrlR9Wy/OuQC4R9nN1mS3XjsXcbqTcFk/7A3VNQun6DolE6cwFWpf3YdgdA
h9cYpEMRLv4jhp5+4eD3dAeyt7HrNnVnL7w8n+Txn5U1/l9npJGWntaO7qGTwWTNb0797nee4SgR
hpC6jm35xY7lnzfMnuiulnY+yC0cMOrFcxFB9KniW3JoAjZ+dGpGZlqEUBu3EQHngFiQzA4o5/1k
jYq+pMh8hD5UIj1Jn62VPQY+mPRwATyjXJ8POiSBmXv0A7ooU8IYPPMOjK5cFP7RAWPV9vky/vPp
AkdszCdWf56Z8xOZBZVGWM8SkTgV6G7WPwz1ANlTv8WwClQX3Ew/2pSWfcQuNjhx1B7doY41bDU1
/cPm+EYQawRujOT3GxG9WADyfrO3v60Elp6CxR1Rn6q5GfkIuPmrfbKrBt/FyO9TtZ6dnnCBuQwB
ntLKDFjaKGpNfF+T8FPzipVqwo89ok1wegEniWDZz9NK7/xFforObiebGHgRiIwo/3eXUnukW6zf
i/Qqyzpk5yBnlScWymvhe5lCXpXRXAfBxXnnpk9QbhOfXUFAySJ+1TwZgC9BvJsCpyWQfxUJ6gfK
Dm//qIKHqJwxlSQdqdGefOr1QeM7U7Qxr+KIImyHhBT7AJs8GPNTwVghCZ3n3Gu/CXokPjd0kJks
kd0LMrPV4hQPy7eGUtN6h1Z6Chn3bEiFWxA9isK73Y5SdtJIor00oeIQ2fSuEpWT7T5KGt5K9p6g
h4ISb+DvQzito9x6PB8OEqWETKCBHWSVo0FuEQIH1ZGlz2Lh2wyAmAk22B+yqX7pjfu5OWVZH1QZ
5rPF3T8aEqjV7DmNERz4cS1Z5E9qlYRxKugVNLPhcsRWYJ7KhZg1ApYFcqQRPXIDiB3hqEfI0b3c
EmdTwNaLhWsSGwR5wedF8GFKBFlH/gpdF1MELgx9RZ+9ooOzqr9X5BiCquQkYvVDlbNiqGKgnaGZ
W5NO9PHSVI+C6mB2EIlY+elUbLsLv1cqyIcuSLy6PXQKq7GVB50WnuLVw9YEqLs0K7thjBrB6uzi
iDJYCwlADyadcjN8n9eY8Cf9Mmenw7L8sM2R6oYG9S8ojskGP6lO0q7BQQXJWbcwB0r0A3xTVQ3e
OgZtbj84EghSILynCLjo6DdzSoav5PD9G4pgCa7R51JIGucRBbGcwX1lo5YI8LW9gMiEY+OOpV/G
aWK8V416d8ZqsK9Zioy045hdv8G01U4FstSYRSPVN6YeQGYEy9PQM0vK3q5nOlPNlguh1qpvPyby
y6Htd8/z83EMKNdjEk8oERqLg9dBqqCUDA7sFDZ3qW10bRA9M9WMg6C6G+Wt7iNobzfSkNAtE2YI
KMzKvzdz4Dc+xc2z6R5/Y2Z4JYID05b8qnihXsZTwdwiGwrqo7Q1aYRW8RgkWQwa9z+ZEeX6i++v
qXKk3wYttILfyMN0l/pbDd55rQV6ASa6mEvj45SZ5FEq3JuT5hiN0g8Q7hidpuzgQMxvV08NuJRD
j03lZiynbqqVUXEVeMOASUVKcKuZO2OIcrHG/OD/8h7K68exXtJtU8klpW5yujaR+dVzO7lIZzaT
dX+CtS2ZJIMcT8c/usV+A9wmYpOJo6E9WN/zfl5fcFl1HPweF0YwM+qQMPI36EvX4gRyalDhmx/a
1Hnlh/DOSnxqBcJ1hAkMIxsU0jXn/6L1FsQaZ9v3YoIwe9PU1nugmFsAoOe8PIQJjQWR8m9VM+JZ
KiKzaTpoUNk3ekQOByB256GcQCos37HLYYJR8/d7pe8m/jpomb2nommQ+CdLnjx2LQaFmV/JJFws
kJ3BtSVd5Z1CADCa7ePsVECMdtT69VDuyvZp5WURh79k0fj4VdrrDkMHndw152UvssHzBdvVXqLi
rubkHlh+6Zk0mfcQq5FntP4WGiVyR8hz6vDcW65wPTFf2ywnSDyH7c2qiX9bgyCCzEquk3NtUP4k
G4+3iw1G0Nv4nlUAlaQ6sQ9AflxKTYcyL27sgcm4JdX4h85uO+349zQE4eofJlwHwTl2UBp9FeeP
EXTWeVOgAHV+gs1ZOXodqFl2b5T8x+svI+q7B0l6i3z4st2NCI3Sw5RLIFQzgtLe/PcxLavvoY/i
vOwTWTc+uXDuwCRgBnRAU11aZTBDjLe6YkyBLf5dzgFpEY/t7QtAYHe5cXo6MWzLBix/j4X9uPDO
20kBpY+cD2JklRT9sgIV7LU+KIvPpkJyk/MXKPoCiw/YiteVIpYWXbNroGSYJsSHBd3UO56rvGMh
JTyFLlimmzdkQWiMYt9eNlolQuQBoRGx+UIMAo5qqds6yn3iuODNNBkBogW1C+toLTXkUDzY0XzZ
fIHxgsEHWR9mPLsULGwEtncLARk5ZFXWEy6RLiVIdsA4EZ6UNCufVnMU90yX1GiF+rjG3HOtOmOL
gQ0qVCHBQjjlt9Vm3VCHdSssoRQai0IjawJ1NVjL3hg8c2sWxYFPhgalkn+yIVKiFbXT0c2T/Vbl
McxOPD9l4P+AhrUQzBffjBfZ6M6meuq2LfXu66qhBcrNCVpK4LcvdenjWXbvk3RldQjMiLSRINWd
ghGf3tyGfjoAnEgRNZq63/p3fqB4994f7VTqcerwZEsEkFzK3KolSTqui5ncwzRZKs4YQV01glXj
/VZGFGL2bpRgueHxFYXVZqmGatlN8FAGr0gaChHOIaqQcjdP2/Wv4D4AGSSvdptyho2GtjCskQDr
aR4whM50qU4jCDuxxQwOYcb+7DM9UDaukZDwSYmy0WsXOIPCUfWQPZP8JTDcC+0+DiE6NHXiK7WW
YcZ0CvSmW0cTOnNxFs1rDelw3Jk8KjQAsAq49KVNk0K7kWnTgwBIyXkR2U1EeZL3al1OgNhsmqQa
rM29R9OawxXnGa1Fhlw53cieHH4SycnIHRKTO+7xiK5Khm6bLn8XHaHywg5wNjnxWXSevU2L1pay
RGFnRNeTHWTAq/huU077lroorwm5hg1dlSFM841sEbW+UKEEkd+OWrlVDMagDvOq89NjCDuxXDPD
nTkBoTEAe5ROzCfJC5itWa8iKtkG/Ou+VBxw/pltwKkE0AezdnTcz2H+Cr/BvtVe6Z4AHNHIJsCu
eSdCVaxLoG2SaOE6BSPznLHirGuDAqipUCx2pDFVNaqiSyLjYZpAJT5W2h4i0nu+ORpDB3GkbfRa
X5L1X8tkNzooqe1bSNAEclpsdwsLQVk8ZZ//7VWB7K7kjArmENGcITkNElPFCeq9LxcnBuROYZKO
zB9UVBDXjDS3QEpdohqAGu2TCSqEWqvIY687XQZ5T5EplPaTR1mRygNB86QYH/BO+8MpD5FlrCK9
1ALXw4b9Ja4znlQvJ7Pzu+Alzyq2smbu2M6/nLdaJ3GRcNFHdiYD0toCBhRzvXI0Rl1/mTdYiqFz
9WwJ1ACn/cm9NyJ0L64zaGvxPIMf8f4dn+UWBzv820uTEoBoEwHkKfbtc02VKjfbHlY+KX8bEgHn
h34a8iLEj3vpt5IJYLtUs4FrpcnBd3hv/MwJW60vPTqOVacztH8493ENmxvdOjE/lSW4eInEQJIo
Zg5HOj1Ehjvi/VU9l5SjWB+EQ8JdklJtYKCBLA6pKsDVUYzFS2TLWJM0J/YDAqWRaAh+q2uh0rAk
qbUPLUd5n4h/+EGExX7G+RyIxTXT7ugL9m7q3poved4wGKa2e+p+BNtfopkp6PCHriH49SAWLwce
4Bsu6xlRtBawzCWEm22AReZuaj/dPNSEhYv6jgxuUY9QWTy3syRXcaOes6rpgHWZftPbHsrRjpRp
TDHkF5FcPy7Nvrc7cH8tveugnB4QDU+LSTzMbzyWTAEzbFD/rp+e1M4Naji1nU3ncPNKJAekxMtK
Lv2eTeRhnsGYTLDvOeZ2ux9ig7eyOsAFEPJITK/3FriLks/ra/QeNkGSqmmFtQTbp/6eOxpBJEGI
+v7xX3ExKyts1QrK471jFsI4K2j831RNpRqjAuRtFiD0KJYIHVqqL/PuM6TqraGwLcenrRVumUkS
lJb2fFTo/GAUsO1Qi2gUoS5JDO4pvp8psokqo46Zcvbg9pEIpnrSEgPm2XheyZF/fzAOWhRTcvEh
zAVkVv1bDcu2ZsgR+mRtytiefeknGT4jk2xJhTIpYUxcLG/R8CspcyIHjqS+kecq0CSwz3F3PF4D
LgchYj3sD33oX3fTCFG4LS8L2XOUJg4KyDZDw0Yb3HOSwK/lCSQcvM6VONXz6NdqBHfe3voDPWlw
UosKRMeHiWWTLSbPH/5iyG9GeoD6eR3LfoG49lD6GceVgfISoKnyWOB2UHfznsDlkoRcT5BlPdjk
6Z/lPKMw8OW1DV2mWXyAQRfY7/9ltEHK5aw1BRVsDqXzUWZI0jEL2XlAPg+3TRjwQK3K5YRY/x1c
IsT2A1WWsJMmOgfNqAfEkFZDFIteRYcJp3UqbjhpJ5otRxQaJEym9ZVjypx7aMZheHit19aWbB1E
+HmjE3HbYiCAPPD5+btAP/zYPZJqRvfpuet+imkC/GCnhP2l40eR3cI7MSxyF/LktHMd4UP3zBil
HOSL0R2iuftt0J+WPQhfERdqOMMDNtTeaf4gyD6ymnCrwXEaNRl0ABPNlaKwOm0hoVBdI3yvjbzB
+khhWVJKxQjY2x2jibxc3TKhnVVrjB6ysRid3RHC91n1pqgu2GFeATVbtydKzrZ/cZtlhCNsQOWm
6Yt83lzytNVTO3YgBZJDikMPJdL6ozDvvXOYkkt4w7vWozFl8x6yhmjwfV/s2kHfwq99BRbyRgnD
npbZf0ZV7nCe+8DiYYNvEGO1e+y2CKmg6nV+Fi5dNHgyjOxYa+nQWjruXlthfEbF5PWuhPzr4BWN
xysYSscOVh117q9kRWzCquPeYX8QRHYl/fvchY7ljQtJ5JuS3rlhoPCkNLN+9/rdruHclngUjj7Z
IuqsWmDEHaiYaUiwC2Szk4hHDGRgWiCBztz0W5UlEBsaeZrN1mhV6XkHx/LuLSRDY+q+Guyn4sQG
t4bUFSKvBq5+I60cNOy5YGKh6/aVRLyCLlcS8CXY4igCRhye0uY2itmDKfRrN1hvknwIXo0ab9YO
irOvce4GHkaL46Bxp6nYzsv0LGU9LtMkdZdk/5D7ujw3eBtDaft0wQn63tdDAH88Lg3icb+zmcYR
KgtGofDPPszCH0dcUlbadkKagvfAx9dOhfEUrFmyOvpyOPA/MoaCHMpBKNElMwmm8lz1y7HXTCO8
VoI9vosS1b0+hQXYP1HDxTfgp8W1Gf7kEW0Ug5QHg19pEPyoYfL6hbaDA7mnrSrDisYffPOqrX64
rKPc8PpLUsWZC5AZzeTe/QH8kP0787sJIDKpBLRq29hXIC5cAHOxZZ3ok5EuhIGG1irRWCWcPl3A
zEEPRUhRQFb05SDc89klKw6YnI5ujYekIZcsipCTXta6/Sn9MmsjLh9w2CPEVLwlOCC49XcmZjVs
jogJ4mHFw6qsBMuwDsCrbrL4eYAWjVDYzRhaGz7wC01vQlMy1+nGc3CXNhYjExUixjJYLiFy4atu
Rd2iZhr9Pvil0BcPdDcGLm/gNXY8vTNDFYlt1CwoGGtMYmVLBTHXSMbFMUi4zCyp9udCEHwfFD8f
IYR2erQdMpws84jKVXeG00aCUbDp1wN/FQmrkpxGLcQWunoJX3jv1BuS2mV67K134HN8ufvs6ARa
yMHLOmlzKEsWiL1L+F3JXHFwBPxDZlDfpDt4WS4KEPqo61/Om7QiYUnicZF+5hhr9ULxoaV4zvxV
aJkKtfv5ILLQb9UitMxLUWd3oFQGEMj+GiyelyBzO72FqVNHod8I4vRqxprTI3YPmcVBEppoO5bg
OKCRwDj+LS6Zg0yxl5b06oF0TyQCogaPgsXo+Qh5IWShWV1MWZyuZajgLhDuU6D3Of67Iu0jvYta
NaTzw6EyFkZiCNHHbezbGjO8mdkiDVoZIPD9x4OqlkLfRlUB4MiyEt5R5QvkRrvu3RqhYdNI/u3M
VGdnh1FAH2MP6hakkpdc2jqgT1wmA46kYMy3JR5Oj40jXHDLuRRrZ7/kA1s3qsGysZoU7ULC519g
ykyTZrOG/DtFzPhd/O9whB+qgHMBnz6ovvabsm4pQOhBGUw9g1U+NUaQ8D23ptTiTakLZkK7Kctg
oqmbnvKOFJY6GFVuUM6oF/gzAqfqwIvUZdkCZpjYrFKaSgcnROzAexk/Gd7a9JsZ+4h1kCzeiUT7
L3+ojHYgXMY0cVQ2OxkkiDcjFU7J6VhsklQL6lf7E1YUpEX6wkcpFVSUe4a0uFk9/FdEFIalP9hX
Rrv/LFLXruyaXW7UDnQX1ZAUgO+mteISdGfZpFW0y3OUWahinINDYEG2p7/MeIeVoTqYA6BVlUSV
cvXnUamg3tB/vb+dAWoGOrn9Tf/TDnDZ8sKL7aQCqNaiT5zt9LJwHsFqyDkHl/MsVo6MUW1Rsg+L
Tz/1MiBdmKZyAp+AyvQmOClZvVQUUA5hKFnsIfe/gEGF355RcBGgL8Z2BPi2u+mc5WqlJFqc0arB
UuNNnMurmBSHOuJ6T9jjVav90/Lph83zjnTow7Yy5XQk64GVgKophO7OjwpDto7qEAG9oTCavl83
hEZeMbD/D6Vstj8YjQk1QAyplMS3xusmWnZDAiHOXs9QY41nYF+NVQjxpmxUH8G4RO8lAPn8AyZ1
QmVzxJIjOtky9uXjuYvUfH1Jd3Yd+0V7RoHGbBOmhtpXvCeHPCrarmfMsyJPp4JJ+wCJqQ3y7JAn
825vlvum12j2CRkBKBfao6chWdetiMVYRyDKWP1MfzqxcOkAck7et/eFA43TsHXEa281b6lQARlP
tAx6z8z221oxsvaCePTyDIhUjKPCUEavMo4B3f/efBkkEK6kp3T49AsBv+LT29iqYJs/OV2QeUPC
gu1HgZfK/9Hq+TszEcrwHaw6JtKd7VBwJW3RjM5+E7jW3zIEdhzzFu//MGvRwV4t5uonkhQoHydg
4tNfSUMUns4yWGLInh0UF/x02mcrURUstq0q1C5r+2EuEBpjtUdN6ASfnp4dblXymqQ8DXGt4d5i
7v4OXQ68NUYzv+TkzQCStmjtYFFo1N2iYlnqtX5rQlGE31Sno4tmFeAj6UGijNDl45DEiXM6+7Rz
APwAYwXEK8mVLRdIWXZSZHrAgxc2DFxEhS/cfHHYjljUn8RcZ1/c2e1Fy7iZmB3huZ37KkQzV8tD
hYM1483Iv1gXYYS1RKQXIgaFEHSaYG+hmsgGU4dMFjU/dtFHa8Es32LvsSqAA0N/bYLYZhYwOw5C
H+X8k6Z3f99SRY9gpKqXbbimda/K8OID3HIclXe6oCqyGuemxo9heflSB9Mmc5Ake3Hf/ioBHSKO
MlQ568LCLR7hC/uWA3Byvp89OpycyQFFWGPIHH/Ap/Barp7neUb/qn7+OeLoa9idGd88wpWn3mux
5Sd3O9kfIOKVIL4sIsRXbams+V+D1s6ziaw+4DVW91aJzvs38FlcioRnBvrz9S42r/sR8j2M+3TF
jff+nFnbCrvXWJpRQfOpz44kZnt52XaAviQu+u5kBNXpU04lmvmQXKMmtdrHXk2bTXSj2YkEwefK
Up5IurTu0XvProdFeXi5teo+buGr5NNL36WGVUSabHX8Zp1KYpl/XJ6z2HzxnES92YljRq+U/y62
FDW/Y0mPcKg+9xcZQ1KvYSDMG+Va3Gj8f0Trw+2ZhHrZCD3cdbWMAANfql66prFwwESU7i9f8qXN
S3cmLpVwx5fHuHyMlUgo+m8uWJOJXklYiPPmijK3c3ED/OiaossgxnD9V6G0Kz005/iqp/Hv5fAo
jndaL6tIK1SQNfCryQS1ul86HdgVAOTb4B3YdvSwT7DmVIvJoEGkxsQ3HSEZHUxzLBW2/PLMHFm7
jRg1BP4ZDVUvMyUUWLyZP7t8mwQRnv/m18azDuHMuIXsszMhpsODAzf6IFgHG4qQXkLtFhR1MtuL
kqnWbKM6vEjRzmdu+Bt6RHOrL1/LuKZT55qVvL4Q/gWBXvWpwQcj/vYp0OZq7C6l7Jo/s0i/unMB
MMMdTWEg/CrWdgn1gS1w7A8KR0X8TTlC2OyV39xWiy/B3OS+c4lY8M/T2pqVfsYvxkOYzNKM4WVL
gCRMcYzi0r4AcnhvOkonQZX9KECxc/2he39B7KaCjlNaDf3NQS3a95ryHBY4fEtU6zXP2h+pZvuN
a874+LYRCvKSSOTiNCVd20EEuewdTgID5zINqbjtnv5acGeEjIXyveeUJdAPOfvbvfKGB2R6c3gI
Bj0r5WdwL3rHMFMRxHVGQueWptEn/aJmnteEHMjUJXnoHtVgUNKR75Iq/MsqCuM0iGZOPG4I4QJP
Bue8ZIIG7hcUSsk9wAbDB4WgZT4Ym6xbmApJmaBGKDRp9e9DJ/+JioO4HJGCMbNq2e+yJg9/K0fJ
Lh65TJqsncmdhFRhgKiRXJaRCvg/n4S6sf6pKvrFqBqg5F52FoycZ8IPwyIvYKESIM/FZoEarsu6
9iZlf7Zf4YvBpKGNm82SBJ1nRsVrK1+AGu1RmhhIx4wYpjSWzihOLkCeMZBZBDUo/wXajODvAV+6
buUmpBGNWVEReVc+elztfb95kr00XPGyCTzaXhVEyx926H94dQgx2zSkw0M70r6Lt/YfdsIgmAU6
tnWftjymwGAztH6EsSlnGhVxKz0J+2oKhLUvuC2Wsg8PkUaubs9vfp42nf48Y4t5TaXdi1tuFVEa
RFp+29hGLrNPP5xfwSeWBQTSQlHL8FcMDpEMPItm+8KB2ZwwgFwT9oM4JAs0QBT+CE0INm6r8EUU
vAWIc8shj+DW0MYi0B3o42Gl0CLX+W8VBRA0MOkkbRDBvARc4vNQOsO9Rlh0xwM7f4+7eqLWbNjs
1yWvVf8V3alwFiHO4tnz0vpPs6rMYXenaU1i4FTycF6bKY96Z2z23T3h0NC+kbFEKofwTdnyiyTi
+SreGX4OsJPC+77lkRdx4KJJUjhHu763qt30q8nNgtDo8YtiIkJtErtM6fiKosSUoOqnwElRwuO0
e88w2NDzELAjOPa6VWIuVB75F2hhXRZyrKu41M/2opuMXh/yrQIcHM+iCm5XX7QwVshhGTdZM6HL
KFMb1ZuVlsVOygpI+iXucaWXQ+FdyQ1sp6///cvCaSQ/1hUnJLUMDK3054no9JWHuQmW/40Z57H5
NQ/WGx9af4/daeECh9/Y8+KxxpBS9x0M1onn4hmeNMPgtAfHFsxO+m5jcpBtYgbhFDF1/dNb4l56
FOn9YG2FFjv90YIg7Np21X91cQN1yfTXOSvIOn7H2uZfAecCrzwNt6dxD4jF7AIahE75p6XzQb1g
tTzLpSL0cwQwZkRD5z1ReH/RqxKdaaKSRhMqjhpd5N0ozBFHZC0GTuan5a+K77vk9dDvK2ckwMwD
GPj0X0damOspKnqSPOPzeQqm3FFzPpubCAJEVB5v1yMu6UU14m8dSIve6Vl2Ci/wnmN0oBM99giU
6//LFK2pGbpSKJ6XNkMv1QKoBIue+DxO0Dmf0AxdKTFFm2KC7us8U5WlkLJIfHuu2skDLJTYIrkN
qFZcE36cyKlsWPG8hV+i9dX3fl/f82HLV+2Gx9xRGS5Klhrjui8hLL7R4pmthHmID0LRASS7LZk+
3v4aUMAxQtBKt9FwrmLgPrL/1mKZRen3TT5t3fjOYpnAGUBMNLWDjUxSaqKPIa5qiRlyRywKAU9v
fhqwCN7sC6XsJn/ZLD8fAM96ToKji5AOkan3vB16ZXb9N/URj322NJ4tQlkWqnAN8rSTIVjwys6e
rftXbqSLb3Vm46f9e2guz26QoOE1wMcL8uTprYmVUMKA08BvinSgDlkR+1a9pTRCdnv9TiJB0tcw
a5UbKEL7sbJTD1ouYX8ioeSXyIqfEoSAyykKLjQvz0hM64zEJYqYaodHzLNzIRGyJ0gi73DMCPtY
9OE8jw6FEwVr+cQq7AZhqYx9LnzfZ+JbDhC/4H4NCyOzQh8/0JyeQMM4rmxyZSkLQ/QyAsRkvywa
mgdKDzTtuTLhqxpE7nj0ADxfM3qiD/EHEJPa4tKZDEwiawwm1RIsSPz1wWcD/CVGjaQc61sZZmCM
KinlZ8eDErANb2fmdS1yBIByxYV2i+yYUlE3ff73io/PB0fgbajrRxlPYsjWFrCXwqWmJ54TUNF5
tB9tbkgFsDvuLzQMqaLJC7bIHXqNfMfrJjrc+6woFWgwSfcXjjB9c75nYRuhAtq7M97kuf9fPR4r
vU4K9utGWKcl4Wo2rSRjMG4mlndViFN48HNTjqAzWHt95hl0M5Yg1uXfXNDDc1LWaTJdoC5T/F7G
HHp7GEK47zcVpEeNTBjYX1RYwl5CEIt1oVIE4FAxNWyyDO8hAG2hulrmBUsTT//rXD53oVv3xbVo
kEs1Q1Uqp3Xc9KnrX6Qb/O1181jZHyCypRDEFr+38K710vqRZt8vEdHvHF7IcM8TANAn0QsHcLr+
l+fgc2LGoztOvscZyGIBna8ZsZdt15S4p1kl5m8snRsOm/7ZSqgsdecW2ukixzvgm0Z4U/4bpKKs
wiBgTT19n5m0XLnRhZPFowIenDgeNGoQP961iqINi5qAZXBdfhu/BeIMnW9lKsc7/fDgNOwzg4yG
lXhp+1Bqollo9raHvp3FKb+SD4KEIuFNY4tcTDDBOchiwjE/r+AxI5T/6j8HbNnxno57sS0LZK+U
eTWNkhjKqN7Vnun4csPEYQFunfLxtytI7gEflnlXqHRzNBfVxhqxj3p0LlCHZFtUSOCxgYWiw7FF
UgqdUGtXUDC/XsK9Zd0ySjpvFOzPfbtrfQMR5YulMDCiSCshXOv4Z5rBWfOZNbrBbDACNZlmljl5
/QvON/RTUuBf1jIcbmm20a9eUv3IXtPcEvda4heFeWxX9z2RLbkcrUceGmX968CUwC3KCCC9cWkc
gnEjdbQg4ynkUP18oCKIGDdm8jqdLPaJEBPhlmohlTQZZaZCudtdT1YH3o+5xERcPiN5kaCzxbME
dttQ2wS1drdC+sAylULdDfCiLHORmebbay625Al16VtfWu2S+y5/LE46H/0EKP8yECwMJSJ8auVj
P5TLa5PpdY6ewNWKrevuF5yFB06lHuBLLnMSPhelbkbjsAJyX5R07pX7Jd8NriWqNG1wPDOV1F4s
lJJOlcndi4RDUbIzxzU4hUCPRvs8OG5jwV/0sHx/pPwfuqo6BW2LGGsdDUfnVxevje+AhKDhby0I
gXPW7ptt1TbwgvAo/wUg+2laEBYFOgZ0EP5m4Z5c1V0fioK+Pcww2ZzoZEMGcOyU4PW/FoQYhGtd
ykC/f5PY+Uy7cyMY+FzC9h0lskCYStjOfQsiDWsjJ5Ibw0+BIX2ISo37OI4zCKnq2XwbJRB85FPb
gnOatMj22VBpTM53v3GaP1XobqpkRASkmPFCam+dZ5j8WJsj5P0EIa61dfN3HkD8cRuXYm478al2
uS+XmkeVodowt3rkgyzXgPwd8a6fkh1c2xzN+cLrchhCGTASUkf+Xagx+/6ugx1HJeemh++elZKZ
8OrjjjExH+uWJDOtPxf6caEni4twAAmWHtdGkUxkU7gKhdNtodneGnARPDV9C3dPm8pjtzZ7k3Op
aYlH10u/FH+4DLQUOUBkY/L4AHBv/+D38N9bQLhSAMHQGKMzcYPPxksV5iSsngFLZ4PXhfhnWThR
RffaJN8vHb7/xCoSC4Pj2p50kBIsuj1CLqiuSS2t9YLz/d00LWi/62e6BOAzvrz5bEuZZWmv2zJ5
iIBGChoQS0J+TnWCi5G8JSpO8lQVns0oSTykbRXMZjxF4YADF4ACNi9UZXx1GRTysVeBklhhFzU+
F6mkZANzQCzCfwRtErlBO99IUpY2wKBfLbaEAkBNHdOSQEANe7lC4cOuEZkSrJTYWVyfz9TJUrrD
kO7jrxqjicnqvOTbFefCXBnSwJGcG0zpMxS8GexTtXRobODjQ8eL8mAr/jF9ydPrioXrw3kfiL7K
GDZUdq4wXLEna8xZJyIzqTHT5pjZ7YQ69cnF1Uz1lMxpQT2O4KfJjh3NLWHqaBWK1hLnByS0Ko5t
RX6ceYw8IW+8DqGpJNtiNSVbCP7TdcbEitvvXL/hvuhB+3wb6MoEFIH5lHFRyikanTuzc/zPa85g
/sz826wi/xX++kTN5TcvEAtvlrmn2lSbA/tv0Y7UgTC7ENwrOH9IOC2uqd2OTNK+xj9aE0qbiXCB
Bv5zLV/M1It3az4YoflSULtCAnYPX7EJM6noPkIk3l1awbznWSkB9d+WmO99iphm6bWmUTJB1Joz
zwquqUV/B1dPBFvldViOEVr3Tr5rXxXGvmQjXsmHq5DPsEivOsv6AcPrjTB0HUCG/e8Wls6y2dt/
vtAPp1blFj5KY7IuN34PKzp1T63lBZ86gzGxrJfz+xZeI0sYyD1CuWHRxpxobxtzlk9eg+cSifto
T+CAJCI5PxqXjC2PL0A1b3ec62FSJAf+i5Er1IYkcK4f+Vt8BD+RwqHqw5+uCN5XgNM1LmBjKE0n
y53zEX558Pg/YlqfPQwEVAhFb+gf6DV45Y0f1QKXN07b3+CsOGsyrq0TWjhOwYF0vGRgNCBZQjE7
RlVU2nSXVirGN/buKRB7ozQYa1i2MyM6l8YG2gFkDrHar2hrTqFe9B+ST0rPdPC4rMHvG0iY1ajZ
CmeNRy30+xZ7nhU/RF/c18a2wxD/Mll/AX6+4jttZpq+v3gwEhiUk061z8sUMhb1VXI+z0LuPilc
VABH9d3M2Y/lziH2475ckq+TkujTyFQm4pPqJeuTkUTK4HBYJWlnHzP7agSXSxUpHyaRIM/gf1Qb
aPCo19TNV9qLKpfwX/wU+lDWIw2Q4+uv6oKj0jsZU1+nrLg4nFBLzaIzucN1i6ReV86vwhc1bt3Z
APmt8MH8vyOuBZgo7oaOsqtSgirOx3Qg8lNGhiwKNHqqAjKJlOqXxG/YRg3QwFSEbdfuuqv4tefY
r1X+Ce4bwBg1sRL++/u+OEUm6TOgUO7cbregSB4bPouSwKkLIRXtp2bcm6E1KdqqI2YkRFEHZEqa
P8BttyZOZjzadKy/zgiFo0RfzG2ErX0Ezplf/Qeb7wZ/DXUcac7LY3/7q4w/hd9zWd3vGCW0nRu3
51xNBU0CBEmb6+FVx5xsaXGfQkk9CCeL8Hr3BBEAi7H194Ax31Y0JPc5ziO25Zwi6jyDf28J2grU
yvdVfkHVj2pxTwMgSR3dfwAzEo8Lz++LFB71s70K0NMu4a0rW8fUJkWa0Acx5a101CDL44VgphPJ
/Pe3/IWioYyLjXzRL6do/ncgwlwUVKfaeKz2NzlLkidheTjzMBYN7DHxqfZNgIBZAyJ5IdPW65cI
7kvJNTYLOxXCW0KmWJQD4XW361P6B3TIQHEIKBymFZH7xCQrUps3IkWfcTMGDYUy7+xwPi2aWzZd
PfB2/9fqmuuIufTSbmMsky1Ur0+t5VCun1MizpZ7orLtHUVYuM79P9QKUl7D/+gySnDB0Ewc6u7n
DEUrtixOHvTrYP/n1+c+ZxjswDA8BzBdvHURIOGGeGTBHKOFQD1BTy3Cvd1mINUyURQwXZHI1loM
r9UpZeC1Q3FwkdO/WYJZEN2XLGAerrJAtu3Xv2Ekshbkx9uRO2dOW85X23wCxQe+cqcIzaCIM8Yj
hMFYJQG+HLB9fMTO7lhOJmVIvxPtEdTQxlGEAvJMxkN9eobN49E17MX6Z90MsRVU4oAJ5V3ZoCWw
PuLkxCxRGQMNppEi+YK03D+92DTA4+NaVzdu+ko5uxdwSXqkIutVdWpfGlg73JxnUTyL2vmC9WrJ
ICNHD8KT1ZVRcTlGUj2r9a1ZBaUosqy8bUad+SlzUwKDJRsG1vlE2DQMZCOtpHEXTz/A7TBA4IES
oiE5sQqn0g4OBoThPTywp51+UISKnTiHcOkKQt+xSXV7Zm1n7Lbr74EbzBF8LGogAergNfkBb9V1
GMRVdmFSufhbRXB7nIr00I2OvDRdknGIRcvGMdxsOmD0ku4nlOvIGxalI4hN37YOpRlXmiZpPt3f
Q+nb8KqG7vsing5j8d1cgsiYMRjaxxjDHWw3nlTZlC1t1MbuTUK+2cVJpaC2uPqeTmpUmFAnsMbm
uwUXRlpYUjaewhSXxTjvGG7irt6zLmsakT6PxC151Ud6bhQsTZvmUudZqa5/VCzVoHOi6YUBZE2Y
zjBgw6+2KP1ye95kjirMnMXyMUALviXpI45b7ubuPAlvSbmk2zThfkqe3D2F4kI8jugjTQR/eMDw
VJcuG4EA+Hld5okv+ntj1WY6L0ChZUdRWx+KKDng47x/UauFLFUKbsnawBa6rScWn7mZqZNr0BO0
wy/wFimq3PYY/XpvyIdmWwb8bsn3Ur6U6/0f1izBu9qTvTl6cfsCtJCKQlLTe4aWVtr0cbGmVZkC
e8ooNdSEYIhkqyi/lgINfkRfR5wQqLQHk3HqeYlgXVTp9zo9Ga3O9JKJEs7UsgS7VPHaDcP1I3jq
wPqD8h5svHAklp21DBj/WSIIV8qhRjNu2iewjmK+uRq/zdRTEhYk0h1hTthKxgOfLIa+yzpnfEwI
3NCt472vUDdqILi5EYsiIm5RddmUvCdMF6QrqDNMSIV1GAx14fjjl/BZ69DJaS0RpZM4TKT93KLw
QDgATV9YQGVB8F6pABnTtGQ4UMPHvwVANXp3YyqjCHWPcENPpQvwtZ+Zr2i5q5uE6lcpMNdPUfP3
qYC9qHmi1ElzVIst5z0Ai6FRbJdNChwfpp3QPYl4R9d/iYoEQs/zeHser7iyJK0RpGBPe4zqociQ
XoYCY/fQJbPGBDp6jwkyU5EuVbLPrAe/k83DO+MkDXHzWDtsB1Q8Bx/C13FkRMHG7X3GnelbPe+9
BG563L/MC7J/c+fEeqPGebQ91n/USQKeereOp6xQg+ETCjs6B1LKePxnyGz1ZEmmvN2FYrwG7VBa
uAG442MPQ4T4odbfdvYoPSUSooJpsEMPbYQsRIkW6yGOiMPNjNfIgxwwfRjGME/ytkYt1gJgkHjd
w1dvM890nihTzR2UHSplruv7pMHMvm+Nsgb3R0hbNGvV8PyyR3EeXHcTK8pf20f98E2PgfBh8+mX
dnG1tnXQm0r+o5cZrLJuxO1IBLSUhrllvyWl1swNyWlBSPIj5xO2UiIxx0UJOxPeM9UL4woxdT7j
Qm7AJhGVIb5uOhHVvEyxpUQsKE5Ce5H99buUylY7JCzgTYy37TGV1sT3NcItr0ZrubJYrPwLEBfc
6x9ZlPQWlC+Gef9R3SjBlWk0J4U4j423fk20cVjysaTeNHKAqac/Uo9Szj2oAIhgKDbLlAygird2
xgvR2EBPV+ljIkUqwuvjEDxLbcOcZdytl2PwGzKxn2wpbIqIl2ltFisuEo5Iw/6+COTtV2XeAntK
8X8dCYUpQiGF1xt94uHuykSnSXC6Y45FD54udOdD+hRJ7IYoqIF+V5Z9udxGAZSDWEAKPdf2Glfi
lWkAJS0ufEg+HX9EA0lQF5rc/dFXKQf2HHpxgUgCDymz69swqgzTqk+KRc+9WnYMfg4bu3/OZ31b
sb4AZBlOslsXsqfwxm1V1SdWDpXDN9RhW6vSYJF6MHfvLd6u9lFW3CBqgoD1itky01+xn7Fn0tRu
ytjPwvHF5tdx9Mwvbh/k1CxCJZ6IxrwgB+XIam/YQP0RUP/+PpaoJLmMg5oH9FafVCAM7z7fUoFo
uRuCKU5PmmjUQ3iWFfKrh961RRjNACSR906ShgJpfR1sevZ73LzfmMbchtxAunfcIM5yxlKppCcb
xwXB5SgE/awp6wY+AKrEb+rtCNMnCO00BDr8WNDzvpofz3tcqwSf69S1kVoRLWmflqSjoIzMA1J+
E2inyQAnFtlvF8ugia670U0AJ61yu/tG1YExC934zCbhL7/qMcR/UesQTgTjedUE5KLBkY3t2Y7x
ulQDLtZWfILjrg0c72iqcUu1BuavTf5O3by/pOO9DKmetb7ZPeY7v2NWnHwFpaKeCGWrP6PMzbww
AQsL6fV5O3/vEh9f0/aA0/0Ji0KvWCCyUiIGalplG1SUjq74Cn1STqycYX+UZwohK69SNxj6SH3X
MBw9XVwZvXKM38XEmtvsE4vsSg0r6t14vRNTWijJVGI4PNFfNe/FhZ/wmG3i8RW0f0nBdOVntscg
JfCqWtIWrq3uIUgpDMa8wWlINgvSuy9aS8F1p6AL/YRaRHTTr+AZ+3N56rUOZpCRGDehYTZ/VFOw
HBQToEgDNEi8RNBmnQRowu53AVmGeID1JaKQ9BzjmMCNf9jCy0wWPOKyBJvwXholZHIrxaiaMCoF
qQs6gzgqpLh85qRCLBiZArT/l3n4efcfnoISn7xU/UxJX5b4zDuGbqsa8apSHBxpdEEERESKMYsC
PpyRfMx+E0RIqpM9B8ookkJTH0c7u9Y3wwYm/5IZu6aLX7tYf0T7eNkyO1aB5xE8GV7+RFtgU9jq
HcB78vByRk1p5edVEwG55Qfdxwsvoz3XlMJTTu8EeP4Dicyfw3D3LZXTIuzxFaS88hu5CBoLoKMq
e8wlWfyVSOqQuGtBgcGgE/V/NK+tYcF9IU28kjZLZO0z86u2x8oaSvWQ8h0DPSNLD2UHkEZzYdQM
cJU20kY8GZLlK6PJVNkQPgkbL3HaNNsSiIukrr0D48niIPd5vytblj01mR9x6aVHzU+jAcc7eBiH
eJ8LubapwH5qfF5p1FwR02kMbbt4JMDoPhEEQBJdEGiHdaWhYlbpbc6B5GGeUdTHcTEzuIkaDiZM
mhhFr2mWDOBefCIVMXn7t5V8+ZC89NYe2tWy9L+9BChQiYCmKdx60sPyecj5/SCPiJoAXtEHPZep
WTCG1eOVOdv+HHmYCTIRvY+e1SqykoAr2zL6G/zWTMfzddbGYcoLTIcOxr3EicP19bxoVO/3l5Q2
9DJiPB7Xpr4KyqzHmAtyvYsfU7KYWS4A3GjI5xyBjddPw0/dI5SRPguogrjjR6pwVEE2505XqMU/
Fdej0y+2mSQMr+GOwPx2S8PDr7PcafEF9+DLuXNQWr66XPydGuRRblUFGe8bZDexg/LRywhN9kGM
12QkhqrDLCJ58ywFUVaVi4kawWJLqekKoe0bu09iciC0JJAtKO27iPzC8pinbSQs/JfnQXEQszBB
IPpNX/ebkoLcRRInk9+vMqL3emfiiCU5EKiwIT7IRUgViiKQzIHw2vI1lFZMrAbCWRS6HfuQh4+F
4PAsM7u9I8U/BbKENP71zO5QjEszwvBCu6BpR+oHDn66EvmDq4XEY/TxZbBvb4I0st/eO7mwfOTA
x1C+jPhKif56h46ncoAIOMq5wPZwClzZLfX3LtXQHe5DKw8pve7/ghjURr7OQ7RAktG6vyj4LtUc
f1AeGEi9jOlZuuf6jtaJqaMaS9Tn2S0vCVpZOdXiV2pc/eR13UZxvZWS40XKtiXXam3zTxzWOlDm
vi15YaRKIvXYPNK4Cvja9lwlJ8UeF7nXgSQi2Lckqjuo+prRObAeYO9KEaVIAeoWFicnMmppF4Je
1NmIBHp7g08ML3ijodCbhgtTvD2Kf2wrF/Wmg8KCtqJ9VQOtnj9IZDbGbUmOMDoOfmZWRjg+ZJsb
DTI0eKBIdwtQQzBT2eph6/bPTiWs5MUn458nRRDZjU/t3/d7SBiHDY7106+J2OfHcFJKLt6RjshC
nBRsKa8Fl/6sEsVNHe1gZQCFufUCDcRXDK9xobAwC/6K1UAmgO4jl9NSJc3mbfs8i+TsHgrisfbm
p6ZgjCrJFgkymy0wSE80s35tMt94UupHW1cAy9rdB/QQ7p9fVeaC2rWdZW5uR7Zkq3LGCLs4BxPf
e46WGsATEEze6S8MNYnQTJkswriPboQ60hSizIw/JFfxDNRtVrl1rH+K3g10GPSzNbInsZ5y+7k9
MN4rSjEr/Dhcc5BjcR+oU8L4iH/2VSza95vpw1s+mLrrlFKmehhn1a5h78P16GPr275+690+K5r8
PjAh6VMm1yq53vv23GOQzeSEgKkOttEtQN8UZTbskrw6juebndaKIq4d4O9+ebgf8NCtNiEWfJus
IvBRchEyxUWvRcnlJ3F5lY5SI5gXJN1lAJHCSYfrJrn2hw4mrl9BAhKc1raT74xlF1QwbeEZnSF+
Jq65YcLsVYvBgMsgCtI6K0Npj4gY6KlaJXkv8z++EJCZAnKxF41cfRCm28jrEFxFyoeXxhiizuoN
3rF1VY2LDFF3KBXktrk5MT5if2kBZsyrWhsZ0hPCUKJzZuA4WisTkxX/0uKpM0edWr3smw3s9w4G
f3yKdephRUDKFlZCRanw5YOaShZhqoTp5dwJOCY+I6bb4sHOuIw4SgcXj2vOK31dc38DN8Tw7ZyT
up83R+GiG/H3CpwWzQAJIe5d2xAuKKvbKDHO65kyI/GQokTiZMNrD4nwARiRVZkbQF/s2YZnlXbz
O7GIsFzBgTdMmNqBItR3O+IhTW/llaEC2VNyYKOS0TVAtcEB/2mPiDNEZ8OsUvXWUGBSJwrJZJju
nlDuYOm6icHfQPPImymWbZJQatQ2hYnPIKxkVjF0VuKOLBJdQsL4o3vv4Ay+KQ8/eEcRag6qTkw8
s43pUrU8DQp063ln4hpLZN6JVD4KxX4jUXnswMwLpO3EQ9xE4Xh5wRy9OAM/0Z9WTH1rh51WKPqd
qgPlgg1BDobwE3iQLhqEoDrfEkNvzuEjRwn9eEln7cmCgbfAYSkRNTmUi+iJG85zVyiYv+6odxiQ
+6ddUmcW72f30r1LVeIChHS84Dno1/aVZUltKgRIa0EXk9zjZPF7XdWBLMCPLFwor8qj0yLFxgIX
t453TsJ/Q1yB5lMbz2w8kEvsjSFw4vuicjy9w/ul2/pFM0IzIi5JqwJlCwomrrEqq//N2cPMvn5D
xWpgIqquJ84jI6mu/6fEbZzm5VOmUZoNgOLmsaLXNoP3yYzqZLmRmmVbryJ5n5WcO2rZLTyUnJUV
0zq7hj4YVv16sMtxjwHtEUe1nrVNLppWu95ehMGmmHJFXluLxvfWNoyBSIi0qVMTOWmlTNq48Bcd
w9wuKWTC+QYvXfBHfzjDW2cAZw7NSD8k2JGQvIWRygrw97Fv9q2vDefdje1aOZvZIHG/0NnxiU2H
a/l2ek0GDC4ii1IHYGu8kamtt6bujSUI6kRoiTe44oGtTiaDocxZlWdMINRTLBJojWQBsJ8hUH/y
JTqCPCT1Xs1joqvlUn2nZqvBhtXq/IZjmww0zQc2eTCVvrnyxDd5Y27gOPZ3x7wnpDCb5qv69mNl
KTyjEHeNovNMfcj3P61W0eVk4lMFWC6ZI98o+IZZVa3YZQs4Ntz2OZO+ZwAAZ1bKLJwyhpwxbFF0
J8xSI7uVaOdtolwuZTqmIBF18wqjA9HRaC0pSDYrABBt9WHka4suHWY4hTwHfqU/sD8NAd/x/QdE
gQWxOrXCoT7lx+ZKbmV+QRlh/a00KaHwMRJQc7VI4d9Owsvof6QlNatI3rlqgO01l1CEDOCSe0dC
mb+8M7N4j5mcsMybu6JA/3gxc6MaPl6lZKytadT8NiTLfAFrvUdXIgQak+lrs2tQZKIEzskVmFjc
jGGR3L2El9gjc4zLtUWL/xOk1zC5JWfYK8HFzRBqnVpjO93Cz7fdOasNbGaOSawhqkjIDLPOEpRM
pUw2UMc2Yg8Bhakb9FIj1/EiqovrPu3eCaTkkr6QiG9ZyE51mNpdRNGVqH/fIvxPSs1FOsFJYhS8
ghDm9j3oq/HiupS39toS4xXFDNEfn9pQSEDuaaQcPFhZ6fhbnnNI2faMcQHakQi80J0OJeN1zPSU
q8pOUVmm8DWirpbtt+IDjJoDffuJhN5rUumXNECJQeNdEOUQ3UUGZ2VqvkW5wD2uzpYcLtMJhyO4
UauIswXQ9TMWq65fkpN3v/Fe8y+2F0L5i4xZ7Z6e7+mmpVc7Wi3dzFwPEWgYZgWnBZEPONKD0OLu
T/TMLtLr5r9SeghcFzxbVgeYZgPSUGif8kSHpBN1ydTzjZ7tTulkp5uasrxmT6Xk+07uyjNRtzrX
yQiE2bjUKlp/9GYn8ki7bPy8pJ2Ua5/3n5N2yPrmIsV3kBWUaKe4HcClNUvB+nnC8IPexWxNUzjB
8Gro9Z3igpmk6CkmD9hicDQ9yW+bRgZoN/T41C+EQ3IaI4w/hNgqFXc8RFO9d67w5vEHmJ75zHJ+
+uOCpmcbF0hbbxAh7QydDQHwNjLDeH/vuEz+9eJKOuDnJc6wZR/VAf0+HBZb862vFl1KxnjJa79Y
WEiKRfmgb6bmZLQt+XApMTOCWIWnw9t+BXp8r1kX8d50B7LRxW9KybBeJ/QhxYfBVh9Ohc0oVtso
giY1rNHyhORMPzt2OI+C2DMLx6R9sF72m0v4uZb5ntY5KVgsl/SgG+6KTgb5RO0IesLmwV05v26l
ADDfKr+V+QE0ReyttWQq5mDZv2ce4cXChj6XCSG50xx01w2N9ZvZ39+ZDds+2AKJL/kuarfgcC00
b+vH9+hKimWIsIhE0qesKUpxXHwYupHFBFPnZGDpOKYhyOgjl0fpgixzVR7GlWmT9X2JnN0Hillq
oJxAqjxvE8PMbq83lw/MPHeqCXkxLxeH5aVPC5aaHsH5XPui0h5Ft1o5dgaMxA9pcZ36JuHm5L58
tUxkmR2dptR/P88m6hFbF1dKNHQ2KFVk0TbysjYfUbTQ0SKcfAaAggVe2MjSOOR15SmulmY9rrXB
T82mxFESwlGns/KscKyB2f8fLOS2zwxRUr7n/ytbNyD+dS1PFnQ1xQylncswe5zz5Cmv3LM1wtru
CQj2RGTxCfFjRUjk6nPFfRSRursBRLvscOwFb1a1aBVEWAr091EvmG1wPkPeOimmgTBNNIxOTCPy
XYnMlqnwMKXk8fFgaaoq3wK2qisZaZNyQwBe6nbVUjJ8+miQJSx668OYvPthR5JuiBQSE0uJGmYm
5cmcA7bqQRiNtchkZb/615mEdqoc3ow33p1WGXkiNkNyuiJMMHEJZUl3ffX2YD06ovaVPN8oeQKY
I/pxwxMhVG0Ullh6yYuLVDKfrV5yljdI7zc4F9AtetSm3BXBKT4F1hxUKCR5kuLHnH9F4Ozj3WKm
1D896sVGPBMxVtnYUWPwC8bNA3i9Wd2Xv2Dns1TB+MK47JOQFJ+wAVDyAADRQMYTfCgxi6F/VZB/
MnNuVXNBms44lB5DfHPVpRgMF04dnTopHae79NkuM1Xbz8us4Cwv8NJeZw7f1yf3g9lO5r82MxYW
m0X6NRHfixW/TJZ2hQujnnZ4S3y6KvmZuAsJjXss9UrUpwrDnH93fuW3wLzCrmLfBYi+cSG1J1iW
AUdKXW4oYq1vfRV42mEfE9jo7fZoHAYxTW5A6dQykNRrdyCUIBUsXstsy00m2tsBP9ntPaU5WwnC
8g9RFry9NnK9fokpI6UJ3EgikvJrvMRKEjAUsBG/zpAv2+jV17G2HaMx5vOawn3p3UNczY61vina
uou7dK4Tk5eu7K2Y9KoWHOnTDnz0al68mxlCukz9ThifjOtzURxhFPDwjEVIBPo0Nd5Jtx0ZgqMN
njsmH+HHhwWoCvHc8/3TxVdZ+eiZbmMx7IHac9iDE5IYIhmIP/6QF4Cm6QcRL6VhHhd5k8LBUoIJ
zf8HQpODgRwmV5/QtxhGF0w2GxvNK+vbL5C2ajI0sOEQ7do/voNqTCTzxzOWTva4XWHO7FHaJgQi
eYxrGxuUjhDRXjUxEh67OpTq8oBYrNTmklytMxL+O+gm+vOTadA4Y7yFZAtgPdGVT4FOFLDnKvCS
WHJEYbry3Ofiw9nLJonbuDeZvhd5s2AfrgKOwQVrAhY99IXGOcbXfWPEOWbgNLlkA9FfEG6qZt63
J6LwcRI6Kr4wCeUMh9rUlN/EzQ+DU8o3YZyCnermnx7LCWB5kt6mqpdieQ194qDw1U3vkaqKyU8h
ijzbWMgqPU6DvhcvBQ6lfkwMnJDo9Im46s8ZzrmAA42ouGxcLt8VW8nAxrTEmTMWz6Kf11BQrPCe
cC7U9hRUw6e60B7tmXHe9mTp1CiyO4vUdvotnDEobCXfEKqExwya12zvxlZMxrKGBSbHBfAM1VlC
1t6QoUZPjU995wuO0Gqmy44kqW/29FNQbqb5w0Khy+x/lswqGUgb1Gs7vyV1Kq76V0+WEa1l9NMT
FVaxS8BI6gq54OEnV9fVLzcJfqbgXhmADEtS8YzVyHLcSlcQ1fYI7EbTD2LV7G6UuIaE8leWbmBe
JH6j1dlIhsIkoqdKldb8L2Diih9+q7HhOuc4yJb9hKgRJSoFnHVju6Xpt4JHTKu/z6ReU1nAFuh6
n7TajyAgcIyZ0o7GNh2+Yx0P+PLRGAYirARHERgYRebYlf+THcVoyS54SPXVXfg8GMoTkB0Cfxcw
YsbvoPIiWu/20T/qVWwkZHXJ0QTrhxPwhuLW5uBVahtELdeEfMPvya//LqetIBd+X3Vi8VBKDOX6
zYWr5Ti3EQCUeZb0fOxWt8f83PTz6M38AQ9FKe1ZTWTDUyTRJ/wWbz5xcF9mLU7jAQxdduvHdmvF
YenQPOo5LWjzfOBgoSXCnYqgtAMyFUgDzVWIjdpZ3PBKRu0QNyfH9UIyoDp9AOGPxzRboOeeOXLn
XtJWTE9kdFzUaLH9/HvtBcISiBxr+paUDmjAMRKyD/svSuZLqi8QlMWFNs6CTvXuXQkQTKGbKdEg
U9T1icO6+qyXZm4NbKN8nbcZDWRIiy/GJ8pSEWOqVAxxpl87uJ/FD9c6VdFehZcyzEchn2Q/zdKN
1MzBO/sG1FCQYRGToMjTnw6gRFILs80mL86pWAlLd35lCm5BZCLHxt96Mw155O9qcociyl/j+sDd
ZePYBUJHHD8BG1K8RN/wH4kkZztYp1G7wgRvITGHorVysAGCZ0TcWmlS5N8txetA6FJu16CDeJMz
MYUDZ3Q3uOTnmP6Vz8GBPDTPoj3D90OKjQ/I6oC73q2x83XI4xY2aXJqaMvQs/eGI2MafJ9csXiL
R9QdXULSu9g2mLkediC2z4dmYkOfdnqyzfM/le2uem+ecUXhhLdoL7kDsjF39MomH7zKNSQBe1fM
XYIXsD2Ge/FIunHIQ5jMA8u82tqnRpBPTe3cVdei51Ew5NwCq95YYQEkMtG3HIfNUEjtpX/5V8Vv
EXHgCsYqclmjjwR6PSsq/K8IftRV6we7qIKxELEEv7VKniwM5Tbgv0DWRhVrqG/YlSMB/DuyzMEa
BNyTUlN4jf1w6VtGSh00Uyo9T3tK/kLBM/M6G7l6tCOtfO70cETDYK3FYABCBIvJf5ELJcgYNH3i
beRA1MmsN1bPOwOhc6nYlBw9H6ScnkMk6y/gMPIIHBQr0fhqFYtdKymyLUm1XsesJvwoDWiH4v8m
QN2c7AVzSS6CiMOt+VomQJEIRVHRy8yAqcL9mh3W3lxOm2Gf5AoDYZjNb8ttqUqvZkInyhWzz2PV
CcoIlLKxgIo/2JNVU0/AHPJkBxG+PhwkNwocAjYh5/jAQr74e31xU+kr7UGFQIG565ULCRLqklg7
kDoO/1I3AzcPTss408UUuPkGizAGgvpeyWzoizlAD2pDG864pSzMI0iNQc1TOnmxPfITgCJjd2eT
WG2q1AMdgKJs/Jrdg5DtOkS3qUgZLgkqPsgrr3bIbnpmtIDZaf6vREofnLA5skf0Z8WoK6juzKKO
0j38Xi18rvUxrBcSeXn36iVxJQwmY24fB6vDAHGvebuU+d2PU8XrFOJpFil0MKW6VFe1pZCFComj
zG3/dAXkGpqOhHzcokn7ZBlcABK87c1iKmiYmINZwwIanYshqwrgYRLeVcbcBq/bcKO8IaeSubda
lZnmNqBHTjtINc+t2QMzI+676W2z15S1CETysPZ3BlUDSHahK9L+wz32f6nJhwaa/hy69d4XBts5
JcFJpd1yTKJyNr0saHZkPCkGv0WVuku5N0V2oEjLC4OP7hss38MSx6ITwsY10iXeotSMKE+oMzHP
X5A31rBklXdOIEkVdYriLQXvJoj/l+qwHPTTB0JwH1NOn9vGwRIwr2FnEK521oFtj7wFsA4SGTvP
vz6bJGWiO49HIS4tH4guc5HQt0H6STUxR+BN/pS1YYMGzbPNLSF45B6OcuAJ1yyzHTrKKGe9vUr5
IT4LavVBdyrqRPUZ6+tvgvMCg+jg4804IEyXXosUUKeuR0e9DQfoTbY5sv9I0qxpPOKbX5jgLkAT
1FO9A7FcY9ib22oyfzbKLud2UYIoI3dh8GqowT1TYp6AmyvB8+MwoXq54z88YN78EmKypwlpMsO4
RIIF/nRb51m5G6eaBFN3+K+7PS97k5L4tEYYPnqaSik1Pzj0Vaia0n1BuAyLtgB9yMSyCIiI0yiv
8kQpiEZo0cwMD5Pjdu4vkVMCjQOvrMN3SdcRvv+SpjVxq6Q6+Qr0ch+Ca/XNUZlf/iS8a+xCCD7x
w3ulUhPicprll/g3nTtJgv4B57GOElw3kJg0M14MP19XeY4PmkIvabVJjG1H9WKAfMEAlqiQIwzK
xsFipHR+O+cnu+ijwL0sXBtb+X8FRMEB9AOlxotyWDfb/z7PpPe4CjverlsqturZvp9fHp35Akx9
rh9IitpHuEE6q6faIGK5NIGUq3IMudvveaDWpKfxFpFWsO4axxrR510TJtOeARLptr0AWQmYrHuW
CgLT0IYsf2L5gGcr3gu8+pRLbgKKCJLhGoY1cxG3banF+3vlo0r5rquAjKwYcZFXDVtspfFyLW/4
1jbdMJpAJZTs0uyqfeBqS2CDMJexTUbPAF7JdQyiGamEINdh7HmIO6nWNvX9TmtIivYp/zjyawoz
4v4eV3Viw5lIqDe1NbEmQLwsqs8JhyWvhH1/aqswkOv4hZ4I94OxT2WRWw0ascynsnbh0BtlgtEP
t+XJpzUwqRXKDghokTn/T+Kl56cQGytz9FpamHzjeSgHN+9gVEs5PcifC/gU7zzHEJjMHntZ/z68
XVQXA6fLJLHU7YBCscsgPC7dHWFimHvq+GSnjhULhMKp2xN5IMEGiPbiiX8kcO11JcqaeUMu1INx
Nse/uNAHwmY0AUuRSWgmycdTIIJ+J5TYhYfF+i6mBSZLH7yqAUNCm4M1PQLnAe3pw+n1yfahY0ZW
evZHBTkL7Mr2CHnlsARAxLnbwnCkBwjFOV4g6mdOkbq4Fo+213O+UOlRffLTLiTPk37ReSqx/X5X
09QG3rRaUqRP/vkcnS50D6QjR7PxGInm35/W9aVpciw35XCwPerEcTZfsyngCmC2vxeHTPMMXYaQ
o7M/+QCt4VLKNeVPiMVLE4tkGbTQOzJU1tyjfZDIAbNsNz4uONaTD4x7VCwOhayWtj/qNBSAztLc
7BxNPQfsPumS4/AOolLLnADpMMSo6zUHC+FE7CEyoRcY0O/xz5NeHISyVdvFWDZaI88t3v9Wc9x5
+UiHohW2hs1ip7UG9uSNFQ0GuMTfLWrAA9W8BldKq27bXNZ87N+M38mQT9W68yHsNA6/3Pudu5Um
KsU1yw+K1tvTf+8XlxD/I46ITOkIFrodbx1noI+HIpPmCCscZ3KvgD3js/AmjzSgtu+pvDIHuIy2
zILWztlo46jLTwTBf0ia/+MjDnkn1k3iOwROSZNcLpPCABI2MC1z1zwRyPf6TZH9khTTv1D44bjD
jxnw0T9RxBBB9Sxa30mELM3aYuJAez9yx11z5h91iVdVN84BBEqwsBsaba9Be+FnMrB6Dde7FVgE
PqkFfy0UbaHlkTrLV9NTbKCniTV6sjzEzHVcD2nrTfXzbxqSSN1hpaEX86Psct7ngMf3x8P+goRx
L62yze3/xXQOLB0kcZyVGp3rzk7TOkONZUA7DjavzXYEZqPTWo5pi+1zufcDE/ENvosNK64J41oK
OXagb3hvV3GiElaPZaL7266dJNsE3X/XDgjIBmEVs5Qce2opdWMayDljHgW3suWb36S/hcVJq24z
Bkqe4Ge+DUAjMhc4HYH8HC5T5jn3wNq8iVsf5nmpvvLeeWj4NdL9+SFylIUilLkYUEYOuyHm4RHA
OaQmLIL4ucA4FRmq2zt/N+zbG2yNjLr2AbYT6f/bpTSr4bxST1OikICZbTRN/9AuzqJQRkyu899p
oaWYtEtJgDphGQWTou2aVastBGZ7kJBY8alCORrFjmBzfHJaOcD7fTD4cnqjPG1T4ItlcAu/63Nj
K92WTmDbiCzxbxEJhYYh0hNoGbwyBIUzJka9SIT41B9vwnydeoQRTJSON2s3HMuoUYfMn9QG0qpC
/RqXYWbepk8MbQ0aY7hzeQIwBQOjODxRwJYMiGMX50W3UaiH2im5Gu1G4xqV6RKfpttoDcJBMqRN
9Y6sOkDMwonwg3IMOaxJxX4O/ngg8t4QwLrUuvcRKR3XkE0vTqv7ln8EPq92ut5OInVO2QRO/1VO
sxRVhQPRexhnuKmRjIAkP3W55Ylt9yImU7gQkIk9PRD//EVfq+yaPJ8j5sdpYAEXYYE51HSEkJ2U
mNdKa/HOtiPRLvBJRMo/d2PugQGvk1atlxvjYTC36Di+w/Z/4jWvmYbT1xgweLpyhTvU7dH02ZyJ
0lPcAESWD66EtAMcM2+CfOOsNfDKTFJ2M3omC5+D6koAn2dgBvsDiwC/w7c+9tvpxQ0qo6lnV24N
MUZNxmrH/05w1L9mfPjvm5gnaK/LBqbsrK1Ojw/Hp14jgIDHh49w20d5/mofC+yZGBgXdabYwP4P
KdpZw5pBYIMp2OnepqvYEwg2LXw3J5jzZm4rYy8wrR76M3YcDeSZgIOuzamgJPNN2cTVyiXDYrqi
XK5xKNy+xBVb73nrlxXKi50jGgcnqrnptvJJU7tqkftquGvEVtPXtiPHrde2S9QUEgVjEy2O0N6S
i+7NQYpWYMVJZxqvpIrt8WwAuivSxnKA5bfpoSKGO+9PN3kex7FbIeq9Duke1GKG0aClBBM4gcxe
8XIdK4v4FIu1vLeW0ly8LMUR9Uxo9HNF1HlT84mxz25Cqjp1XUUHmIywjQIMjjAPvRDv/bXSuqtI
7Mg1lOTnPROEyd4H4/XgRsuNZVgPdj/aKqNPhv1bh66agpHYvGmuHvhcm42faA1EMggQzhaVi5TS
99jY2ZBfaFi+vI2RY9vp+pf2WrUbG5OEqBc8MWLJLSsnF3CZBNxfkq3z5HRlpbm8XSZGFf2fogVk
eYu1nsGE6MrOBTfJisMS6dfbB24I+4rp65K9CsHezqvYp41TDf+QS27QOJTn8zx0jv1TufYAaVkD
JFzAhWxb2btY06MFTFlGq9nMNhDA7ysjFDB2/WSuecy80geVs7eCbUx/bqpU6kbFVRw8dGeiob0f
yMafrtrgYucU/x+MFoEsPC57yEkYLStEUqjt30JhyLTIanCxvGXBs305VcupNvxrd4ww0rCsIwnE
eHcjCsEQIxlu8D/kvdzRPyhzJJHH1I1iDlD8JBEEQrwSLouAlnTK373T2GLsGDtfE04lXSXbfOKX
mqiJOlt3360IpGSBW7SwuZx+i/eqlrw+JsfxnkxblIXjMvuGai6o30EL+oPndKoiGDk6B/pDpCtf
GvT7D/RbemYgN60EiJE3crqMlvD4nkuOqFPJ1G2DyS478G8UlBLipwaFKiLE7Wwh5acsHyQNbeoj
/s+l80UEtdZDvGyBBKriTXd2NuoYuUKMG6MP9lWu9XfVV0XHY6JVPTwFC1gMknB0mvyxnkB1Ntja
em4zdTCTpCrDoClmC803fZ7mdKiWoDWTq9iXjpHiFvLpvm2Aqd2V1ab+KEo+P6FkQC39rBKvEV7B
zkthHBJIeUDtg68BWnU+Hufe6oZbYs2ESOAh0ab+xlgpQNOA3oFMpvLktTSzdWYzY2dSD0XVFrb+
Ad2kbXtW0k/9xc0e6lAkRM94liIHiiuSEr/zd3zze8JzOaSVtsY8j8xsb0VlRlD18E1teEE6hWk+
oHE3rcgMshew0QYgVAPxSGKWU8G7pT1t/fduOrziaNasa7YtU6rF1Fy7h1ygo/wJB0v1KzLKTj0z
3QbMM/7uaaQd53OuBTrONpIHsY39bm5pbxVq7U5DPmACMXneQ101LpNTUMoV9ebFjEQmyh0lOut3
bQCMOtPkTS7jSv25zHiC5CghKB4Gmi8y++xtLfIZCRvnpQ1Bm7T6DlZTk3CWoJi4C1cH1nkDw8yb
Qs1dyeIa90JrFGlbf6STztXr7vjj8/zmDdNIJCdaC6ksI8ussK4dgwjxa8XIfXPI2zBGCcKcFBIp
o7kGyNJAsAknIqclI6p3Cl/2z2jYDj1GC9uHPoqwDhdWdYPxmdSKTKZ8XSe/jz9KaSG12FHVeqDt
8aOYKSf6njlenXJnasqLMSakTM/XDiQ6iUgzslvGJyFJdaxVTyX3qTA57tkHkdQp2f1V+PYIjHV2
HeJIt4iVD7DWOvWbxAu/uoNaLC9NrJElozTq0h7FbgapxLqM/nxLMYmABCCeKLGm2K6jp+f0DAAe
F4Z4RU2K2C5xXl7KTjGNpFTZmfOnUknlP71OL7a2SZ3Kvn1mJ7+VBItgkiSB9ya4ygVNsmXWJVNK
hQoogqhcbpCAMa3y1gTjLiteeoBKFc8hcmBr7WkqRX0WfzAlyMQl8az89iSb5C7+bPPta141GRQV
BmVxGmOkNxq0BgtgclGZsOc8gmKChWNwkP0X0vWD2UA6O3YAvGedl4IDUY7ua2hXdKfMPwItO5IM
YPs6m5Msuus4OE7HWRCXB9K4G6IcZ/hb7oXAXJiDuMpIFKbGuSq2XPOXsH44+YzIky0f+S9IsjR3
yZDrLVbxc49TO7RIr6C1ktE+MEAw8TcJnZdj+BiLJBmYuMf1OWzNkCEL1DsAdvjdSI9GTGi9sUme
Gel/vrhqoo3+CY0T12EZO7MWZ3M2k/YZDamWAZTuZp1GyQS+HALC/m8RDOIny5RucHlSvnqqXTSy
NMV/e0algfNvjWBk/T+cLMmjae46gG3l1MvNrHVxRveiIRGnWUmY68CY/SINLTShJGfUZjw81nv+
YKMrtM2tC06/uPdFqeiiQV79GmZ7EBI8MPgGxagqwGIv/0pKw2wB0lcphrpqDa8mdtulNLWhToxr
6Wmjc/IbrlKmaqcEC+zS7h8dTnXH/4Ffsj+b7L855lKGcvjRGPC6s0zfB/tG90sg+GtYnDhpKMvD
JmhYRiWibRxvqZBKl88Pab8wIIx34MqmkV5t5altUOJkbPycyDmWgfHVwlAAM4VauxQF1o7IID8A
S7qhkFk7OmL9AhEXtPDE1OUC6p69oD1o8zqajlCpPMTzFuxPoFj5ljwuUzwfIVufoJxUXCBhXqy+
Wa8kCOMhabvkLl+jEesbkYfGb7Z1DaOtbtlERm4BhZt60gfg4zLKL1PAWJIyO0pWz3u1OidiPdkS
+8teo3Q6oOSdyajauxAs9Hobot+b+c+YJYUoi78ez3AdRUiadGzb84VHrfUZcabx45ItLcD8LM/4
cX2teL1pkMUPvZa1UCfnBk+rOwiUrMq2ixk6WW1EYpABz6nueJMGfyQsQVNlrhwWGuXLE1XA93Ly
UR1Vss3a+CWSQe+rp0xIpRCsDBz+e7F8l2c3E42DaRSGXaB/cxD2LrtiWfYWb7KJbQPuWavig8j0
j7An30gtp4UUn3qALAArj8G3F9uexlEG8NggSQ5kqRkNB7UFTMaqQogkEIzqI6BEK59Gc3jlsLTw
uIhjTYklNCFdDJuXA5hKdTplMzxOQO4pCZUxve6AWhZJE4bMPXW/oxw6cNXgZlaINtNRy7fKDwh3
Af8qcGrDqcrJxwLmyfMkN5Z7toIt13PIurnZiAo3oHlQsSGRNZoNikGtZRscPwMuZZI3pSeX1fDg
d1i7Iz0xg64A4e22DRdea+uwHja/Ujlh2C817jFiuq5yN0N64TiNaIgawv28yj4rqY5E9pdtvNZY
1XRBApWdEyPriSeochT3eHFPbGMvodkKdUqNm3Vdpcc1Z6+cPGP7TPW29op9O63S3y5T9WWoaS7l
I17FQETsJCtCOw01LyjqbR0FQCsPRjRZ/RVaGWvDjopelSnDE3Tbf09PAw2nSY8ITEI6K6mUArnP
i0KbN5JYvlVKSN6btaR73vR3lNEcruqB1EvEE4QA+J0Nz94RHZ9CaWOtwh9pm1bDEpqLL4JcRVeg
xiZYWDY7QLFZrlrChmjPPTfCssAUvMOJmSPLGAP81f1zmpSTVrutbDN8bQhIs+kvZsmRMZYtPjoF
csiRknvtRjXi+VryPKCaYLF98UIIxNCdE1SjlS5FOCfYA3Ga5ffmIOxlX1v/jLkOgJOyyjyK3IG5
NmF3QvsxHf3fJRpEJethwbN3wh4RX7w6e5KlfltygcSfvL+7A9r9XKITFnLROH/DJlbKGjiyZt9D
VZMChVWWLwERzqwVvdmH+Lu+t9ZZ9kdlPm9v9OiJInwNVXEiFWKgujJJJSD5XbboEcjJr2OpHSqr
7svmYpYu05t76uMjq8qdp83pA+mmXegnvPrXe4tC+DEEpfhSu/p4C0byok7itvzEkQzILgqtJ3KL
NO/IGjR1BmYGyGTbOVwKeXhGyO/KI3ppRYedKcbhnvHqLbWX6NdVDXqscbWn+TcNyNLyk15yDMfr
pXarRzt9cMtDqRDDehW9xShtyLPN+H7lXw8vlp1Yd4rfv/QWuVSQmsSQq6AlO/K49564j5RkINxE
XCjkMDs0CF0z6Cba42l6X43JujGTDfubqVkzK6t5eJw1aNs+cdg1hUIVhOuuE4XolsJGVXjjnvNc
ViWj9BKLC/QU2Cxz8E7N2ZmEl/9RsKx+srvgn/L3TTrXcqAwhVpg0uCTWLVTluwfAD6ZtkK6D+Ac
gvaJ2bWO8Qp0RSVeBGtwTsFt5J3yavVw9fZuRSrULk3r9gMnbXz7qRf5JMekL59HqtfdQafIP66F
eIOJHSjrM/0GAcfV6fcGiYI8WG0tLF0ve3Gl/IDedn3zof2s7QkJOdbAMkux4poGdhqcelGdImhv
T/fk6UlWgLgO8LNwQantMdMyz/61qHuk2qAfatflV6gMhWQRSakZrntsg/jp0rx4pD0WQ+8VcTdm
F2lqpaZqu9vVnMnRy4IzKEUqUaxo4V21Hjh74P1bi3Ac7nzqzPKX9ApOrKFmYd1VP/qsidRMZqFj
taNvxfmSlf8E4KL1BwyG8IuczEFG59kUX3rXkEGYSskybRgkUwQ5o932P68UHfDEDUrBDxTyW311
ECqNDr3v1wS9dhAYmOo5D3F7vHKOb1EvSwwb/f+bPvVpUIgeLRS3ixkv1693aN5PfC11nAPPFGh5
WYEvl2wkn/2rG10dNEPqaLTwtfW9foso+it72wpSeJPk5Gr0TP7IqgaTfdSdWMAoIurcqcSyxrid
76Gt1F25NdX6U6Sw0RRCGaR8iOV2dSZt1DomYD/vIHJC3f9/LfouLch9OKKhU6jVhvMzUJIYMN+z
XtINsUsVh9wrDxHN55Pep8Cx7o8MOaCIP8ZGVc1fkpjSjdWg1MzhOdC5NgDelIucK6cS1gbDJ2uc
Ek3qEbuen2AckVgWJDFZftjXRluEon0CkU1ydw01ChttF+yUThJadFvpynfSzZJ/DmmvwKSZ5/Y3
q/NtvTa1n7bLpFxgivMYGggfAhmChlV9+voU7EIbxqaz/h3DxxhcUnf1Poj3h9V7U2pReoDclWfw
eXrC9mLeAqG/ifYnlq5CFhwUzAS5FVgMWAT3vlGbQYsXZLpuGQAUhgJFmBcOGSgDIWeskSnF/k7O
PRBweWXeTv/9t05f3t1DV2P3UUJaoiFPogLhTFn6LhYnlivtr2DONQ1jbrv7peBCy/YyOlzrAci0
bhIxeJFTa/jvsAwQXujEFyFPVdvnNX87O8Gjs4gaKWzIw1M5OGD0UmK1MXzJFAEUCSwnADOkYLbi
41zehTWGV8hvDyKd/t5rSVKmdjAbMsnJ9+0Cmrl6mzpP/Bv3So8r4IpuugfJNScZC9mkiySagdWy
d417g5nPG/li0lr0cjcGxcTZfl89ThJN0Yj1tCvpnHGFpCuUJkTlkdnueBnqHcslhPrKF8tjAipM
kDTyCJCnNOYQ/oN//eahHB9+AZzw6DkAXoKRWNck60l0OX/2mhAZIG68va9St66peHcozwOhI2Yy
wWrLHMR9+qDDQJ0oWkHhN5rgkCMsydQgjbUSE+v87bwhBW0LM6i692QZRFVYrxikfoc0OvDlOJ8Q
GQ0zLTCUOioLZYR5C6SYOlcfnRx49QAXn3YZeVIgdjAxfv7sMI4hghkd0UtD8T70fGj98XNtL/ZQ
ZDJQxr9IKAPRMDG9IjDu5pWA9l7d6paDlorrBFvI5PmPxbK3TiLbQtOb6V/fd7S38u8vJ4HlycsQ
e7L7eXA44dCDGSh9Fir7SO8z/WJ1XVkDIL36IWBeCB2FfqRZxBwGK4+25H0tCWliLnw9eNzD7Nhu
y1SEDEiVG8G4iOMV7kUXRbRDYsrXkLaDnKkGPx9ZNKq5Lgow/8TgxpRWOfHxiyIre8N6H1Cei5ca
LdyZcFzhxQ2PlU0Pn0CVE2dFx2PS57BKMvvyZEejCbydiRWwYMlY8Y8lE2Ocy5Z0WCL6SV2M6GIO
RRTwMf2412tZAQ1a3ZArAp7k9RbhpxdkJqW+bH5ipiuJ9vuW5q6cW1NPKXDFiIdo+AMB8loE2rYf
68wJVcJLJNxZLVBKFrlc91q773ofsW5SD1ChXJPAUpFdrirLaRgqh4Fx1RArvQ8G6zyfAY0p0/kl
UoXVC+UV2IK1CBXfEphrjmNhzMyz0dHWRRBNOa8WWnXIOfCiHJZlubeu6IDEaeMzxkz4WEJkTjC0
gYQDl8Yc0eLOhFGbXC4kqW9/lPnjxQvvbvSUdJl28uTzPz5w+TdnitsfidVzWgrWYRmMuf6Dqm54
OJL4eQHGDVEbWVHq5Fc+JS18kgEqo+RhuMAwlM6El4igsMtw1kVMTvNG07iKaf2NJNqEy7pobM2k
3ZINePLJpd8Bc8n53KRWtYd+wt6UdQ80MOCvTJhiQ2GQ6srkb+p+w231dbl/QSPbWSPuNqPsSV4c
J2UNvWISv1MK3gQRfhKHVvbvLgWRNaxHtfYIpTd3Wue/3/KoUKzMDC9g7ZUqV/fxdx8EYo3yt+RV
GN022YRnJEcJtAkV0ie4XMOGGzGC1ke/VEpfu1X/0Ew+gndAOVBvIF+r7HyAsiMtkg7HKAAUlidX
Hg/cF8vn3v8x7MvIoBW0+f+uppS+bbPpa7KtTG0khptdyMsgbjLY665y+HeywX8hHpMt9bauzwY0
4ndoS2Krw+6KR+hzzdiiO7ytZPKovZt56KjEaIL7pRvyv5fSLrnviLaMyluZxg58AXo2Mg6ePYyX
IKn5vcmUxMQKPi6bOJwf8rRZeht3UzSI7frTIN6eftchd5oAcjAc+VpFTF5Q6OMGlMn7dBV4OTjv
t2234z9XC886AuFFV8lBeN4Ux71yKLQAY8S0JNKBgehnPiwQcKpN+HVJ4+mwy2+1Aji/EJTDwjBO
ztwCWnnEG9koLHJn4Romxelih+128duF2hYkmMHS1RwQXowphYD4UCghBvSMiTNJ/oSLpmRhOUdH
3QKgLpXupoFkMoqMddS5oOUannTqZ45KUjZ6Zfz2uTij+WTNoDdyd9iW1XKUQMoixEngcuY2l64z
EhVv9qvK6/vf6zg8LMahP6pN83RSQxgqD2BNiicDvl6fh7sv5pTjFP4VHsrB0Z/vW1bLv4Qk3tEQ
rmZpPCGpA2dE+/smyWEmxpntGAR1L+Dw2YWOr4cC3YCQnHP+gZ89YcKVF4iPgjpPuaPUWa5BcxKT
eAU+QaIS1dMHtScdKiHT1v7SQpm3JrhrdPBy1ALPkbMmQgwPfD99HkHDlrXpWXFFfUjyyOdkvwIa
W0n1xCeUEddya0yIerje2CXM1Cm1bYIUrWgNQGaLXvh8w2WteVLbcVAYKtf7N9F8Ys8Bi9yJwGcF
I0I7u7WcCj7SEYdjyQIT+0xm4vpvDnn2ZW4UB+4Gl4HWRtKaoEJ3XqLV4mDuksHCUowsXgi1ca7o
Yi5wgXHLnQr/pOxa78vM/3CwM6gkT84BuW1tQoRBOIDX9+C8nI678s2uA+NyRfjG9YmE1e+CLhtj
DKQU0nMQjStGX9fqFh3FPUzXHh7yLH+7pxKs0pl6Mv/DPU3B2DkEL6y4CodKpHRKOxFqUVn7+Of3
hfw2Tw1I7HxNxOvn/ZZ0dD1a75o/NpxoRWzvp3spMZdtmebAYkCQ6CIx2i/qvozGLjDRHp8hMsGD
Aak7o44IhjaEPDM5e3xoGJyiG7yhPqh/+baZlKeOyp153FflxWOhcmh+2SwIZ9SBdC70MjB/dzfr
dwtHBJ8ols1JYD6WnvwvCbUdtnDWkOyYnupIWfp1cchEPnLWZzoxwUemTSWWyhutNCRVaEdOniDN
HaugCT2XogEl4zHDaiWDoWq5EJGE7mRnP+FTi0c8htICwkciR6bKmkdpM6vGL0M0m83+hgEKsru1
4GSjqSymkfNRFBqyq6M+gN7SsCXuOwOPG+al3YJNYGDyrKh76yKDY7cQf8uIexYcmYLYcLP1WjWy
tfohp6PPoZ65alW7IrJ05xTFHFB2YPOHAMo7BYfV+Dl/ZDoaQY0zRMQXmTXSZ+c+sstuO44fNfso
1n5R8qhu4DyldA/rdaZ1/JOtsFnkIqfxzfq4lEoDmMjTcjKizHW10hUiPD7qRrnvU4x1Sl3GcEw+
Mtcwwgr7qgG12D+emj/SlgGdSlYyU6uGhA152e4xwzz4mcmKha+MlPIfYB8myYMkotmsKy5Ec7jj
2itwMu6tKL0PqKOTsYOTKw8kxGg1q/HmDeSRFp8/qXtUYmlFj1Np30jb+2bl+dgLd9g7X6x0DTbQ
L6fAi5WxB3KrTy2jMR3pYxJThoQsQGZ7/MTo9k0uF/CcVzYZ5BeF/gLUtO2Z6XiDy15Dl9AFnh6g
r66EvEpn0ByUrrIkT1hhD12mRvYo+kVuJrGbJAqoWKTnS3O0S8eA1+V7bYxfdzWrh+9F1GMrF5In
WEi35jpriCSrrZ8ow3+LiTQ06jyaIhtv54sXMRvMKp7XGh+n3kojOqQqBFgvEuKTGms5GRtN5WK1
jIwO06nejHKn7CDzL5KDzkR65VoRsyWOF2jihucrQV4k+qrmZYYgzAW3PprQI1c4JUFSA26oePYt
Ekb3ZTuKT+cz6CrCe2HFViKC/FGOSTpaxSCQYZ+rfFGr1g5KWz1+ss0hODJfknq0u/P4VESSOno9
cjnrFTN0tLwlSm3hKosV4d+Zh04o2Mm38Db3LqgE0s2j+GpO7oFR0vwZl/0oDHcqJubEnNFpS50E
xPar3262UJnRV3MP8mya+grxBWoYzmGFsGaLbQx2m0GsrnNXFk0oM0np3fyARD/HtlpdLdKcjTAm
ukjJaZia99ptIL4xkyTwudmoLssoyNhC+OxksZM0TxZIAWXiayG9rK/EzWfGF+X20pLN/ZEA714J
LvIu2omXvE0qoGic8MFUho0j9kbAgnnms4Bmy5iOJgqc26fsUGnCOqACvX0NT0WUiUbQU6FHU2r+
gesvvbbywc65jlwI/nVAkGXWxgbZ6Hm3gD8piKB619bK9hYS1fvQ846vqO2N8rlMxnbR3Lq+v66/
Ds4Oh03ws2nBFw7CI8kyI1uRIkamfvcq1M58mKeaqX4Qtci8h6RnOHTxB02tPlipjXWnNaU5kxr5
YTwYUPV7C63MnIVlFshMSiKzH2KiQfdUbgcQadTOM6rpDGDjNhP+uy9Aj/+qUrSTagZmlCSgADLu
zfhvfM+olzUitGn6ozn3CMoP9cPKIJpJy0s0XMhHVGBGLEhRhnGFXX0h9in9E5hgbKoJhEyh7MjT
ayse+xcCTykezWo8ikqjfdR6SNpXUniZozJMeKb/ta4SbTJKP48it4RkfOdCO0PnzvWodH4tfyU5
OboLhSupcM5GeXgsMtWwVOrfunHamWnr6DFcvEIpC2B6GCGbNKJQsUn5uvtsBbEPqa8YBnMEn2UC
0n8dTvWQXx5e+R0Gu5ewvrWDWG6qY+ujNnR2TSUNClsn9+4/A5SpuRAKLe45QVizJosfpN7H82m3
VBmXpr12VyCM96WqQDqtDBG/OuOBbPZJx2C2DXlpbYrV6Vl56oo7St3cMI/MH7NN5ZR5Jn6S+T0i
gaHgOnyPmzumpiXv1wnBMYZMVTqFh/YXv0N6xYENSj0sao4WUKEOf5UdIm9fA4Mg87G04gcFqffr
sOFQF/dwYm218gBFhNi0RNRoA9AGxFbZQID8X5hOISuigsIxrKJgXoh2wZqRQ7K7eJIqUNH3dpNI
0IQtUI4CbSiHMaFLD8Qjwsk480CQE8wfPyEaLoBW4Lj+63SRRVrRljO/W4fNyBKVEpR9xJ9FYFmU
reBWWneb+k/T6tkWi/fBMAe8J9gxGEMP3hjp4Lta6eu+L0JkfN5yEGp//RGXwT7SnLNlSmT+3jFI
wIky1HB4WHG8KallRngcvQvjOMXfZelzXfb4jsedkrbh9pM6iE2VkAUAjD5P/Mvr+zJFDB28PjE9
ydnN46AauELl1fSmjaz772a+81Tjp18NjEC4TKdrczI0bv+07R4XQHIg9UvRa4scBeyBuwoORDIy
CFJx+39N3940fXe+GjZ2TIcTXEU7Zrid2yz6GhXEskp8Fve5ijDFnuPesbQUVIXHUmVdPvQuSzvC
AMzGYsQhymG3+tHltiqTJ/DFQvFI/H2dOZE61rIiHA+9aYNCaK78hCR9T0CGsOpHbGG8ynTvpeK8
vzdpztbF++R6ylIKel4ixJ04q2ZwjBpDgvCdg5bJC76QvYCmzHp3rBrpdk0SpvtkaZ/7EXxlNhPw
4HoGUjbMqvc0nhnjqQUlY0nn39OZC0w81v4D6x5CJn6Sfqh2vA4W+w+tatV279u2IFL/kc+8Ve2l
82zdCjpKNVPOxb0Nac0tFSvmitd4ct3nRP72bdYRVKREzfmNE6Di4BEF8zCea/JuixftfZRVTxN0
fhbAeFnVgO0k0SI19C6hkMpM7o4Wo+ERl4LX2RU6OIcPGMTg4DXJ4bPt8smmArrIYXegvmIhu0yq
PpPofK4a+k0QtCVBdOi5DFGZwrXWo8UaBLFCIOQ6W8nrPS9y7jcVa5p29uEbtreNuiIvMkdQJoBS
0FucIJ8PkzD0jsW/FkDp/1pNt8Rz13wSRrpqkdc/MeXJw/nDg/Dh8eL026i1iWcJFBy9+Q8QwCa3
yqzqFdvL+Ny7IQfDXaKjdjEnN1MewnUmP0voGGcdPeKXbfbZJDl5h4qMF3c59TxXnlUpVrjYws5+
3/SoCiDp9Gg1jKCiB9GKZzlKqcSGamrRqgV6FjP/mJDIups41kSWDccvr/GE0yZeNgR7zjdOqd5h
RFk/zJGMl8SzkXut7Xo8PMnA0q6/VQuQl5hxacBAQuONX+Lean4VLsatMqLcn58vy6qQiEmyxQHz
mxwoGySBsEO2eokB3a9qmStJ6XOXqX2hvBZ3yjZTKid0DFz9UMTeDNVUDc8885MLYAc1BPsopCLt
BtuZ/NWRucWj82aaocV5cGbpjQsRDrSslm0n+27xaXXXzQ4i7u2Jk0/3h2E9g/OCBkD8oPOtGUTD
LJ6/FdecWjqqvCR9JNpgA7z5XullxEEomDM3N5CZXEFiCVh417Tp6KtuU2s8kthMV3xWEIZMqNiM
cyxDF35KHdqlMXIr1tEqA7nWU5uKUqFLnTOrWHHNpaWcDCEO6c2DDfNCOeT4dU+6TfUHKANvUhOp
U8Xq2r6cueaekVp+mtOFXSdrMoDHsl/OjWhJs/DHYpu3DXyUddusHoLPeynsdhYhSk0poOhV0SaO
yh9yQ7HIrKttMqfpEITkx2SoxDr9ygSbQS+3GlHIdQlW3YBhFme1geGm3c/9cfZyUb1ICGvUmzer
BoRXNu4lMbJBDVgYbiWy9MJf9uC9GwCokHNlteE1iV0N9aMUwraXzPtwm3kOephLdzLwPTvOILkb
c+CGLeTTPGlpfJ3JrryksjLZLEqRkdVJXkgdOBB32khZYRclllcwj+TlV/AK14U06vgb2xO3TjMk
YT9afM0V7sZXJzBDss6b4MhCWXmKQ4z6cZCXEKbkPQQbvk3YtHYSfmwL6BkhIsspcMpHCn7S3qpK
yD8Y308rI2v/bB1vF72m70gIjGSu+PWy3Kd8vRwxgPsYQBdVYJc4C0gXsQJBnnB+xltaLazJLWcl
hzsnZjrozy2M16JXtoCtcv7c0smqJM5JP/1soQJ/jDmDom88B104BBveDbxCvdAJlhSofHKYQOlo
T6Ia0AJCUeDGDvwrj5n4pI3oXipOGNRCugjQ7IoLOK3T9IrhYRA3XOVBSOr0frj63bqzKElvupe2
DWtK4wsFVDFYZXJBi25U25G9ZgcPUci2Lwk6jA4iJR2pBXTSKDwrb+uK4xMdvkU1nA+MGsWxgT2X
mt5zD9VyMjcbNSGto9M1KnENJI850mnQR2pKQB8PfWGrAZigeMisUsH7NnndNwg6ENl52vnx25Xy
1sE4VKYCL1yIm71FSKtqN2xJjiKKVHZxEiqOXhGgeIUVBOM2iu5lV1b/qhzjTfh6h/YNiUoApqCp
Zgu2rXXZqEcUAtc2irpZOdTovy0OLlDFkBvbZvuQHAoN1Aia/8qTzxlDnv0U0LO5GP2a00eUr6sS
PNmL1AUEmNWnunSd52pziOo7BxioW7Utjh0jdXjpJAJqLoDYyDNwWT4TJY9i+CZKr8HvCMwwV9lA
uBeaoUFJY89QXXz/4gKN7aeYTE4Ug1Ze6kQ2NYhh90uEIedErGQ0GUeAUKGHv8ub1qG2BCbsjGsW
2r+9VyAXP9wDTC0W5GllG+MzRubKIWpoKN6izoDEI8GLJUSN/USJ25MzoY5BeuHWL/pefG8MOira
JL1qATOtAI9zjPKhtJFpcyZddC7m6DDz3oKFSr6hwH4RyqbDGfQTUNAXf+VKVh2+xjzNQkj7CvcO
92yVS5V0zLgTVW+OBm3HkIhiOvEuvM/Fnh7vyZm7sAIxonHYBnKhQyIfd2i43ywoEUHQUfZbTNql
6QKYhu+HvWPYDaHvKM04Eji815dmI26+xgS3l6fufNxrYM0z2TCxGokMBNCFPfOi1hDdPATAdMda
xc62vmTxiVP2mUqszW5zTEt1ASYRlQu4xUSyu9qvD3qSZutiWl8ggu315EMFyUVmBQo+NOBcN/ww
XjMrr6YaF24z3uGjh+KStJg3Peve33j87HxrIPEXcg52blR+FU1P8EXDM3clLeSmoNGmDVYvwfEm
cPEARaBa5refaw18qat0H4SNl3Omfd5fFNcAmw+6JsLF4dmqVs2lgkwd9fieW3KUtqA4dPfqTbs9
p4HcHAMsv3iTUZ73waSZSoFLKCfgrz8Ci9Xj7SXxfZy5gukA1LBPRuawT4Qgnq13yRwbpi0gdoCv
nfMbcO3E9OagAhNYmTOpwST2U+vogHN6j75b3A8694FxHE9NCRY48/+WENz/4KDz8YH3mMP6QWc4
JiL2k4FLRk+jVLpdIkCQYMOYhNHXgRCq5+L0kppZdiKRl/P5yQenjMA4ZQhKckfUh9ReM7bTXM5V
AdVmK6Pps+l9rA1vFvJDImo6XRfDw3cq/GlAwmZGR4U660OeV64ZmM/0ru/7p30HkzEBm4CzTWLs
FD9XdpO+lm5253L5zs4YFXd6PNk7mapFLFihq3UFI5tyRA413lh/JYyom071k5oZyjXTkwJ9z9n6
pvNImInp4bEF4/e0MuUZH+m9cs2MQLD/dF5Ss4kOH3QUB3blLp0O4fzfpEX/dNP/izxjJsQaOUwj
M7pG995QkIIUJS9tg9+rQkZ60oEG6bfjtGGbtLTAMyH1UiRn7XE8uYpi2t1mk/N/qkv10gqjCG+7
lJ0AQT4b9NuZ0CkPDMMS5e/afqvTtMGy4iYY8R/ZCt6CRj/DGvtrvX2FtKNuliLICQF4/2WumX4h
OLIuwIhZH6JH+ZPYXpwUtZKe2Wn7egClqBviJ4pK/CxBBp7Zs06u2HoTUWNMUo1pUpCAeXLAgr6r
K7gW7CiNZyHjYBzd7BEHr7BjxrzuVQprKpmV+P2liCygEveYfgxJsw1dvEDmIQm3FPuxszAMRmL5
I4ZdpKPvx6L+pNRGMGfYvfshTuzG6dpUFtLcmwNbiqLlYigjZkf/wZ3Np+4haF1uYRToQ/AfY4Ub
7aTic+Bh6hlbocjDPnWYU4yvtgwStzI+U7qaGfRflO9a/EerVRDE+i6LXDGadHfamiVGu4E2pb63
ccor73XSnES4Wg+CODCeP5USohHBXfvF12TyKXcqi3JmOk+lR7BDTGOjL2tHb/JPiJ/XFJysMlcF
UfTQuSQJ5o2z+rYqcirGNtbnAlPQUmOJBdMZeTlena+OS1E063cAHBTH7WJz4xi/vhIAGtbeJDfh
BFMKfgaqHA/Yd/OnTPcC8JdoZU1pVuFTzhHnroXqQtJyA1LUObpOwt0nS04bkfQhfkfUdQdzWL71
7xrwF0gB3I7yTVlV+aDI2YE9cf8KvfC3R/esS/47trj14ffr44iuQa4/VJclp88RWi7/AnblkIWJ
/Q75kz7t+/XsBn7HaVaszSSpjuJ9G5JQp7LWq4QLJAfeA1xISd7lP3kReOMK/gdZzEr6/87DKueS
cU60VsXFtIh9kOgNc7kF8Ys3z9rKAnODkRB6jbL8IouPqMh8+EOSy6EOz9wl2h7ocGbDAIZcYrAU
PXFiU3s+ABZaNbrTOWZb+0mp+UDmOkZFAP8SdDZqrrkcuyRleF6jPj663BMfT9Vn+cVkJnegI+78
5qCzyg/TpwAKAjzi3ArszzXnTH6dUqasr0FDTBPn2LWGxrd4duBhVqyeWc3Fp/YLtmp10Yh8ku9v
8nWHeSnvMbbztJPJ7skGsfdBcTvHMnD1ZDaes+YLr3xT+IUlGk7H7Q/UvqPBItNb6HH3hBL7DgzY
n/3O7iO1zboGomTwQJvGlW6jhY0jLS+sMvRqItBgBfFmXRUWqUxDw484bMgGOuYSkNOm5L3kiwBr
mxgvJWUD+g7/J4hMeknMiCP02g0zaBrhL4p7C6L/bTKD86RJkr93e+yT6Y217+M7WYlnZl+UMXjY
T1aLbulixTpdFkKO/5O20L/olWC9fPksd7VwQTzRzvlSuyOZWOYgzyJtHWsQ0BoNb08aVwbfg2eK
2FeLyTwaaL7koyQ+IJfB0DIeBf5GWhahor3hHZTI9nVgUeLg2WIjeCrJwWG5fydepSnR3Cw6kLau
pPmN03lGG8g/mOhkKencQQZlJk6EVMBhc0EsLUYA7sbZMvSr0FTEpvHrm5Tm+1moe+r3MZD6ckxf
F5aWQO7yY47BFJ2pxeMuMCMpBua0CJNhNp7u2x4Vh3gHnlRwkMSmQzeohEwlV9ll4rtMTp28UYuh
RmxYe+3arFyaKiydwJjkbmucPaE3Mmqlx+g48yrQkz5fePa1S5nhDrqaG86BUlB8kz4MvVX9VUhK
wkqzoyYWiJyi71PMcSB+6HXnDWizdSPDfPOZehP4qev4hdhrw+DJBdg4bQRtzSCDsBq2WG2wIya7
PVJRyHwxaEnxvJs1WAwOJLbnyKrmXxJRRtVlHeFkJrpZlvKqxKPjCudSRsn5TWNA56mT7vSrL2kp
n53EwDdnIZpGsla+ZCi6P4bdoT6Zu92V/iIgvTj39QcVV4YSM9uC+AmuZvQHuYSnu/dqfVQ4mvHt
o5nEHelu3bJ4XLSwXZnYFNnbJcXAd62baJRwCwqEbNZgWtKZWGWrmfw3GECqzWDKw8Um8haHiER/
E+T1e7Z+15qGu/1VeIPOX3xnuB+haDGeca6kqmiw/R0dv2Y2oTeDLLKqR/84bqXzgAUkJUnpcdUA
4Z42vDytaVI4Be3n1cSUXixwFPBPXRjgepQwzIcnZjJbxat7nLSnw93PVyAmCZwwhlT/ChGsITid
Zg8TzT/C0SjyYVRKWAIG7lb38OF409PJ9GOXacIBa2cjFOt8ayiRx5bZ11+K6lGtNX3LSod3XWQ0
UrcheS4qDgs4CLqTyueZFWYOSgavj56T09jTkDVJy64Jro4eIgVjaLRA7Yi7U3ZM6FJvmsM/boGw
4qEsU4MISOr4btkvG4xcU+a+0ljN78byZA3z9NnzJ9dp19cCHiQlCpw1lZ2XIHrryrgYh7v+eWvK
A8AZov6qtQs3dibpVOWjWEoCsgg/lOY3xKe0bHcjJ2JvYkRimuyYntn8XGrks0vlFpyirDSIr/Kn
XIZFfp+UBUrUctJQktmEoFuEeevvRlFPsS058APQNEUV8l2i867Y4bx+JsSb9DBwB8bJRuSVStYc
IbBJUoJ9pNgVDZAoj2gchgbi5QwMJShVabb2BQly4/qCXmhWWqTh7GlzhTc909tt0oGwNpGMboFx
i/6J9DJ9FYQJenPBdc1iEBQK4qnT0mjgsgZpei3Q7yXDCBW5zd1mr2gClDM4HajkKrBpRqRfi9Px
5AKfOQEPqihWll0vg1mKIwANalywqFWA0zC00J5phSlNQVCxLAV/2T5dCraUUOwfOaBfmyWZBRur
m/G7jz5ZDoipjk1Qkh2nIN+Z//aym9YyNfP43vKBQBaOATMt/CQkMNt3nmdECeleaIUJnLxGdHbg
Z59v55+e4aSnIuGukTRgd2Lk/KZc2Z3cQ2FOe6TaFE4zm3BrNgK7YQ31EYi2xuU3TaYuyBA7oR/k
8+C05aaRmX6WZ/T+tAjU0I9ZI6jIyL6IUlDi1CLQzJwWrIjasAX+AsK6ICzwn70HqspvYPPrTFnY
EocdrzIQp4OF4KJG3P5UByarqFUrSoHSbnWKnhTYh5qUjTPctD9hasal++q5dskuUzXdoBlVHPJz
8lAjt+ToUH9fXxFtQPTsTMs+1RxR6OS1P2YagKRcMarpcLyC/yekOo9zylAEcz8o1B1R51RZsNpw
eNQcKuOoGRNmGDYjCJd/VK4zOmgdr5GRAT4fTPjVHCBzUHK4qNNYdjQrhIZYUgVUfzT+BhV4Mocu
ty37861gZ/Io1NcbCFEp0xPKjaM8cVCqdnZT2btzHgX7CwmPFw75zGV4CHTqL5zdz83xGjYUS/Xt
OFFC7Ex80fL+pR4H2HXWGObGxbC2M5+5iUYV3xoxi1hEiFYyzIxx8kztC4G8XFdmp4Zu7ot26u5n
jRMtqkAOz5l0SSSnPDQo5JAG36/o4auO4ML8nWJ3Xxj6gskTpGAf/RAR9YsV0v80oCtuSpPWTJKJ
kpdel5qxo9ru4skwe74g2lKAxdWbeCX6LZ71Xx8AgLyYwUamzyv/os0qakEndDGbbQsWMGpIRQeK
a3jF8iGq+IQATYaZkTIWDBjVryyzRvLwQvg+P5QLtEIyMN7MfNQ5mZJxEXcUdSaqOJ6+xbXCHM6V
3ZYrysfoxl769Dr7y6W3eP3CZgzNPbnDDxU7fPPrK087ws35yYdA9AyTzHPfL/kfigSR+Ll2TO/x
Qqn8nYY8gabEdt46Uu2Qgjxn8AFqi7SJW18QzLK38BXMqaggYDeeAX182Z8HbT+2ttApuJFK3PFJ
C3Vhv5to37HLPrlyLvGhMexlruW/kxiF5lEiD+qEBWDRc2z8cIgSRTXwtwTQQd1YPTR7HSVMkj3J
H61LlUBsIRNkeer7d09Uyy3vltrEdnXWe4ZPN1j+aD36bklAUDPYCvCMn2U/CI+dLaVKQ45SRsOs
NlXCzEWHW82iiRWRfJPkxH8YbcM3aE4Qj1Mh1MOU6rhckupkw8nWEiaJhvJXSdiYwbeiqC5fHkhS
X/Kr7j1R/RUW4VkxZFol+mOFkXOE6Ne3GYB0iSnSopGFNmP7YlAO5frAEDaYzwKUPXPNeDRZb1A1
N1yKc08zgcO9T4e2QxDytuzxDhNqKQeRoo0dldS7PHuAOT5goDLrQZtBVbje97JIuoGPwImRPq+0
rGl41FoeZUDBtCWReMZgL0irWOOgpVPjUiDDTrbfU//xluHQ1YiHeDKi1iIlQX7B4G14RHHjKPtv
8sdL+BG8S/3IzR2jc7PeNnWxBUo2I4oAi65W0lyNEMy0aNlB1lzwBS9ToJfXiQaL/m8DPggZuG6+
3PY1R8L1A2lG9sa57OxJNIrI5AX7xS7eaZVuoWTaAPm4Q4hXPS17WEMp2YaJNVHFmK8vs2kG5E2e
N0vXhzIpemIB1sOcTan0d6jPXCTeZQn4B/3SwCqUOEWq7K1cBhJEzRscpRuuGCy0c6JHJcjKRIYq
7XzbmInojwphZrKEtddPjJeTH815JRj4PmOgzJnzdO3tShZOuwBIunAza1VZ/vuY9nycmU8oU2FF
ihzJxi9JLTCA77bH9o6HRb7m5OUtxFWE2/gsL/GwH9+RPVWqCvhZTM6nSN9pKJLw087phJkPqDFv
E8bNgK8TWLR//zVszWrWigYcoFPPEkNDepvCpuGidGSSOH91I4AwAE/GFWDoTnbg+qT592lqNMcK
6EqlpIlUuZQlNwUd87P53ASyilSWCN+a6uPNj7ZSu5gvZM8ebtZEeuf0hugrYtDDwm58wVrGz60Y
zhCnVCdXKZ4FWZS1P9NuRFeA3ox0eZFbcVBtFuVmJkVIMFV7/jKKQEnx2vLWogR1tOXbRfDWU1X0
n6YT9utvoEm2PImN58hjjcCHzhBelLEedAo1zxNCkFhIeIOkfgo5/x9FxrM1JT7ha2CdBOaULC7l
qJhKZBqaQQkVK/hqFrBhcCPvzxZeNgP3JivawYIVONy2HD9rqFqMwk5soEOYieo4JcxOjuAAt5q+
Y7Uvd/UOHdzcC2sD+YokKkcA40b9UXSeqfwDCmxNskgU2euMuyPgf0RjJvVyKHoxbEslg4j4JMAm
TVNbYlyAOjZoX6YQXNhahGULFHfhY5ziLZ1b8u4WvAnhbupNDAOZW2wtsGHPus2NyHSlFM+By39v
L+OmoSV/hJZ6AluRdsrzDrinrPMvmzJmQDZPXLQLqzYqKRQTFu4AjI+gQ+44J6z/HZHTQZzPOr6I
BeZte0KK5o6iDiaMwUh/jTYUx8WUa19NKKNbPmuYdK48owTrsDS/NNYVqgCVlaBWvnhMe6ZvvpUZ
KQ7HQXtDBFw5PaRu8PCD/HKsi4eVIzSwypS2u/cnFI17F/8fDTG3mmC/UyTcvGen2667Nwds+5Bc
Z/8zdAGMcIw/BVw+P3IRKhVFnGd3L5moQ/qPwnhmLbuwLS2plzi1B+7yo+eLSWmhe5SmV6geM+7u
hx11UluXKgOacx1BDoRB7guw+l8PqW/UvRrbY+M+vz/Vqc0XNKsHiqu1qZYR/XY20ucK6iOTn5Y5
Kkjp8tdPoWHEXoV8PRN1shsHpS3+GXDAWYCRYdM9whfhtEHSOCTH5+3CisuKVHDm/n1z5QP2TPnO
3OvBPItBmych9u5WRi3m6ST306DaCkRgSEgE0BXOWMaipTFSOC/0yeMiCc5rKXJAsX9Prqpm5HkN
NQLVdpowbBoK1qcjfaqAp6kM7KDUcetc9QMmsHWSqFudOTq5wlDkmmIlzO03Ld5ayKCkZZMpOm9+
srobWf8SBRbKbW2KDBqc7jZlVtEg861Hs5eAcD0UPi7smehLssBF1n1nrz20cLuQKuQJU8VV6cAZ
1HeUEsl0UiGA4hvB8NkczTGiTraJDA7MuH5c/RuF0qi2ETU5dadtCDIZfR7065sERymBdv9aVkxQ
crmAsHKGt9fuM4uCfdWKuYJY9lqofNVJUcUZfdHAA99l9BdBBNvZ1jGI9lls0k74r388kwIdnBBn
7UYqbr1+JXc7DfzgzvgleWsX8BSgl5Ufdpc+pMySNe8iaR+Or8Oe2mbEk9jY5v54aWwqu129n0iI
twmTMZOkdKcAozPqyztn2s3tCaHPRW61H+P0SkZPC+rwRI9SvECTiVyRkM9tP0X4ZSXdhG+sWBXt
+/oyAQQ/Uf5RDW77yLOyRJNOAtCiXBbl26/b7h7Ucgkz/fV1eGS1xHh+SODPaT+gyQicSuU03hnV
GWT9sihSs0fFSZC3XlS+7Lh6N9XsPgYQuKNKESaPbex0xD2aA0SJH8AkuA3gX5QTeUaV9n2UZh22
HCTQLY7S3qx4dvjdW2lvUtEZAElt9ZrGe3row1Csf25etv33s2WJRp3Dwr0rFccENJcbPtJWz4EV
ucfd9s6Y9wBBG0yDFPAYricNVkEzusmR4O/2yRNya2jVpddd1O3hoMaEVWFLSfJoFY006UQqAB63
q6Uo05AL8m7rvIQIbI/kGYp6Ve0vr8f8CdbWkQD50wGOc6hfFNVmoAX4GGdaRriDHmhTVSviCFz+
woBsv3JBT08BnmTGFV1S5/5RTsz9TDvviCQVCaPqCOW5RsHlHzYV+OKClACGYluC9M2ouibgDSyZ
fYMao4IY+ob+I/fBp7wbxRmBS0uijm4d0kZLwbe/PD/20+Gc04f3Mw7M2MeRCqQcpyZMq68ZU6Ik
0/WVL0Nmg5htxApQqlNwootrxB/IamTk4A8+lYWa7JUuhPPMdIYcQKwzhzkkY+OTx3grsDoOnfGj
uSlFz5UbW84EnOD4r71rY+7ctB0ewxPoUX4WM93ZCNY5amb8OZ+N++Gx1nYvpHVIHSOzKUDt52g+
Ksit/BAdAretNAeQT+qWyWQUkq/uyty8Z+pMnBNq4PKS+M2g9nuNwQjwAQTxg27N/4X15811PTDa
fXGqTbBiof3Hwc/b4uq6UUIJ0+Okp7GlQX9SlM1MkSSfTH6Cn0a2RfdCdog/1jP87d/gWuKYsRuB
wMkyl6muIfmQu/5ElEGN8cmutYj16okkywZVGB9PknnSf3HlyY4AilN1hn9pkN022WRvO7Mr9k2z
LqKK1kiNYWYzKm5BV/im2pD3NY7vg7tx1GadAtYAu0FqarZGdyEuXsH7yVCwVx3gagVg1dj+epFc
2I20H4FV2GT4uMQokcI67SYguYK8zMyi9FWid/Xe20wZyLpQAWjdBJ7Anhx25bSK+qDeSAsnVTa0
6C0ewnycG7MTsLjy3ZUQXTag4UKVrLd6koOSDeT1+IxtHFsNEryVma51JjsXZJKePOqpFFROamvN
Ju2rgTVOOjSG+hLjkG7jfzXkHLg4TKVQZlnbTdm9TgC3TGYuGiUEu3FiJnlFTGTl4d07aNgjOL6B
1l0Iub2AWbaodD6XsrAHlSLYiuBINUHz0+2934I++HgdDkEOwBoNloKUlJxOnaTZbCZRKl0R5MOz
tstS0NQHZNhtlNGfRCPOp3jtW/x75IUdBHBwCIwq/5YIGQGYRe3bAX4eVkKvpPKmV8JTZzrqmZ38
y7j+6kvQ63H/V9WL3KPTou51D8NPGj39krasrVJ7cHoJZWjIgScy/FmMCDcYfidutldqZqTVr+oq
3C43M4FfouWYZ2T+e1RtFVfWj4Xd41yDCX44E4dI02gMOJ85Ws1g+l9MkNnKAbMwjD7CBMCQxO5Z
PxyHjWDYg4748MD0VpHR8GGBx/+tWbAeVcGj0GlWR/22hu/Dc/PBUBBc6VFSqxvMxVCf1gDjn1F+
4cVXNY2//UIdYKCt6C5T3upV+gRIY3XLDYNIQ/+TC7xCyK3LtsRvrlKh7+Cu5NUevvWB1d02nh6O
Cq1y8E8tRUSVIB+qsOZjOsv7KqXlvJ7zOhLNDzlmGdjDKTgfGWC2ugqg4G+fJoIBrzpFJIz6GlFL
9JHalxh3dLVdlgJ2Bs+odwtKu/VLt48ahmSMK9KPKGoGDki9H/wmp5KdQ7OGcaNbPvS5JaXjpUMI
oymv6iOxBzGbAzLxdLfOcaUrso+rcOkABHkfCEgdFB9iiHv4O7Xu9NhHRJTqJxKOUrh+u6/e/zmC
HgEm1gXR2pi74up0k22OM1TD9OP0VAXEFFfu/lkTQoumVrFHAYUpwyu+TEmSxurrdeqPQZve+S6x
3gfJ+XehyGCvVB29daVxP7Vq1KO+0/4V4xN/TLI01+rRCqzG0B8egbELaB1fqTulN0GbW2nRCn6w
3rcIYA0nLD5QFvAvlh1U9+JrN350iNA32ATfWHCFGaDzguzLt8SCL6oQwV0n0qPXxoOBowoldqnP
z00thvRVYxOlVCi0aSocYU4o/lKNqBwd1G8wUnkDs7V99bjuhAkcNkvOUNkJoJVUsKObiV+KWYo/
SQcjs/3TMJoYq5yP2J7zk9w1D1e7vrLGK/m0+rP9APVy6hUN158F03n9Xcyy5IG4rFKHLiGddvRd
N4r+CwsgFaNOtrcG3Me6Wnq1cjbXNSQKMAmL0V1mYHWe4hzD7+9J4QLygoZzzS7mTCPWt++sb33/
TNXLEHgA+f0KAKMyrdkBkm2Cb0dJoKWuHHTMjUbzacWzQYETPH2RewrzbtQnt+LsK8QrkTkkLc3u
wMJMt/oI4VuAAAMpcG0aBtb6dRSQNDFkbAUAXtOh+MqPt5ub7qZHxfccm54z5m0Q2xXftTDNZ4sv
EZyqLJnJIncXznWK/36O0OhX4Wd3JE2r9y2H9oChlPs6m6NxOoLW8dTvhwFRpImGBlJMAaiB6Eva
KpeCXq/acfsbKu4LFB2bxq/568iFtuZ635mRofs+wm/ginwTitaGzcVHxmJcArz7CGYtJbU7+yZC
pDu510jlNRulOC1N5B4+AdBV5rRTUpg08oEnhSkRyzPUKBnJOXPmVOZfJo9ktcPGW9Shf3WRuD77
qA2jdxKgDapplX/50CcyLI01wak1zVXL4Rnv5++Ti9rCe8KcWZrt627qCuJ4Cho07W+PbUjL9eSl
nEIJfZKVptp9pzM/54I+5RMNZQli8WDYAuEVE7M5I7n9041L9cbdYn50COYHSpMlYtsw4SJCWjGw
xfYbcP/bMiiUGRl+cpmH7uatq0UgbkNxwqKcQzPy8qz2lm2zhEYt9KE8b6TTgOWFW+V++B93rkNo
VaVT/RlAR126DPIEoN7k2kqhWHsWAAVgqpwBiH0TrMsr+jJhuF8CdpEXvfY7Yga1LP/nPqMY7Isl
2PpKUogEanFslGo8PXwhI6gb/CXjieXeasQ0AvKgmfY+K7d+jXihKYjMwwd3MHXZILXs4EischIA
ESUzKiDBqxH31lRkeZQt6FsafPy7iIHx4weeXsfjDZb73B4u4vNZ0qXCOkWBGk/WrXuOGX2hQyu6
E2Zk6RTSJnzvWx14onpc+Of5o4gMt2UkDWghvj1C+ep/K0xWXcJqbktFYbTxEwdECWMJJrURjuoi
PTqxsEPifF5JPz5FVg/bX4YHAECL+3uBEavgnYvv+wqEySU5K0OM1n+8inl+UBmXMueq/HkKWFVM
LlGSqpbS2U5H+z/9HluIsT/wKIKOoFfEgamIeEQqvI4bXMXoD7jGpER5edZiUq6vwKMQ4dGAKmie
G8aoOlSyL1BEuCbqd4r6kXBLzxup7L0zhollOnV2ao4wOGEOgH8B9SXMFSTfPoeX8c5TtG7jrLI6
hcusTKvk1XAZ8ZGBxUvTVdPNn+6oT8ljgJnZrg3MmGF9HiFxl4KNerYg7a2TiOOqrWF6NdLI/nsO
pqfA361Jt5Mbljvarm8vjZ1EOC0mFVDXwtORvq98e4HuA4TXyafP+gO7HXi+SdIisOx4iG7RJj0r
Siqc+lcbx8AO3HAVzSRFuJZBcWfBc7VRzfS35racnYmw0F5SDDRkm7/GnXvJamU7cKoag1phCY4r
wlGi4nrfuoscSz6hE2/49mj66AYH0ME9mGyBFh2nS89jRXUciO46WnaVvqUsmYx9AU7TZvzPxrl3
cJT5vi90k/DXr8nmZ1ndLwkIhwp9zZMlbMi5B53//swJf7pIaMP78mYxPEKz+aLrUyCHqS1uO5U/
JM1cmcFncr170uUcKJLAiFMiQ0CzUAZpsmwEgGyJe1cmR7flC0CASD6arGTstSg8F8qFIIXq+3D9
cQEY0N4pjBmNRrWJptuZMHkZd4D5IaXWBwOFfe24F+8ueXLceFlbNb1rQ7RTQnsfzbnhsRlZPclP
SFgP+wxi4kqjOiK7DIvQg//6CmGxB6jKJzDC9RSblLe9qL5TWeiFwIuDyxTjIXGFnPZv9t6zr6NS
pgQlmBtVIDxcxBd1bwIKKcwiAV2lKG8zntxvAuJk5uEvYn1C0OTbbfAMY1vuxOmfV7nFS6j0QXZa
xOjbTKI0qGuwUg5if81kkHO98GK8NS6v0LZVaDW7t73v26LN+ZAFQAv9D57kjmiTAG9o3K2SSUpz
5QDHnGU7ZC/bbxtEn7NxrSZTtshwgAwU5qaPYnJQk7hMWjpw4iHwhmgXP1tPKTwI2sYqBd4Elpwp
jFWgd1A7gXz2JilmEgMutlA23O0AUDOQ3g/wV5+McPB2PJ4faMjpbAK70bkkspUdZIUKR+OsapeA
gEJE/1GodXfrrU9JkJaQUF/G+ZGGuHbmb2xw/UfWmjNWAF4CKKOanMS+eNO8RwNA5k9U94vxH1rb
47yXjFES+TmOHaIiRCZp3tCIpl0kHz0vvq4BVmiIMG31j0zE/6ENeK3C1+pylCZr60qLS2mUUIpr
3XVyxiIPCbx7/qBg5bSIR57QjWDcKrvoKw0EyXmXE0MHOcSxJKFii/EE2ZEKHBupr17I02lv96pp
lqQ5POMp0oajl+b3tKQcfQ44oXZqgCJW62ITtdEbagMh1fezgdX/2nAanb8BjCSAJEraX8CiNkkM
JH2qmxAij33qf7WwE27oUvHxAKwUWuhS59YPH6VJmZb7T4nNX7Z1DSWKNomaHftn4DcCs/JVnH1Y
+uIm2+E857qDkANcWlinNZFRYJlMkK1bOk/VmwS55oYyqzF1vYNX4+OLaOaBQQ0uuxmj+0x/IBgX
z1PgRkS6YK5ZcmjMg6Vw3+m/Q5BBXXwWvbc1QVOKA9zkTsin+lduQpP50IQA3MROeE+H2hSOP9Bc
zBXQv1e/hNEyu+ifoZKb/Dqp/yCwFoNxicD1aCWRMgSkv9JeBR6k4jrPePH5m1kv/IpJkR0e0cqv
eWqnk9RYb4ECsOxQZhWl9y2CKsJb4DQUDH1VsQHG2CUoGAqrXR1MOwYWaS64I7e/CuynAq+6HRr3
xwHOsl/YgzOedfv0teQqC/pmAVHEFi8k2EPDsXKH/JiPpjPIZvJR59JT5zhv9o46rFfbarQqJT83
u6uGYcC/gz6Yj/f1yPElh8ZNLuc8TYGMIX+EsojNaAyTzmu3kZxQ2CEbh3RwVB810u5EdgqpQ6bA
bCbX/+8aVRYVTgULV6v8A64QpBw5+iMqeZ/WjqqETRS82dG5N0KyK1EvZZraGoE5c2xlB8rsv2GL
Kpvg/QoMPqIhHWGV8rcQjxQMrWA6rGsW3tPDuUC9OzwVH4HCMeGJHEL4Vz6loao00OxNMteXVHRv
frEiU1l0afjLAco25n5JlK5MMpMDqr4nnjmzZF9XNiTdL2MycLTnUhLJWyFQeH88xnsq2ygjw0xZ
sKRELXHbHvWXfpiAXGTbLqHpLIOOqQ91v4PoKs39uTTfPmnLwX7N9LmhQEYKT++Oe3XykEQfRuG3
XiVZy8iBBQDn4jJf5MiZpKbOj/0K3r3EZVR/zPO68ZpXy6Je4lvOPPoQLHROeOQaiWKaiwSnCCto
dkStrRNxOZ1gbr9PfXZeRJdJCNLVuz+8sR8QSKA5e9Zd1Z5taAbuHPh+j7rGs5isDsJXz+L4PFpv
pIIy8qxdc+6wEvTmLkNYpQh4xK5G+6XxXfRhWdDyKj9aL2IpSfA3RabU+ni4IEf4z/MyzrDymYAM
95LSaIIppd4DJVmk+3GHBBOFjqVq+4hTuaw/GLUHoHEO+vUEKMxBhsVu9nG7XJYns5vKdKBM7h2z
PsVGatItiM6lVlEs5e7R6dMCTSQpfeZ35nch5BQtqLPi89wVB5D/2UgYi9JFb+oOOZNjJQ8WO/SZ
u1rqbS1bvLN5Qxuj5oYDJwFV7TdYG0wlRcKfs/rHlkRHUNuEyPyJEzL4W2leqh8e6WEE4gpB7N9s
ZiHTxsIn+jWzQk2eJl6pDWVdRdEvKNR7PIWdi2l3kswT9cUeJ+JRA82xh//mW3n4OK9hTd2iDaCe
l1fI7+t3hUT066IRANqp8rajvVhsqWyf/3hJQzVYKETEP02oRAd8waexubRyFWh7kbJfSukTB8g1
iFEBJzHMVdpzrshDnOeEMB/5H9CB0HxUV4YY1XDNTYegLVRg8vRRrYePjLcHd5OGIITWtYKR8HDk
/yviHuPhqhsszEah3s483Zvn5Boz4h1ZNK2jKlBkY83gH6BujN5ti3tgKWjA8QryqAgAqVFYKyDJ
9CN9cjsTdBz5NML+ssZigKJnPjDucAbXZB5EnsQotcrcnorSEiXGkubCCEJQ6yNvWZXwgOZ5UmUw
IiBiM6N7NASV+4uULKCmkDm/mdru+gkzM/Mk3s1sReu0mb50u4xh7T+awZYcZKJIhJof8BQqKLAL
vajd1Ax3DkWqrOeuGzl2IWpWYp8hPckrl8jB0MZnE4GuH0OQpdC0ThgjTplCxJ5yDe5X8EepIquo
HFYuYrrIIhWs7N3NDxr7TYx9snPX0lH92ph2CqhCc6rW1tAn3W/vtUXwF1Tc/NSWGArtnxyonNQ1
48xv1LZy+lMBwE+ZZE1XeR+4csz3/2Igf+n00cjZMWotLLbI9VHyTfjUmVoa9MsY0fx9+nNYyQSR
MtWmx59OuLKzoP02muZYcKpRzNgLYAwYNCi19kMNO7RIh0/kZ1Uclblh3QAeUYttYNvPGR6sD2U3
bO5yuYR95oizt7SW21NGIQ76RSVQD5Nc0lm3gqViO5TSojmP6LzGjTk9iMxKquRgAwAN5olc0PD8
s2suPD0oS83SHMtxP9eIp7vESwsoRUXImLmgIDPZS4K79RlPgZ4ScjAACUpDRt6BbBbbocCnNH2B
SYViBIs15468EkBeF0hG1h1JHRFPh9VNFvEBAOXs3vvfITz3ODDBI3FgRYTW0gtAzn48eFqwoa8C
fdIKgdLZvNRcQQ9ivpCDJI5wFjhtvMWA9sjGkYxcZnksdEx2K+FdO86is27rnbGLtuQ/dXfYYcEf
2+An84CHLw1u6xxAN7x5ahIPSV4UJ9aIxfqJCfq/WBeMVzuBv0rcohUntALr0pZAlOn8nZsZoHcL
Hvk5Y5IKY4CRjHBCnwOxNMHjuVA6yxnJVEE/G3SUX6dI4r+b7c5SR/H6+rjM1EBaZEsJiEMTD8IO
sLVBv2YIBPczT0oTB783xzbWdwcTJbK9q0BI3u+O/kehdZlmISK6u3fZa60yH8AjGw+nN7IAAh1J
dCQcBbO64fsq1oOBZ8Ae303jE8pRHimYkg+GHm2SiQKvWUStYHraVboN/SZEwX9EkxnwhJciqKPw
FDhyFiwxVzoxMiKKXll+3kUEjlC1YQ8BPEJP4vIUmWp2QZVgsBYHJqJYvnXoYHnF89m0mox1m93y
YzWQTvtAFlFwF3lz/2/KHIePO5Lou7q0+u+YHE6E0Vj07GRC3bfnkXACXgE5JMJvKi25AURB6WZl
0iEGVYs/7VlFQxSLi8Uh/Vc9OB9t50OgZWbu3lpE8Ief5MAsfBiZyoFmQ0igsPzbRpFKJFYxR0+h
+hHRpT+/8UVF7Fqm0xHVDzg0XFISN1n9fA3gq/9Xqne0diAAhShSm258wFNlbbSxncQFU81yGMsy
SPPd9YyrJW6vaBu+ConwezA71YTV0Y4/SXg1HeT3Wz/LUytOUsp0BPiA7GC+ZGq7dSqD1b8+xG2X
hy6tjxZv3fQ23WFhDwQRxMX96EqL/Kg+Lt+qgNXIpeCByuALlMZLLC9sY/bD3pf9x7Nt5/uXG4nY
qezzLj6BIUriT/Jpz911YToYyXjkqhBdIRidG2Oa+Nxgy7BNbfNrYypELqpLPHq461OxA/0Ym7+t
sXuLKejZeOQNam19YCfa86Km7h+Nbcl67B5cFtVneR0T1HijSav0OEtmcjtsmrss3A872R0yiw+o
NEHBDM45rO3vVtfO2PdDfruUjeBwzdUulltXTKcBRfAoekHzMREtu5SxhULHhQ1AhUAFe3ocOJc1
AvQ/MAYxAFlB35PA02PU2knjb49F5fvoo3SLQ9cUHjIL3AXQ92qjGsEAtQgTmjrXVmTAGL1kaNDt
KTQ2pYclBS4VGPPv4HcJ8/yVHl0wdctLTp1FRUEYQclIa0Dz6F8pi2a8B9ItcY5xqMFBY1q7X/yx
owaA3yFChqG9OA9bhc44qyHXTllvUM/2vjiyt+yd4I+i6DjV5JEDOxqhO4MVTx2ZdF0XNoVEKcLG
XcMDFRFDT/FKGBg6N8vQ+V/nxdBGYUK2tfq89ysFOebZSJLef2K9LByWkpeWppTqH9tpnkDUNVWt
/D5YZDyaBIC44v7R1M/Qnl72QhtcB67zhMUCWTVfi98/lurs+BJCZona45+ZPojdtAA4TztaswAJ
AqXch5tAg/dJn1sJ3lNpgqg8R/opj+CXXCcF16pgCWlZXSPywDQZTasIDx+5r7DM/gUWJqM4inDB
lU+bf1znPC0vxm+u8SbUli8/1bIhKaFqx7aqxoxirmZ9gGHRGKvCHPYwzamjPllM7TlXJwX8yISC
RTngumXR4nDPcRPhMidfJT5lePgZUklniI0pKi6RFqdiQmtOzWEOfzG6sKOoQbhw9HV1tWMMCmcX
eLGz57bDnAhvut/vVaVq70njacNJIwy5xzU6CHdVhOcJdxfsdRTRr20TkHLzbs31QEDWG+pW2KVc
Z84wz2W4wpezvLeuxOCs16fuxpitofl9OzpDNKY+fbKZ4ZJnt94W7csF8lCztq6IYIoqPXKFG84g
gP8UMxfSX6CLkC1Id1D/ZxsP13SflyiAc6MRzS7sxTKJBFP+qG7/N1LE9bKY0fURaq1NmsF7NVIM
M2kI/hoWFRFwPVo+PsgF6y+7EkwYOOOHsunBAYHpOKNO7MAG7tBMiFzHcUv1sfjcWJxp3dawBxEV
CTbkUWBDCuiJkAPzLQ4UOwZQ/rG1yQr0YGBAujKQ71eODkSii78C/66GYcDRTiz+KsuJlNqu6h65
U5lxrVIN74qBDzRyJNzbbgorcwJOuPI8bhwdCLnkPEp7/W6RWmH5JEUerb3cUGNBqg6uz+8ZH+J8
VTwuStXJMkrt38BEImIfGLsnVW0ZgtTDBFoScjLqzVCZ4+z8RLsGSx2J/NzpBx9veQpghZFl0OY2
SsmjrDc/te4mmYx+S5+iOKiHyfgi3jVkKHCYA0MXzEKUhrahHOc3naRov2TO7L1VrRqKJ/X+3CPw
PcpuRLgmTdrs1GGLL0A3JRFCXRmBH23VNLiAdxSyJCQx2Gl2M4Py02cjzolZa9wtgKHySZfU4gwm
MorzHuONfBP4icIiH4xqAL9n8q/ewS0sW0W5fXOAN4rKYboQ07R+dKHKEcDo3m42BMB8s0WLM6vp
cfDIKJsrWkt9KArxLDUvbI+Bi7GqI9WaF38YJ1Tk8fQJNs8Ou0/uH+VMIWx7be4ZUScSaiQLuqUi
UuuOfQgdadoxSnifasrf9es9UrNVZYEXEbCqMXLboHOCphxr/AcDBso+y2ZZbAy2gcFLyFWtev4M
lkEt6T/mOSXzMnc9yX84OnOX+Ahx22Rd5fxJsjWKid8KmMb6EbkNV+H9tWwuIN2JC6jeYvd5qkzp
Ttf0b+jAKXU+OYfCHVikLUCa/8tvdQniMaRebqF00Yf1tPcJ+nAH73pkhpfnPczALq6tlymfFkPp
zBUs6g5LoUUk+VPIilcfHJq4V+2CkMsswkFLyamc9JXaXb7idggVEr3yyDficrL792LCBn9qUFnT
ffBxepxw5Umpt3QHr3hrNsR5I2PrE9TqGRLS3/fk3nayxEBq7P6a9SWFFvymsN+uWGvdLztLdlTy
i2YzRzjeLTu4LhrAIXVEGkpFv7BWp8ACFc+YMV53FjiAYbccX/JjY00edcbxjljtLcGEtNQGGTka
ZAh5dAnO37LOlVAJe8fQ3t+b2NQAxI7KK23ym7cdRe77q4UkZEtBBLz4Rx9lMoqMKvMnbhqHFT0y
Hc1fOTi5Ap44M630LmE9yy3qCbqYMZ73X9cCEEiKaGneipn0RP8HPyHvMyj8tm0uX1gMs0KSXHfh
zWQi3O/AuOi3ainXIJKfSTYVU4epqVx91fPj12Ap/m87VhYsc6dYMha0jIWPEpMMn4zQy3tE3gTK
KQGnnSMdq0NVXPPF0cCYpFjTAwWku5tVeQ6ZFPIPV2A1mxHYSvxUX9SkuUsOAMKQOTqcmzYI6PXj
vLA9YNM6Ie86R4BayPNEdvQv0ZapZIG3mAvaBgDnpiKuxgfRJYk7gbjcSGFvesEKLfFhqUL+QHrn
dz32BeZre2pTrKJXBDsuJHP6YpIIWpbfGulHWM3nInV3NyRRjIhNjJ5/vDG4Vt40aXqLltVfbyUn
MXY6npRpO3KEt4l0+v+Z1ftLtYgMf2DVKNR4KC7TZBBS0ujF3gxH9ZZp/Vs+5omlfcESwzdyipMI
iV4qNzgzZ9j+pfbUQkYoXCCSNcHal5gw0+Y5naK3z4g6K9Jc29eFLSTysciNM/aFUPUkrDpzfCtW
b96PnOu49wPYecmiZ1nVVCRtfWEaHnwtCz38i7hZ9EBbzysoayWoqq2Y7PZLQI3l3K4nOdycJ/S8
oXHXmgPzlW9jAKuhUvKpZckcUlBAwkWn+Ia+4AfFBQkgvE81qSAyzuLW7eKHIJ2UqNAVAnPpR08w
/q89MQRtTpHPCDKZbVA6HqpQoZC+D/Wob5tFweSI5lAucEE1vsi2Twgz88GZ/Vq3fWs8aq3BPcb1
Mam32A6e4H9FhX6qFYnUKhQbguzAP+BYIGjM2yPFweVljO8akBkHKHNUM83c8Bh7UeYpsysqFqUA
EbiQfVdB+VMaCPTmNVbPKMf2mzvvKGktMFyNYYqY+xvkMBjHbvbgfCnxTytyLuI7ZiDmrxZncZNT
nbRzG/zw/YDfQRUiu9msy++sZfo8OO01FVAUPB9R2al+HNS81xVCoe0F5Iu8JwnQ2CFM88lFnuGc
pZ3nKTbh3GcULx0SwXGDuI48xczEeH2MLSNvJ5j7Vz6zXhY+udNeRPF3whImKOK+daNxr4TyhGUw
yE+U8bP6UAbC1kt9i7esJT7THxW4VpuuJ4Pqa54zWtohGj5ja2AwK7SnDLs92wZKzxt6ivL3nxye
ubwp6QajZ0fiEhLBFdeAgLhMOQ9ASR+Gc5REa/bcC15M8Vn/sXgSM/TCuDik4x75GzPcVwwlOQs2
NzEtzKMQcQz6fTfUTOoNCepPHQbXCuC2MGHrd+SAWWzzm0Tcg2rSqJcR+RGNg2npjiolu7cFXY/3
U8+3pEFIY8HH3jjMeiuqKSKUGFwKI7c6jSKnEu1lzaHbuT0sGzbchtrn9lgNaK7lvrnktgI4/ER6
o4vL2hNaZXOSP38ze1VNXbqffKbgzliWLKW0nX+ysL4ciMkjLsQSvKYj4t5Q1FDuhJMp9InK93q8
cAbPPtbl6VzoMX/EXmiK+faxWSdWNCIcBYwONPL0o2ZD4G6BXWsVvIkQCDduQv5oay7/ZWVAlL8X
JPOH51nvjKD6Lxbx8kbvlKLQUE1ys7HCQZN0pw32NlubIQEq0EWI/7pIJY6PVC53YZtbxPMV24QV
HOSLak+HaSGaa2PAnRwNfLFZcY72G33pE8MWeeoWLye10ype6msUw7MzuHHUPisMGlwnzyU4BzbU
RpR++P1SUOWB2AhkIyouvFFm+sJb9pC2U+LrpcK55C36MuoPQ1BfGt4nqYH5oBtMo/hhCEsOS6IM
vfhLHUAfbMqqYd62FruvUFNIOiw1/TGTLQ5r8SSuXtFvvOm2vQ/ofZsas/Ko8FTXP5TDk3ABQbBq
tqSusNP84SMPC6oFsdN/qCWVbF0AdUJm0phdqJA85bPchzaK+qyqWmI34d77cl9HZSDADTslKANg
r23hI6IkEW6lWyK51BO4B5tqCDZMHTkCAUozbCl2UoigBazo1LJts+OUypgPdoxyCnR9WS1S3EmV
znjTLaTH3v3SF5Zwl/11EGkgGHJ6Iki7Y/ccPkwRy3/2p/rO1m2+HYNJ28RTA+V/h4ZuIK7WYpm3
IzstTC2YI7DaBKs3YEPfpR2ZrwECXtf50ChevY1X8i9fX0fdEGYbc4TpGtNKi9TDivhux5hXLbAH
Cir6otpigeL8o+iO6Jbifo//TOj2nh7pRcxHGjkkIzlX7ASOpGxiNuLNR+dTxZzjXO2vvVUN5p7t
ZWWliKODLUY5yBfvCEEhzlUYw1nxZmKCFMksEoSEYbJYJg4I3ydZPCgkjTBuqAm1UHLI8eiV2yTt
9aEBW0GLR4RClxVqCf6XWu3wgymbM692alCSHL05v1+HTsJE1R3RAlrupRQqkOr/w+Km7F8zBWsy
zafLKVk42hTcICpoi6mLfdWvPHI7ioljuVcpWLeOIO7Eb+ZmF/3s4yL8AvOMJKuNpCoqKlyVG/dM
AAdbqmG0RPQ+12vSfxOYn8zSyE5eHP/I2ni09TA7loAOfOU9ElPfnUMFpryMx2IlUwY+TzSDq/kw
OXizNHvfL/s1wVcpnp7XhpBbDBhGW2BfYDHE676OC8FdBZ4jI7iRKMozyUfcNxcX7p8HgY2VZIM+
wN8Owg/FSqC0OyM9RZwNr+M6WlqE7hs5AzruJ3Acd3ze78MKu5qHoE1Sao6iZRGy9A6ixwuE1SxF
qg89AAp0J6elsLubdjyJd36J36SrQIzPcJ8W+ORyGnTvq+0hNl8uIDdWzZ92v1NCqz79f/DROSy2
2FjBYLjm1SzyOLpZmLD8M4W3XRkDYRFus0FHKr8xEoXavfQtitsBcXrFXIB9ALx6xbUoLU1CU672
bXTejZLRvVWVGHiLvPoDBFNhyhhzm6GrBEkIZ4HqLVXdR61oqmpEFTVjDkNviaAHBMwFLCh3y2dT
TMT+/egnJs6xrR4uE5CCx5oTp/PTw45qtOoiEfZPRprnRb+3K9sr6JxOoTHh0sYF9WJS3EArvWg2
AIAmBA27LG+N97jMCjlidPgS+seWt6yekcT9O7avX36Kaf+cYDVLHaF+9AdRGX9Y4ylNzyNCVx63
b4t3U+Nf+Lk2u6Ifj5tex/X/SLM4+oo/QFWa5QdSpDm7Nj51HqLGxiCMg6XkzgVx7axvJowZcAMJ
CZvq9991OucFNsCltHLQPpYAq11x6510cJbDCVqaWCV4aTbf0403T8RZ4butlCEiQo7FRKCMCmUH
b6MGMyGzGpdYBuoyD0AVOSbAkZe39TYon+m3OtAxxl5en16dk1YjjjvT+MjAoU72ClEff+DS/hlb
GdG+GnmrsDZmgvR99wgfMdAlv6lo8lxBUyMj7Ey6SYQIpnNDYFNI67+t2xMJYIqOaCrN6Ty1aRgH
4Zvtz+6rKbWNKH/C3BttWh0l3lNqmt+WLzmYJOA1dMRRqbmqP1vl8vp8/qbkDjFHP2bC7k+yF5xn
HwWy8f4iaeb4cU5KLPJAMaV9fxVVwbDj2OxgcdtcCk0A5iB+4aABeEdKqGWWvGCFP2yIBLVxsjea
TUDJP6Ffr8ycL2IZmdrhkZPQLM16PLDVAg5XlkWRLSqwO+/oVe+aksRswno34VeZaeHplXCLn8FT
3glJNHw4Ow5B6pkAEHorGVAaPX4VPBacbO3JlkqpzY2ZX3t/sMX+vvDWIzWFPGDrsm8Pjxn/GWuj
lMFiT2Wtag9F9ey5uq88RfQfQy0q4hOVK4CwsuqslRmv6SCarAWs3CMfz6dgiwvGiaoFKNV8KYtl
XGJB5NX86esJ5Kz913zkYPqSa8hpyoPs3Sql5xMSfaLfXh6OPJdvtf2h9UVfrjJrycmKtVmDplhy
ObuZsZpncPQrGu6l1Pq1k9o+A6WHzRdMLdTN4piX5hlT1g3s3izb2DVZUQUzSp0QnAj+tkcDZp+8
TI7BYPppLNhvrGj3GPIWdEb9/g9Iu2OwYbJAXYdNjFdaAVvoramvliNu8+jIcLSn/xujEOyeT1I9
CQ8Laxtg09rW9kj2094UGtRoZBZB4Ke1bf+Dfl4RSPdb6PxkMgUAqRHZe6UAcMkoxqdAayiEgKtW
klPvSebeYmbcmm7hir7dRkf0iE1YDDpmKPAvoQfHHLUGxhNGBfhnqy8wD1TwKsxPxZMs61dySIxQ
s2gkOrZF+qAfOyx73W5o/nO7gJKpGOxnDW49DR6alRbjk56PZcwEoCNtAk7zRAX4vTb+rkP8JtiH
UsgNGYUopzwqdPDZ+e73UaiuYejBDBgoZSapLuD353XVqIOjPVKvJ+7D/pNyAjAtSYoyU+6/SkYv
xFqO/AfeaxvEsdx8YYJjl0T3Zkiy1ZtLgNeCKale8QfZ9HPQ6x79yLaGKKhXH1hysoxNz9pBrUep
ElGPCc1UJBz3mwwvqU5fMzPDujo2Y6K0VACUIrEghMisZgGEsbfIBUHL7PVc4548lb5Qh1fP1mcA
c8EJ4JiOpQP/B46K61j5N8VCwGWZ/TC/iSpoJr2J5VblzJI4pCY3D7nEjCGO0fAufHnadAjL6zXN
mJT2RIb1YsriscDUwNGZTzw6ggaXOXdiryvWXfIbFu/agoZjbUppIjzWtYHh+PrYJWzVJkm69aeA
Zm4DygtmYXXPADY4tYIzvur84J2hzi1584Ltx2NPnDdTLyRX9E13CREZWJeRZ1ichHC4eCP04+Zv
r0cDiYdBx1mUh1DAYLWwREwLHlQStdJuy8kUcsp7YX26MnUy3HbbYghUdNbKFts2lZ6bFgdjehOx
Q5Zt2HAGrR1qCIgxFob3JhPP/rMaYzpdTwylGWV1fpqtlqUTsUCpC5c890AzY7MWerRuzERbnGnn
aIp1qBdNjAmAWEzRiIsGoxUyd5m22VoLC+z2d+qyjh6yHKJkQ1TXopSDw7lwWBXzMIZhFmz1AAh4
OBjudgDgXMVe9zDxrNwRs1VqrZ3ZYvj7K9lS0ZtSo5OPZUNJlWZPBM+MuSvXCmsKrMdfhOKnAQs2
FS7FdyHqKmWlb96/ddoxboX7hXHp0W0AX1OBae60ALK4s9socjLUGkRAHRIukxcDc/FWBhvPhONu
MdjSubVXp1gVjP+jgcGmYN2xdEg8Uk/R6MIUIwg2h8b9Ql9cf6IxLMzlQMasHFkU8p+FTeqlOPXi
4mgqGYfT3RS4520IcdxoDWD9J96H8hZgJECCVLdv40XZ3Z2fYUv03q39dxlixcFeRJZ92el+gC1s
fnXm4jp8j2wOHMbN3WeAy+HKxYt28V5mQfjYGtlAkHuG/YcqhGN/6/EHlpqo2hy2/Bt3CtTPm6de
uMN2DWjC0i80bXnwx9jj/+3/d4g1TmxE9EMWY0Rr/TVavtQqVehvKHxm47JsNKQCNK2AGWsPr6KB
CGb2/h5z5XZwyEmENl0GqXvZhfXVAQnDhxF9mMmUZeJCfYdZ1etZ84DIbjsat3rYhKilmYK+tDEY
svMPBucP/GUt8j0HlRZSJEPk/wVK7OlI4fq++BPKB+GYqMNTzEprBqYxAiXWjQYoeBVpFywIVhQG
YeokIthNlRbeGM35cyrY76jBVgEizoP2FIdUtP5OYFdGIPwV4pKDzH2jV5Iy9NERclMLZCgOTf+I
8h5CcPNano9l9MOKsAry0Xp5ckOPnGBH3XF3gDsiEeaD7Cb4B+HaKzLISJvrLk88FGUE91iEkFF6
YZDrNvDL4ETvtIsVE2ZIlScmaKPzBgBhfXsQ2WloH82eB4vNHUCKbPgNohVbVd9Zg15Xd10e9XYr
84v7h7yR0JPKavOtuBLpdTW07PFuLD0wTI99Yfs0U7XkIsZcgNCMcv75daIyBlRvmapqgNpbAW3u
3LUuDFV7IK7Aib3E9/f4wZqSHWXGf5itfqcOIAjd+Hl2NS0WU/TAh7HYhbPKZwV9VSF+0i1eEGLN
15rNZMeP3vbGUujQeLMVSHreSWke18DLNBWkkChl2cnBcsP7RCp5duSMkS677HNrErdxjN2C2PkC
OZF66dTAA9tmRhX6GYFgxohzVKK7QgTyMZNCgiruqRlP/7aeuOokLFHdfL8UvO4nEFB7vqobSGqR
gQu44cUwqRovCuewJY+ngX6HRRfHIAB0Uj1moJXWLUeCJQTSYzGxv+ereZKZ4DHnNbkyCfI56meD
OSoBFRKd0ycqXAIjyDvQfTjBqLp0+hvH8UZL35ccuJVZ7svlUCOso7D48R0UHO+B9rUE9L4CcPDR
40DVfvUdI09mdLGpbufJ1IcH5ChKP6/UOPgALbAJBpsNncubFxC+ERsNZxq/iDIaScEpVMVt15mJ
iWG5OKLBsILsN8OZ/htojXt+sJKO6TMH0jzAQ7gYvzsG95u+fyIukt+uX9DHPe01FPPEA2Gy0SYv
QmwWuido7Um0PrbbAjWXPfglsFsgi+68eW06Fk/jg4xgs9YkodTE41tCtoEGrZ6DDOtHGwiyfXAm
4wKwbiAGzbcPky7Cj8PAsxf7XppjchpM9Zv/4UMyqmkF/F1uvngfmtkigrWHtAlO8FO+pVyN+39P
pTFZW62b+fBidk4KhlWLSJR7UakpxQLQYNY3GQ0RN13pkeLH1QwWQbjew71wwCIzt1GmJc8L/ja3
HRy5DKgeRbN2NvuvJcx8dxx06luQR/N5K1fXRyct9+BNTnVM1h68fwr3gqp/xO9jZ/qD+eu441W7
MATf8RRiI6Fs/Q2+nsdmImn/F+GutQZtDJiM72DU496EC+rx7kvRUdSJYTyHbrCLcjgrL9pZT8ro
g4DlOJVUlbx9saSigtFflE5fVttkhpr7idMkKR1V3YshB1M7Tq+2vpytdjeXLtmYt+zUjsv1B7hT
H8rNHKupQlDZTF6yraR7LHQljIX63fLvwW83jJHagKS0RKiif+h5Kc6HXKPJ6/LoaYIQmuRKkkFI
oM7oZwPhrXi52mUTzT0eRJN8kh53pIBgQ/htglwUSVRsFWNnptJKf9Ot45a62Yrq8+6f/91fUC9l
OUTY5HbjEZcq1zsk02i7I39lpFOIX65Dt8oawqHTJFtqBvErEW3GEj5vIKy3Tjw9KxejapUjhmbw
dkp8M7/wOpvm3Yn6S59iTLIL/lRJgI4cNtuo+j+Jm62FMLmg7/CnIqy/M21gS3JneHCEcsAyw+fN
fCfhjS8+HLykCwckHPL8EE+cIr2HJAtenGBgJRNBK/syOCqcl2+AXpXmSQYnmlyGGQL+dNPbYvNy
Y58BNPbFQ9x0xyHgXPgX0qNS9PPIObBqONLxxcPfW7WRH4ThfzBHfvq82woRBkwHYBRs+ALzRsLX
MpdkIFLzZDo3L4BELahd6EDPc3flijon4+HWk2nefBOphJ7Bjwv6SPU1GwYHb2bPEv0z5NOQqmsc
AMxaO3nmdGtrcETf5cgb9thQgP+x1b5zkAJ0mKQIo7BVC6sx8z3ofhUQ6PeZZ/6SJAG7u9yK4buR
LWAQcI7GJFPYuv+AhIrS+0L3dffK0jNWIWpI/UWam4dx0NHFTUMYCB3vzqsCQT3ty5YVEY68xPRq
10pHljDUVN9e3EH/DVMqAesLHJrejxArKadDYlqHPCzf2zaT9INqfSPz0oLuzUYvX2GuQy4IlZGb
Ne5LIohOrbXEbMGvhsuKemN5u5WcER6nboM72JBpYyaikEDyTC4DRAvtjoaRqUxIvVbX79VQfe6k
WBbZAG0R5nJZluEqxmoE89tt+r2u6/N4Ldeu7Wl4fo5PWHft8EqeiL7R9wlpQWa+K3/O+Bukf+UR
wspTSpv4+LZ82Pqu3xI/eMC/rBkHTEAPE+LuRmFi+EbNwcmNSYOzATvrjr0k95Sr6Lg/5slKOprb
KMTpqEg54yrCWU2pASggZyQD+5YAz2odqKlUA3WiJCFyAyozpBcJ60Z9E8nvXxRygTS1D6s4JkPB
n9a/S8z+1RcPZpjNk7lzz3mv/2BrEZuEVwS2jUU0ktv7VfLvAqaD41xY0meQDJc/YCg5k85yyU4U
nD8GtN3P8WL/cQxZRwAcFdD0WwAyo7pLy36tjuQ627p2OniTA5NZ3lEYP/an/tszkMk8bD/RBd7h
EZIWeZGwqmSHlI+tlaZXGRt4syQTXfrpM/elGjjm1tl8uleTiI7CHlOIzkVpsL6fHYkMRtvtNIVA
gJeDWIqShfcDWYPnvW1F96YPommPvAwedtQM34BsiSsLRfmz2ELFSe8ulGO+p3qJUxtYsgPTLyW0
9zz16gBIjURUKC9uuih7rJdX4csspyQxgcY9gy2lbWYFjjhdrzbqs0ut7kvFEYutA1EBOJzciyRX
jNqFwqfPSTVY10Vbdf5BXa5nvW9wTmdbmSruoL0oCif31ta2RJZyRwFmL9D2V6IpaK1QJDkVy7fx
60xej6fVQIRe/HykI2MNw+NrXLn8tPbE2l6QsXg64ti0DebCThZ/vdY4ZwMY+PpQGP1iklRmrtYZ
BtTQmXUe3froijcRwmW0KFMwqIY1oppJvkdIpfuJYMAa/w/7Op7qz8g7D9q5D2LlB/8NM2xRJ9BM
qC0RXm89AkCbESvHCHLaHTufe7ji+IgIlGwRMsbr6evBmeII5ZkEXwrT1Lwb4x5/Ysj7Wy5AS8H+
dzr3EDSoAEmC/4vDc66SeXN8rrFZ8bYL50Kl9n25ikAX0AqWvxWSm+e85sYshU0qvFPeiX1yw9MI
BCVrH2j6O/RE4FEubJlScn1Sv0YxL5Jv+tajBdlmGkXFF1GvbSi3dx++o07dmRnov1reY+DnTQjo
eIaHMCwtO9PjY6/8/6SCt6+UUBoiEQsU+WVs+ehLi4Te7jqcNdoER1wTWQ6wY5gtqYp6KN3M6/xV
pg+utGYDoXE1WcjqTSeOyUPur2eXcvHXMqF8S+4IBW/UsAPD6QLkkeTEInu/iWo00+HC38JxGiBX
TQDiXJMA9Lv5t+M5W8n0YQAnS80NRmUdbiwVaLYkWvxdW3N4fD//MqMb4jrzUZvfJQWTjTxd0K2r
AahtikwAv8mQCYqUY4V9aUOgJkZiazk6a4E6dPyHKPDbx8T4XQIwpCQjdyQ2cVe0ArSMXpv7LslN
TsymzWZZnktVO/pmj45H427l6ckOveQF4BZLPtlg7UjUhTeW+fDC0z6l9EjqXJQ1xdlk9cHQrvYd
3epJFIii67vTd8TPbEZlPL3YJNkRHtUsa3JQaByl+fXpt8xNAfU9/Ws2SUYduOaFpK/mLOV1mYWq
gDEBBf4VBaxzOAH3VVGunMrg9iYVOXNK4waU4WNAOQ7zKugfQG9McvlW1AUBa4AXfitzkQPJ4Vwg
HLV0K8+1CaIWQ4hB2nQS9Fmwjhro2V9xddOtiQQJihFCyfwfYNg2p48tnfojrW+iXsoR8YdxKGMs
IKO7CnheCOchoh2LI20FyKhOMDTlrzL7zqT1h8V7zIiJArBIR+jx67U4MuRmFyaakejC+vuOVIKB
ZQUaqN+fDsa0EQS3Vp+KaYy9WABNpwd1wzYS55dkn7Ojwtl/3Lg3DYuCO0w/AwdPCcHzDy5PRyra
xXqNcafJ+D6jDKxxbMoNuwo3oSGV61VAAQ7ipieI2LlsJAntTVIQjCKIrDK7cGt60CY+WO9k5y50
vtn6Gkelw4svZYEifANVvx8hjbFQD7mtvjiHSrTyeD5GVcNPR3FeEk7lm3CnSSCfqvrNW804voOJ
6NKFjhbydTRSVKBlLyRm4P4EiWLYVFgoe5Y/hFLziJfaTY4alIuj7pFi3rf51JLRpoxiH89NNwsv
PdFbn63qIRYEAQg9jSy6vnVeJIBF+c1W7X4ahxi+NqaDTpcGV5eDppnk62IhxCUrCuYpeF1mT2GV
i9phKpFTEfjVOaxbvkGBNnUHT7iBL49NExUce0lfS33+1iVOBzmnTEQzb5C2SdNZI2lQPPFflOOz
KE+MfqysxUvOxau5URihJUNftS0Nsq91YN1Uw2dmwdVpFNGYCuUYjjcMwRKYfqRwgnLZxQDPE+JY
2ExVHO11w5UU6Qi7Iqrf6bLgJhH4nVHLkqljV0O8R4DlAeJu6Gplbc0L7cqK4B5zg84vCQd9irPJ
FBXXuH0sJi9auA0S5jKOBN35GD6x9PfLdqRxJmWrm+mqciAO/sNxHX04pQN0ucnUE//nrCxGrawH
Wr4VmYU220LWqT6QMcvqHgIpcIpdw+ZVcKu8Dsb5QEqBAigdVy4BIQFQWFbBR8Bkxlgwc6eDcE6P
sIoAofGy7j8+F9RSCOCJAjWIZNQf8yomTV5v0YH3STHTNHM4viDlZVMYjaLsGz4hjED4hLg7j9iu
0MyPOSx9T8u/IGQ4vGpEiA+GZ8Ltany4meCGJgfJyeUIxXV/hceSD4V1pcNo6pNzuDL7BlITcjNu
pIjf+YN2eag9AX1+L0v3BwHfGExGwg7kwCkCL3uOI7fNxTKfj8KinovNO37zhIZGwYtm9RRiHc2k
C2uKd4/rASSQOY3BIctUYO96QInU+TyLvN2eofqJSjMtzUY/IBsnR8HLdSvWtULJ20wtB//V6457
U+kKll4BqFshYTB2RX3FKqNtygwp6+NlxJZNLQsjcbeIjQwieQQUUoZ0SuV+/6n1pAsbk7gwO1Vk
yr36FNuFzDCqgzpUIjz39nXINCzSz2l7oZ231zzBE5nhxxhZi5DSdkweSR4MHl/bHOx6yLL342HR
9tCk4xamXC1C67a8+FyQnu4v6Zirx62sN8h8PbPW4L2BHnfx8IOR6FuaRqt44r8oX+d9GHGHmGpT
16sMVEe1O8MMRY2YRpXJvaJTiyA9mxRR5qeKOHPUvSknk437SRRXEBbCeBJ27lABpJSUT7EzCNx3
Y2xAOjErBa2ydK0oxJn28cezrbpiMxguMu6vtjXDZZEhGRSLANzeeSBzcDI5bKZp42KoYQ3ikdS7
qhMqoWmuNgm4xo0GbkSGh0YYUm1vy84QHspiQ6WgXEdHi2lfUct7XbIjPTdB64VJJKdZs9fjC78t
3C6RHy3BkxhRjqmlAgIYhzkK1zj0Z/YfI07Da0IIjZVIaKu4e/wntoGh0QuL0mT9UlCqtFZ84Rwx
a+MjtiGOgAZmWCnPLQzlIzxR7FcoaDPw93QEakFi2+aZc1uWWzPREymUsVKtDr+LUXSGqxz2clbd
x2Fi75YuN3lecxWyadVEEbj7TCN11FDGth4cZYuPp2xukS6UEktxxYdWjXT9yQj3Lp4fYRFE8MaY
eLiJV77YTxc2oz0KzM8HwltwExe9bI4IMOfsCtcC3jroltuJBjE1nZwCfsmXhc8OZOQaZxkyee+N
jc2mjrud+VZhHlrqCzflWoAu51/Kb44TjIq6WCpJKcVRV/2EmKy9Q+ooTWGTwY2EcEG81BQluBqS
qFgsm4VWhfufA97toO46aQkRffbO9SkcX5woBFtA2S2/XryqfooledPwnD2hGT8+gH/xpYS/fTYm
q3uSSfkgtkV1JPCSsnkw82CLCY+izYUQRflCgUGZ/+YZKqcIlOvcN6pQVVbK+uf+SgxLFH54cTys
Mq4IuPhq2ycYJQTR9RvydfXXDijyHbgX8GDPH6A4tumyS2ps6sxujz6jhpX9bZ7+PNeZBs733Bjs
dEr5RY/FS0BX3I7H6G+RPRz8IAR3MtRuxf3jm4TrWg9vVSxs7lfeLPFrvqLRlqcr1o+THurIAVxt
qioYv/Cgc25p/a90MjPF7E7kEP37O8fp2IwZRKSKSUHWr1Aa7axRBZEjnimTVFybENfBvajGCWtJ
mDe44yiogjXRTH/e66PP5H/qgBI4xT78I8YQnogZVfSwRiJwICR0GS3qpbX4PkKFwzRt8rZZlun9
P+GQ1idasPivkHLX8/Kt7X9yG3VNaMtZAkhyOvBwyJDKmhasYOprKnxnzlfe8e679FrytOw1W+Ze
+CNELkJ2ShDR1VRHj9Ks1B52zuP09+wrpXDf2hO/9W7fjS6WoeEj1XdAOzvecMUMbPAuXPJmuL30
FWPJ8XHQ8WnOma1PpqzYyWT+R9JecXcCebBfXOf8NGFd2l2FmbRTxCRcTXNBdUahsuNDnZnXIXpf
LQcqQxg0CtaGjGd0JsHl4wMklo2tHAPsD4MlghHbbxeaQ1ewDU8qYpXJSl0mX32pm7YK5b5xdZTr
er/TDveet7M2x94/Am2dN0S+gQcYv7l5oSoPDCIjkrCnpfepJZqDdHAO2aqJQZdziWcs5ZAnqZ/O
vuvfbNY6XIL6JgEWDJ6HU1h9ddMtEWQM+5dCnD0VLcqBSNiaUdWBHFfNQz53qDrZIIJi0cS/dlcR
dqD7ZSEwLuLMgPcF/TQ2Cpufy8SHJsEiTYd7odbrdU0O8Lgrx4nrFzmhY+QzsadmyimqPJGWlKVq
bL3yxcdYcOGv23NlBrNfNeuofmC+WahKvItuEGU/ftU0LDleLr68zY2/OYLal7bog6X5fO6C6oN+
NEk138bT+NL4BH541NF9K0/gksbmz8ydleSLA7M6cP4z4A/IS6Sk0MBPzs+A7U9rkNx47cWXswAU
orkKh1mnnzAG2BF6k23gBep57LGNmvYbci5QgMURe8ACLPysfyFUeATnNve23FqlZLhoGObDU19M
5rGg7ccq/zmAVAcxK90p5pfFIEWc8DJPY45bl5wTyB7Ky6nSz8JhNtSUzqxBam+N93EW97XUPa5A
Dp+P33CjjbfxUQJVDXV2ZgrpfmqJ4ahZTsMh5sqEu3nWv+EwHB5K7Kn/IQjG8vT2VzeH1+VG7wE/
VzL9+RaIYHqJ7ZPu4bZMwEBZsw18a++ieIMINp0zTT55kFnkc6zlFbpnUPMgwKmG6U5IHUGffHxZ
KtPtmAGCyBCAtY6WzQ7rJvFfupuz5Tp1szzX46/wTP//iEZ3ZQr5yje+bPfbPCxwie2N675+vVzX
nPd8f0Nta+A3UXdaZj07jbfGXvgC5svS72NWk3mrqRF7+PAKK/0YAPktnKTlqcW4iXWlPFgAdcpz
hVBAW1Lr6G+8LnWoBjjItl6E+Ia+Hv8vJSqp4I9PG/5MsFSuWjs69IUbM8x7zE8hARsLK7dYU4YY
fvGiuWvo525cbrAogSUPKomcu/35ryM216gThP+Z9w9DnxRlsX1TaZKFXYctiiUzEeO0ht3nGSUY
GFeI4+XbtJ0pO2MCtA6ZskCx8MKkqvkvIKrYe2IBT/DyV0Dx9EgJAUN6+DQRHlEQ7h4SJAedekEE
T58ds3PAaN/aAzhXIO74kn2rYOe7hJ+iulS5u49LB0RNSlNf+e6mkQpsMr3t9ggfGd7Wjf3tXQyq
vj/kcbgdIj5PEbyjq6QgF49ZOVht+jeLBBEx9YjMBEibpbinxI8KPujxskEKmrEr9BO69IymLgUm
wuIO2Ozer5LNyshK+8m7Ct/IrefLeytn2jiMd/6oswIysCYhHPL6/OkoJTFQMR7mkSCPhY/Kj412
Li9XZboceAHhH8GsslWXXp/KHNjXcXhzQLnj+eOy27J82W89GNiGpv8NoWiddAcxB3zolm1oL1wW
9ogaqdtC5JDqUqrpTnVTBsTxHiSIoeKJ+5anSHl95cb6jf+j6Q9MQ0wCKXooYDXDkD4hwBcABW11
UgGpznF2rSLZ/q/7SqkahyvKi1zvCIHxx8X5Ky+yZiqfREPy/c0rWOgJyjuOrkd7/4VZUzZmi0w1
nflnU/zyYFxn4u1eHqlwoJi3rwJSp/ihUizPEM8efGPvouSQKXXMtHIiwIdYNkmfoGIgqd/Xe6O/
a6isPTCGu3EzIXsyiMKDTCWthH7ECoc5rRALoZXWPDHduF6OeXbkj6xl79rKHap/3oJ6Z/bOU938
/T399bEHtq8rP7VyLiyJ6HyvCnSY2X6FwD2/E9HUqSdjPpyvlI7svBZk3X80VPSm4O2R2vvpWMZX
wTzRj34sGRN/0fpiBZuZS8Mm5ErzKMku9jPpJ5/lu/YX8X/a0UhZhDFQQ0eG33EeyUOCgac8hTVj
Vd+HvsEybfNQuAMj51PMZVU5Q7KU9ez925Y+lhKR7tha4EseGZldunQ22nsmOu5ujxfwp8oQ1j8d
9S2nrDVDEmHvhZxqHpqEbrMtYOv398ffbFKiZPAvrCK4/B10SfkqAavEh2mOfPG7f6Qq9l6rm818
DS4UGwpST5VFX1k4/xbK89OcB3caa6ZlDTGNUVpegEpdZTOpMU1j87fYf59iUlhQQESatnueWB9W
80xeFX1Ws0rnDjlzrez7zd8mwx99k2GuOQ/YTuNddmeK+2MPpV1/ARcsqFw8A8YQaXAABsT9+d93
ZU8kN8k6cJ1+bIvoGwsOEPcqnExUrvoy3sgWA4j+i+vnnTqVC5gNzsDNhknbZGyWKf7L6pwdbB+z
Bw9y0WwH0PxVqvDfzojgCtOS4qJf89qwyoO7nqkqv2EMyD82gbkp7enblwVde5r8TKrcuYQ411NE
0aa89Pcq3MABAQ3pj5l95gV2tnMLJDkQylfpYBzhBpUnTsNs7CyBjFmAD9QgTl6i2NBgP5C/S8Wo
1u3dK6J7x9Gopl1dlngGAgQhesYXB6WzAQvpzGbwKMzicJJuNCo8tobWfqqRHFVVZhXmEYNNs3BX
XDk+lu5FiMH6uv0/hz/Wg0bmpy3sPxNTICk+sfyPKmOB5VUCR3npSW/sTwq2I8X9Q1Y+yRo8thdy
V+Vmu8m66XyVfTYwiouOO5zu++/1RdDVyySOIe2a3Z6N94Si0Ho0ANGv178zaEC1Tl+p9HiykO58
j/6ru9YwAL3D4yPolLo4DCDHFY/si6EDRNbc6UuxjrpUYoiEAj6Cx2kNWe/0gm30Tmk4AZvOVu04
RQCCueniKdyO9uignvNo10EQRjwclVW9igqgdIeN9zf4og+ByAqRgQr3xhUNnNdnMHdNK4Hbcmxr
Yl+yCDFUCAyndC9b85TiEq/SMRI3M4UaYP6TJvA/UFDF3ssUTJT707iKUXWSVruAbanr1ibZ3wgr
klt4Ewz1IA8jW6mHg2fag3XJq9E40X8Q9RVK5kisd6jhywUIxlBTffUhs2fTkTCrjVv4qBjwmZeQ
j9vXv2t6peIXn4EeuH1jJuR72rkVXChLZJnxY6gfuedtZNODXHkJDtewX0jTEfSEfWm+LJywSn4J
qLe5D57O5cIB0vtEwoYu+A81Ej5o3QPQ85gkOIGy3IgC7vujhjzflxVF63+vjWYvNG74UXW11W+6
NMKImPB+mbJfr1Xv5JJvbc2v/HhGw8Ypsud32JyDhyUHbjf2c8yXyr282l2hETI1hHpGUu07kYAA
EYDQNb5Hwzbh0hUQYPcURxrEs/tabeLmBeUljo4DNH5RO2ljr2JOQwjGkyZrTA0tDMiP43nflXsW
aM/GLmJWyFsdpefYQXtsnWPEBdwd/OGHE0TpWS0/Hh0J+75+hrecYfWrhFH4786eJJtHF8GrhEmW
4PcDymrfGydhnR/o9rFPqkcClTHzdBXUP4/rGCILDsqrIFsI0W3ptKIDqSUACbiOOb0fBweNfnVQ
3pjUH6+VNUvTxntldmSDCNPRqhdMY7EUG6UAoCX5cieh0HhKmavjX/ksfnZvKWp9h9LGB78m+3vk
Gw5ctJN8SmlMyBvK1SUc5sqvb+PslLKnTeX2ExbjlTDkH8NzUmoFcbGI2EGoVGHoGL/zx3DBF/mE
bY39TfcGqgfzPn1sBa1bambVH/HgxvTGHFsCXTQUyHi4rYfSRjm6d9f9Td6xNKQ66DuvKpVLek3E
xvBU9MO5QBbGF4EuNSnYMt47yGAUZOlN7h0Yb0Cv8tKnqZXPSgm3ntro22Ou2nQpdqrDUvJZgPle
0Ridf5MhRKFiHvQ6P93VuR7EciYWc5n9KeCLF3mWWkCmzpDadhlV2hDAsWPhLK8mtpIm50vDwWqd
1lpkd6qCDw6pDBNUX0zyveXEgW/P9NMTJ10RdG51NG1MQYQug72coJd0IIwkAZCcPDy1aSUgq1uo
/SpFKPHHB/NFY1KhnQPw9Uw2IezKBPbEMWzNfj5ak9nxWf83Bba19PdyuA2d7mcEYxyR7N3pSaF1
sWwMmo/RfDP205jQXHSVz6Es6BcwzYlkcFmJHWdXDUaDVyJ84PCq3jbJZ6IIh1oVjkwAq+CiEKLi
YdbpBUrlI408gqS8fAkrasvibkQ9EtWm3/QkrWiPQtUYNZeTJqopYDH+bRw9nZLPgIhHyMwW0GTp
CzVA+nOcfWzcekQpq6EZ6PIKgc9FU/99IyGxZ/42M16XxNFh2hMOTc59E0mmOQLU9gZluZPaIaOh
9e55bkS6oJ2ltklatsJkouKVeeYynbo2Za2+gpCQj7APxL8x6XHaLFkeDIxwwf7PvjRcGwCvCqIn
EAqJBOVZeBGeKA7WX5Iy4FU0/NPuWm6Gmlz/ljKrU3gZYvb7S98fly0YeTbHE1lZ/srDACekqT/a
a8cAhVfTpzti/25m3zFUGrLyi8BSCSAbTc6WVPvKc6WfmMm44T/bqc4fHm4dHF9FGqGlE2N77qCZ
6a3ocb7JOzw3pp3TlHpj9680At+IAr7GizO4egGOBp2cH/nye8/ojIVfurz/RCw/l6vyEj1V7Crb
sGilJtavOk8v/TsQzsAOK+DDoZnV//1WTEQWyn9R033Eeuxy2ZytOTJ6+sfoHFT8GeWX5kru998C
ZfCkquo9ppM0iKntDqtO49R93U/o/7AAILlZxxjyHY+J38woJyjmkIBkY7q+JYVcfm1+YsRVHjZh
3I75N6+EJ6H+b0kIm0YooheQDCYgToMxEdD/pkj5TeDegi3apbGkwRy7PjlDYC3r9v89BNCrTu5+
1kbqmUlYxx4U5gLBcvbNv+sdu6+qGX9Ew1UyLI6tQWKnjmUTke6nXOGd5Fd82EaY+aU9nMWhj4nP
2r+j3GQo04YAD1MD32STj5JZ8PUXmbaaGjHmPxsIGQC7UBZ33Yox05fr26PCX2GTm8eNXEGlQ9oY
WaskyMZ+6ENf6TM7Lrt2xp+i14T66VQzrhtvUWrALwlBXtDxcqR29D5+OoiP+UB5zytuUjFuetni
kA22iyW9XrB3c5oc2KvfB42lOSSeMGTa1tXHjkQRFsTf2edki3iUaIp1d40L2kGRrRExvUsuJpxA
Q9lQRFt74GL5CElPG9pxBv3Jqy1smRCJMXFSRfWjjlWf0r6lKSCbs+PYVwyD8Z+WChShjGC6KHrX
mmxTnvoZ7hrSNF8x298IonjqNva3JTszXDPVDUB2nmlpB1XZL6Jh6dzpH8Kgp7LFiOs3OR1JLmZT
+KaTb2dHxYDZfTo77XgrL33znwL5aqxb5ObjCkz+KnaIT0+azY4IkPhutEWY7bVIM5Nyn2M8P/cI
rgNmsPAPIfsLGnlkeqnD5ZDZpgFq259WMhHf3i50QR5vnEUfwILL1wFQ7Qp16RUEH+xZNmBfzXh8
SRZyCGDxBktm+3Lqsjep8mUy8z2E8+3rCbCMq2VaKSLd4fFimaAl5pOTQYG5H5km09iR62N+/fhL
xB2Po8F7PtDZF85HsgeL92EbdWXO2fjBU9WAj/6JAqf/XrE5esMDeff6INwJ51FJAEUdT39mBjEl
6OlZe56d9DFZsOloIeiOEk2aMQhlPm+opso/o+KGBnWUNuVwq8Hg94fet9vqfijDMIaddNwBsZJZ
wqMVZvg0qONsccOmftEzfeRlsd15bjlhIM5y589Ghqf4LcjZb4XRz+UVbNdpciMGWAruR4Oxbo7l
XKL8a8LW54QLIiops1FQZRebDr2Sduecl+EW3957r1r/N6VRRucbIXlDE3UoKjEbM75FW8RfsWRq
0pb26A7lSDIgaY3jSZULwCAW7nfR9HiURDBG+6G/V/nfOE15Uq0BnmgaaV5n+cW+6aPHDqBKkOyw
XqiQ3S/Y+uLGLXNBs+z89IDlddho6GRrXiFC5dW2cnDt8srs9BKQi6JfUl8fYMduYYw4imrKciB5
UVrF3OYNTluu0JSq0coiW0/+Jma9ndHSFaizsRadTjiITPjZ8pIYXI+r2CPA3dfVE3RzW8llu2EV
DpVRHGuLzXeIHUsT1Go5h+V8fTScm9L06AH6x78ZS9mcg1RZEZY4VYC8yItaG1+3W24DRCIRIOvq
iVO+4ejghA+bvJFSDA/a7DnxinWzUdumBgMwW/vtECYT/enPVkLr1mg4cpS3V+7KoNZnGqlhi3EF
zkDh1KfHDoURFH0BomGgmzlIysfPibWlqnN9szSWt2kA+xejPD89oHMqESUp+eBEfrFoL/uue5hX
XUnyVr5ZLMVavYTuQ5G9pMKuDpWbiURiEcR/upoBGS79KPRghWTngqGT55QV9coSOMctR8zqdk28
DrezjBLTosqYYpO6LyzyWpqcCPqWASzqH8rW5VfQeGoytTzKCR8AdFGdIDALvB7GGLlB9L2WBMDJ
AkEj17u4yYkcTcpm9mUqT1q1A48QLs0gh2qP8+NPTNmPPeJfoP0LznQZz7Clxw/DNenZXu3+rZtg
2WK0YjFQwpMLV8Es7eLmEIVUAoqcpJxE9qQrm97n7R3ZqWSf86zugwcFny8QFjDjxuMmn+dCaZc4
ItRgyHY6Oz1TRvzAHNlWM3fjNrapC2dy1U7phqJ+NwR48PuqNWRlSdk8Ljr8RYji/4WVEA2EC3DQ
Kn0o/fg70Mdz7Vxlpr6NHPKwhE1rOLGWQZlau+5kYyet84jMhe7nKwhy+SaG0YpsD97tfamekRc1
c0BtSyMUR4g3Xds1lq6jKjK5wEhqJzwzX4wqFvI64mTX5U8ZQ563uNx8/jU05z7AUZq7VMgYOECI
Khz6axu4dlwlnd4GrL29izIe413trdsPdCeFPhaDrItKVf5JXt0if4H6hbMf2q7KB7DOfg9hvD0E
2x77phWeyAZ+QrXEPeujLMcWs4tIF0oCaIDYENQm5//ieS7MpQKcRHgxfuD8nYuVhNghlzu72ALu
vkyGXCd539RYv6e73HpwJGogT5fUf2Q4SamVwgIZ6W7dS2+yDbK9hid6gs7sLeIVyRLKFZf7hjdh
7Eoq7Ro3FRHXfAc8R+NOaC7huWmk1F48wi01N7/6UAVNRFuCz977q5lqR2yoMBGNZT1UWf71XGUl
5ILXIiCsDjEqkLyQREc0WUhCcsTu8x3pj2SrdEAlG2AHv5r/gZU4voS5SeTFbIYuMHp0qjcAZOH4
hX4VCcIMvVPv5sbpcyLjAUFuc+P4LyEts61ixl6ZJe9NqeY/nJJtlbmNwGV8FNm6etoWy8EQ0ZtG
fw0ZaXywgUvVyeYmtA5SPFF64ZaVUiRGKGkjidP2qmHyWdHkZMNrT8pHcReHmsoIVnOC5SaNr2mH
wyzEyEtpO4TilrkWST7sX03dU5KQrbTFchdTnUTBjHkJatrnbCaAVgyZVHZuc8nrq/wmBB8yt8U7
9KzN8rPtChlLBCZ1VsteHtugPGWkAmQWdpzy9l98mepZOUyWX+uMf7aNZy+Myya43rtCxE8NUair
/VbRkBH7oraiad6QwrSNRhwP/iHtZ5jhdKc3bWXF81Ldp0ymZBc8QYAhizcnOQ51Y7C+QSUUkLkK
swhcIU+VkLoMfocPCjIS13C9l0yAxbOXZAL8UlR6+UGy7/cK18j9HpPfe6wenoFNzYQidKQCiIEi
t3+TsOSkBkXjiMcCgAEP7pmKvAXWjGJUHD4CebOclABXxDBPz5LCkuNXAro5y8In6vyOhETPeJfQ
a7Kel6DNlg/AGkyOQ4huRgGVOV8tQfAIhck83XKSlWdC7dtqdiGyg0QIIc0z6w6cZJnja6mBqr3G
FRN2RNXQfdC2OJBMU9Pzxroyk0XvHdqoMubOe9+bwVnyTP2VP5y0qzXgjuNxnEG9x9tpJdQy8+uD
+GpiCpraftzD/x3J4QAPT2TA2cfaSbvnyMnD4OedoaRX/le1XVWOjF16iQX7W2R+45+0FvXDETxA
y9JOB/IfWVcEy3M9Hc63l8Mexkl2A+qcNFlUjjcsmU9OV5ksmsoOLLlXNm7NzdDDjxZJYYzVXIL5
c3um1Fv/RTbM1Vlu6QFD8F94iO4yAFvCAoc5BtWJL6kr6lqIicrc2/1t7ZI93xHY4yDm2gr6E7WF
RL6q4GjriKwQMnNyvUOAaddvAQCTwBefYvpWyGBiPhkvri/ArAVIREguuTYzYghb8cZAqBp52Dp9
Kj1kYfnRu000VoMTw7/iy7xf1n4kVmQkxqiyaXoj8f4/sTHLBJph2PVOeMYUeQrMU4jVbMwxiABR
x/wxPUnOUwy3wDVkjTMBgjAf9Ysd/kEtfarqr+R+In/SqfHQnUYReLpLO8GaarZScBWcIFpNn5Cy
n6xhd54S2g+YYXZBej1XdKJEZEoUF3kHzYzOn4Blq996SffZ7L/FgPPdp7rGz2oZqmaCWdug0nSS
tO1UVBwr38Ji4caSqlUZ0B2c6+TWVSfRyispp349F+Bufc7T48TpsSTyyQGEGlFsy3bYBOeeK5Xo
b5wQbOzeHYlIgTIhPFSnZzzJ/sO7gACMyo8kN/IXvS3JIxD0rwciIsdb4C5mTxa2cfO9Mw1Mt5xU
ZDkNHMUrcZVAAIavS+SuHB1kqp3KG2fW0y6pwFXGP6X2t+1aGEJpySG6hr+yXNV2+y3Lhg0xpAwE
oejllom1CSYFu5ctqbXJI5Ktt12RFFk9DiObPA6nURccjByrNrjShh65CspkrOfgmNANCnwhWmtm
TGH+z0uN6teKMl/lRiE2CfWNmEsfiHUFyeJAPNS+UX7sJtTiQikhh/Q/7Mr+W2g9k0qxei+cekXM
WmBMb39k63fwMNYMzbJy7MaPMcOM82d9evgKW6hjhDuKC0FfzJZzYPrQQvJgdtUvvxzB9ZZOx8jr
5HG+1tGHtZI8Cv5/2mTi0p9jFK4o0Rqs0DqURBxunmT8ZjKoC6fOuMggqcmM9nWcjUmyQSvOl9Wh
lYe7E7Kj14ggh+5lZoGiauvIPvhQWJ0Sbor8CTLAfp4nAJ6FFeiS6bVrlpKF/bG4gPUdpuGWqkCZ
XX+Zmpf9jWNi1NqvqZEUQe9SwQPeYtPEHV8ZE4y5L9P8UApNZfMOXX/t7NBWGLYqcbVNPtu3MYgC
mRKzcd63QpjD5A2H1HbGX3Al0tV0yzah/wPQzqjgLSi7r/Di6PojcpB+kTINgae5vLTF5MzXXkYg
BipI/oPp86LNtNSHPN68zMedoXv0Grd/r+uflfXVgT2D8TkPF3mzxJRtzcKW+qfJq1gs1e9+R8W/
eu3nG10hVI4xXFePJb+kCXh9OowvELGENiqM06lK/lziWdC5suJHB/tLbv4fNB/KsjCa2QT60N86
BSR2+paxbnKuZeLgWX95tGK5Q+qWBvTE4V+KLRgT+VC9t7d81XGVfVKB+Yj1SHgVLuJN5bZ3KrJA
F0JvA7NukAhZg+jtUlwxJaZBublAgkoyzclYSH5CeGc8g2bm9e8Z/Wi/NO864B8x3OTG9xo5PsD2
V+jG+cf5wawoxbp74XGP7B4xXr6xsGR4Rk2urC6PrPFxzt2i9H10cvKtdDfYXydVTLo2QkWPTnb+
rCxgzwkSMPz00DRT2sTeiP5wolw9gHskqGr6dtgv02Ux1DjilNMJQvbffjA43XUB9nZQTT8NxGJd
7RJCvdV/ekaRtJdeiFqnuNgNzqInevoNX+d3PCOjGFmhh888paoJJaNdG6QyM2IU/6owO0sTCH2j
6kSNxsWh4skrQXs0hqvDLLCbm53jCgTXlwqxeGmBiM3BCE/ZLiINy6m0s1CoaIFZWZSUjZV0a0bn
Nj7o46ipKajvR/DXCwNvoaaBiwwgndfjXAOZDtyVagNWpS3SWBZID+NWxGlnW3FIb7Oie/ydHpAH
SVpJgam7rVkAgi7Tse0FShznIeGtW5EiEx3L9Z/RUBBPzK9IlEm1g12CM/v+bBaFFInpabAkFRKf
RlbStSd0ZIjfKSJC/KZxOdvwqaiQvjlSRJEhv8/9hhxc8JDIv/oOyw/4nxaSL6J7pmbrnMhvqLOu
yy/h6xFt353WKI86jhEX40ynYm/0NBZjM8739CMJ6gm0iUJRVk4bixPImkz8L+fg3s6Lfp99Z/g9
WzZdRdHwjEAQ1ikC8na+g0SVVlXsBoGN/t2OvfR7HMXo/xCHuGXvO+7y+h7M/hjf0lJRJxt3u4pt
fdpidOB/6OCxcltINJufS211KihuzIUp+p9/ku7+rVtgw0uR8GlpOjk54zgk4wrbw6t00wc4CJAx
ii9J8LO3mHTnevvmSoQ3O2G9ZX7WBFcpuPaK5Vh4Z1gD+x84lCbDzmEik0sruSnPKhT5lf0/3XK7
gB7+QIyJ3nM5AVnyLYg2hJe6TJAYIuRDVREniazAvKoO35wukODoI+vAVRdwp5b2LH9ZFMuuafQJ
J2+2uETgvNojoC+XS3jjNafDofoJgau5y2fjR2V1OsLrDWsYMHVF6LENzP0tiqGqb7NR7jfOdZ4o
W7raiVrLcTVOT6rHgIyB5oHrA5ElFFY+LM0lb6GFIjA63fz1IBiEU8mCgntDGQ+AHGMiFhT/JAAr
69pDgkVk5Ec8whjSXdyffLH/bPnuW8mgXBUEHqk1Za9UTvhojoNZBlmVCaSuhGM0jSPXqqh3J/1H
9H2B9lMJIHbrCOjdRHBwAMr85iLWK1grZu4EZm7kW6Rqx1U6XoIAkxQjhRNJPuuLIDuyRE11En4m
JaY9sDOrQSSPiuaboOod5RKYnhvh8Gr14rQhiXaUulzoM9iZ8EG6iDIQaAj5zJpOnC4bqXjtD+p6
tt/9GjZy4bCn6mtQGsLhNyarN8SYkdDXaDHn4ah1g7l0j75RFeEzxRvDsHjEIyQORl3I7CZQ+OqQ
95C2/2qg1T8ev93jIMFaXMSw9CimyGWfhgtEzZCCI3OK6P4a6UygMqvqSn4ephK/XkrOKS4wkhbo
JmcL2wNVHqr30h6mGVqj2ZCT9AI9NsN2yfxfi5VCr85suPZ5yCQabzZqT5ZNop/DMbof4CTGEuzc
VXc0+RAlbropDJCJQd/hUXTkUfuiWh1SngG5YuUOrvsDrBk7MR9ay615ArXOQtTotflp/W25gH92
nfIzSt8QWrAl5PK+ZosJw2dSRtE5knIR4ad2nY3WkHX/8/npELKw+jfzqBp10F3wKHR34rLOf5cj
r5p0eD5HF26Fors5mnrpdjY1riZexFeg41Y5CmpHZa/V1RYEhCm/s555eidA3Qp4JzEHjFjbHyla
yZxhAC8BWp/kacwOYxI/aHMMwnsRVXhXGF116L4c8sF7KBpZ03pBD3oY5m8VaaRCD5PKQvmpa8at
RHIe3YeUROJe5E5a0QEzK70ZzSWU+81Vpf7K/qTWUV4kKmP0FVX1yj2iv+5NSAJPzBhAnVrQ72zc
RSfTrbPT5qFBvf5iuQpKkSerl8+V1H8tZjKtSJ9VDlugT4N3W1J3FMeRDZ/pH+1AUtPdMMgrs0s6
EQlFduDhsaJIP9cgTVWkJPDQuj+arW9N+/r8Kjww5H+0/p75DGQ9Mcb6CLi+fOLvZJywdoAAzyLC
w0ItGyfFDU9RlRkQdeddejw8WUUZgdlFAzz1un5VRbmprKiiaXsrLcjGpaK9EBVqJyyXk6LOtIqx
vzN9sVpds+yXy9CuvT/aSkaEG8auZOu0NSIbvsoNI+hdk64djWe63ZJPxfIAv81fu+YysThgkt+f
XqaNt7L4AzRqkptrxzhz+CRC3Wfd4dv4uSbCtIWSyBZyxCuQ2lKFF4lQMZjBWtbK0HdvaJKhZLTy
D6hggl0NcmLaM7LDfnqk5PLn1Ns6o6Ta01Cgnhiu+Bp2az0V7J6+0/y25LB3j+2fK2GMRdn+BYYJ
70RiWzATshhWiz6O2jfvQqCMey3sPAT7gfNB9D5Z1z09yQc3GznsOogB27FP9U4iD8UmIp9BnPUA
BR3VcZXkaWYxSXeNzB03zmqJvoXfbFAEQe1yPAcCMUA0hOlyvqFWZIbLU+lMbSD0UcqF9S2Li2Gg
XkLhMatlgDkkCV/2aQIkzY/yiSfnCbgLtmKawaJ4p5l3UPQ8XKtnNoidk2LpY1+5/TI6IcewZ5zV
RUUdG/8nxqVui4XHtvjZMtb9ChzxAFFvlynqYDY+5Zff/uqqAYuiZ5cVuJZgy6dc0YJNiVFi5F8m
InX1opW/WkBkx7fb9N9yTdNNMxFdJNhL7xwPUw17DAJz6mhg2lYl7jOo3QvAfMFK4tzv0okG+AKA
ew0c7Inkb7mrXKcwFlbJW42zQzWzKO4zo8DGs8vC31wfdOTdUk1uxY6hvUdSUIWJSRn1sYcJr57w
f1SGe0fj/ptxY1szedVpb/1vpCLQBwiSKX1ioDqDCgNn4/ipjCEr7RFRlBXwUBI8h9cpjotERvcm
eZqdR61KY7WGBsnB5jSuNPjt875aeYqB3t5F4+gmlYeqGDiJwnEQ03hbX/z7OCwU8ExHJi/Xs6cP
F3z81gLaxfIU5IpbrLb0tot9OxLpM3uKVVUw/SjINJiGxHquq5nvqpWDBuJKpylSxtlT2kcbVKic
JNXkW18QC6+7OnWN83uPca5qLFDBLXrv1H4+pX1ML8Oy/nlZ7X2yE9p1aJOiuabHrf2kQiQL+lGz
zolcGpxoQ2YgWEgQg4Fj8aKKaEl206JS8QlJ3dguGg2/C0YWJ69WFOcda4zDMfpDkOeje1WbDigi
j+xhQxcD4ZSGIXIOvLAqE9pMFCryfUB5NXZ7PaatXk1as90fYxCtKvHXZ8aPxPfctbctjBN+Wfdl
79hT2MomKdEI9qu8auMlCZPC1dCLlMP1fvkIFii1AgpM8rzAianxBPemB3gQYsTNFGfPKRq6W+oz
RemPHKFKS2c8efJzD/AWNWHlZnBuWtJulyisoGqq14oBz50tl/Rgqcnwf2oV2yOYRvQ5BkqPbgpS
vAoxLXT6aiq+n7tVyupkApYGpvgCuwhtMoPHtSCnpzAgj/cXHaccg5WSTRezPeAj3sQXswIvFTUf
RaSJW7BRYq0f3V3t8AhaWhNhETsnsDR3OWo9UTetwjs7PDyvTgvZbowj23bd6kPMCq0xQ+pB5hgW
HQfz0o7sgaR7rnCSH2UnB+Sy4jROBfgBJtrKw7BBktLXqu2bR+3sxluA0h0S22wyWjmWhGA4ree6
5QX/TnP4R7Di6A/cWmXsPLt3jrmJR4JCYC0j/n+YasHLN1SupWMU+m1xKAALkkrwwIWEqaMUJEQz
tF6EY2IaFaT4fT/4D/wMctHOg01GO75rgAFXbbuE72l3DtftYtE+hawztlwAeo82G/LAMT4wvfGm
lGpY+tim6/SUpUuWAIM7XAIKRkM8tIZqLmuLx1MkwWcSFGD5bqUOrG7nCd0QGmIoOt2+2Km/jilf
OIYnUK9Z5RantOG+ZRrERiDue6MDOGucjy1OOmC74QSWzws1nTyEtMkZsjYALP/9eJzBt6X6M8Pe
50Je7JmLXirFxkBYcVAbr4PFSpNk47OQCZFb6unLdJVOF4TqPgQWhF+S3R89g2VHoaxn61cKcPWm
uUiLsFvvn1YLVubGSGOH3009xcHeWgrbxwkg/HjRN4+jF2ydOtk6NiOE+cF7HP1wrNakXKHqFJHc
usqM0batl95Txpud/3GMKSRx7Ia4BeGAM4xV+Z4O3hnCRaWhoRVBWa/r7oKRpJLPYEadq1VGAqaH
A/FINg62d9iR/aJJwwo9d5HJ0desqLPsZVfLFVJMkhYxQczdELcqR+rVeIhq1EMWNZ2rVt3krZLi
Ei8o+ZCXlOL0OzGQUJJCh+jvqRfPvy/G/6Cr1A84YNY5856y2X8sdXZBJRdO4L4xf+sC/u1b9HU8
m82XGr/69cJoAzThZ1x6/pRSj50fhWpUQ2+hHdyYdSs19+PlAaA9MywIS9cJWdFdAUhkPHbhxmze
uzG2DHtjtRWyVo2s+zQX/dZAgtmpJabqizm4SGNOunwOXTt+WNd2TBsJPmRlNsSV6oFTkBon+W+v
5qLNYqwRTTDusCSQ/ykESgO7XYyzvgaqvevh/8PnKITp28Ba70ExFKnkogYR0Jxyu2tF7JBIW441
bYuf5ZQaeHt2VVHxLW5/sLfPyneFXx0GESkPpZ1frxQd+tnI2XHxVWYoxULpIHgn8VUAcR3M7b6/
yoXK+H9yPniGfTzCfz9g99JE0+EZD1I+rzM4D2KWDLBWs5ZHzAye2f1iQWkpVOT2CTDr88r29ae8
A0HBdklz9tjAeSPqDj/qvyUawGbxVZlMK1eTU440RYtaZm/hydkYgSahyrZz0tpQHgHLxKxSh/8F
2fbr+CYP7f3dkn5wzsGoVHkS7WoUMw1RIah2kTg5xtUwjPdYOs3JJSGnO/DDxZNsV+K04d5Fwiy4
Vnz8o2Qoll5tYor58uSZH27MLAFzj3pfNRDbg73HANqgPOkJIgY/GpLNJINfHwCTeQjzOWoTg/nT
saHm/7hX4Y8mLuqKbVoumyYjXgwUj8YQH1DwQ1brXXO+GpAxblGnDY+/roLIrU+mG/aAmQ0u0lFG
yJMraxdXDAnRPVe1s5PEv5pIQL2MRWFEo5sED1nIBlGIxiWmO0xsLcGNOHy/tysCRGrzCXkiJrIL
LaLBKBIZ0FCTwJpr5HKXOm4UPp9Wx8n7Sp5aGPd1GsH224+GiyXKu1WZCyRbQquBPLmWC8fkp6/D
ulbQgKau3GeyhmInel+xOqljJ7opMmKgf050XwCmcKcu/o0QNCIXbGuT9uIp9R/JrEEUBFDbIAUD
AFKosKPU+Dh2Zz8LwK5HvTLqhrK9gwpxiJSudEMDuQ2Rek12ttTaAdyBcx4VKOOdNcDqFFDqnafZ
iJxDif94LnIWIvkBYNBCASAaqJVrO1Fg/XVjAVeDG5k3MfD+kQ5wHFX1rGrdPPt5+DyD3UiEyzsj
imulnkmSIUjTEv5jJ2xfESS/+O629XlVpw08I7h42m4/KGNDEoGmT7uewwhS3jp/NhfsjOav6yyF
zuLXvY9LpZKhaygw2TKRKMJHC3lyZ3zaGvgQm8FFhR+S+4UeNxq1Eb0Kx6ru7DhJDkKdZ5B86Z1Y
MchqhkbCqOodn9oAKC7INSrmXfR9NZgG8AaHOQngIMCON28C/03sNb4nml3ayFrUe3R8U9rJuZzN
LEwxa5L8a0Cx25IOW7IMwaKDQvWc31Scno5fCfG84a0XP62beQBL3jgQqiimca1w5mBhWsWxFXQq
fJWwAPPftrXwNIW0qsufiZ+D0LSRH3IHU9Ucfps01+wfWXplQYTpe6rGlkVVS2dCt75L0IOkZu6w
K1vqXRkc6LyADxtEE1Ip/vnhr7H937Qn58RwKCYw9lJJ0iPUENWslYmHdSo/yh6iDgzxHB171tQc
336FWF0q2h1NFUkdJmhUZsqrfao6yvteUhjIXeixq+Gk19GFjCjpXAKLF6uyCO3vQ720f1HL9AzP
T06Hdg6r4pQpYyYNNsZJS2SN6Dbx3IWiCr+mQMGXOAH73WZCWG1sbsH7AmbV9RZezMi6/aEYAZI2
cOt9shV36adUBcqCgZoblRvd6DzrYdVCt2h4doDUuhLRIZqbnrPwJ8w2PTum7P5Gesr62AYImVch
wilZRGcXapPwxYORd0SZNYRMndq49mhST4OtjlZNi3wQjbHpTUgWim7pkoz8hC87rG6RubPqoEHw
YHMxEs16XM+6XgLBaGhOJ59rNZio4+k7+VW3yllNk6HJbH3zWGyKWteQX2QBfAHiEhrSbhs81LAB
6vb3To6C4hMsIetLPDRWKy4iZyeTVjjwHC35YGTG9rwb5ztObpldvlGi+H9Y4nOBBZauloIFhD+L
e+86nM/De9VUdLUWXu5cTr9KCACmHmOD1W3078Et7TYgrtO9+pdV1oQs5+Cq7wOimoNWtpWjbOUr
B5h7eUfV2h3YhgsXcTFy0mzj/hL7QNssSnZw6+qnGrvsAKLnI4SHXYUPebIkNiaUJtBVo1KeY9hX
GwxX1HKW+3FDicBCttgeFsWXJq8ggfZ/X8p2PRB5qovi8nQtMTFIzBAERuH4CLwGfuDV+iUxRpOG
FHLe25ZnNyqI0IyhriJSF9uSs7ByBaU1zj6GPNe5gG7McZveUu4P9exujBTV+pPq0wNknDX31Wad
1bBsH9+TQziorwA9h7SZAiWG3NNt0CIYs6/AgeLjH254MWbYjbPcvb4mUoYvAILt+d9HsPciYz61
eEENL4z5w60xDDkUvbUj+Ey5+n30SSQxNnNw7F6G6A6fuUiuz15MIBY6NfcOjHAL4FojcQqnlMVd
sjnzVIklfNtP4MhdWZVd4JWhE1CZTO4Q8O+NAYtKhkSy0GQc+go/tVcnP0r3IXCOIK6xO3UwlXcz
3wYnCN6AUKYN/jGGI0ixZ54g+wARDQgzjJnXHBEc+WmkU5md5KfMVUNPGhpV/cetzDaWzu9cdZD/
TrPj91aMVHPhTVOv3Y9sSZTNXrOB3++psXsehNET3rNj/wcj7bCfz9yYZ7wqjzLFEksj5d9+wi3L
NQfRs6DxoiGEfWmwK+NjeP1lDzBfdlJeNZxOd2Mj/kkhFVdnoO19mPDLU4XcyDsfThqQPfwNpjAa
yAIYth5NuP77LEVkuHufNMqK38QgdrygK2t+zj4wW9+7yWepJ66spAjfbF72g9lZq9zivUcwqQd/
ZHIuyPPzIuvg8NV+m5F/hV/X7UQMb43vyX3XxdVDBXgHiXnfE8X9EDeGGHVXTLc7pSomPz3qcfvV
XsV4E7cy5xBfZjLLB2iHO4ikhzgvcPOMWu4Lkhui89rFoAx6BUkq6GMN4Vfo1QAxPH51tpqn9uQc
aZ8LxREBVeF361JM0yLAgc2IS4Rc2hcD2WC58Lm1mAgRew54GuSGLkaFJc7T70VlTf0nVDOPj17r
7CSa1sMjUKk4r/XPHhJYcmrrGWZQwrXwRGbitKSKHym9JcB6JedXvSN0tHfv81fRD8JvWBwUxmLR
DQQeUe5FKdWcLJMYvyp1QGB39DMrm4rJb0LsuCyBnxqHdHPtEAQavZxr1Fc4TO++woH40KL3ZELP
O6RKCAbncShJOItaxRZhOvvA9HgpLlSNEHAdSVn1AGIx+GjY8f/TctgUXh6bQM1NFE3qAPVXgE/I
NHlcTYhhcEZWKjFXPMAGgMv/5dvCLjcV23aQl9aiDM4TLMwYEbU8qbpUHStwZS3R9OO1K6B5xpZq
C5N2KrkqOWqbIjxLYWyTLeaRejKFdU8z+AvAuexf2Nm6lzvH7zz5t99pxOwzqS7FbQnadZNbWqVG
+ZH4IABBV1kA+lBEEIKTTAyLajkt0ZaHWaAbA5+wIopSaLQ3kXweeRDAjn0h0zgcy1vdKKhKcQf2
7Q5yy9zhA5M3j9khMnYIDoBJBJLf2ZMkXidn4/sKcNLkqbdoi7mQyKZjDCYyi6HwfJD5sAW40KQN
gLwWU4j6HHLe24SgjQL+zYJXdkKK+nWkPdvafJFSOw2OHeL87wpqI3djUCL1GeGWJmc4zUYKcjfA
jyIuJ9Y5zYeM7mdMIgYvuqZKwJnrUBpcZ5JZENHfCfzWdoauPEoFOwm9gBBXy7GwlJ5UZ/Bkcbjw
eqpXWGwMs2EsWkf2HvNsUaJwB+jaf4S1ebqwUtMXSsH4zwYSAG+N/RWJv1TwKVHlspSDJs4yK81j
y9fJ/i8Y5ByR1nJY6737ndZlxxQ1Ma9j4fRGw4ZNTFMrqvIa3LDyARUc+RTeZY39daV6EJrpQGAp
4hOsnRZqmTI/FbMIN3GMyL9v+wtGNk/+AXJff7/iwI+veJcE0y2NbsoHiMhLZRgJOZKIgAX6xU3n
Y8oTxj3skyB8xd5yak+dPsaP9NanZWkDZ/djOBb+NX6jwMEB9bMqGTWAsQjbnhrijEn+tIdPZqTN
Vw79cmpcwhiKnRnGUdwdSEu1xOpZiE275qwojwo8bJd1HmNiz4geY50lgsgfVJVZJgeG7sVhVNnI
TMFfxwLQu7pdHMX82MOngPfwLzh7JJcTFABTHr9aPtcSrPAiFMFZk285RTt+EdZUAKmqqzdVQIdM
vs6C2BUWOuAJkTWZXmndOY90Xi1PCsk1tgmXZUTOlD9lAbPdD4zT7NQl2OrnPILYEuqq42C/6McD
MzpDEKpdVBScB39QWSpmOnURzgVpcOX8RafZbbIrxl8ZpcABAvGmSrqdWPicbvIFGxMNt9rkmNJr
VgovqAyUo+kKFfD1MH3uLqTxnC5Bl7Bikg6OoUrQcBtPJ0mlGRBFa0s6deY97DLOTUOA1giFNTOU
FQb+SUzwsZycRWeGwVrCES+3toItlPF5QFIH7gEseHms7WfK1nFO18lr90FSGWhGTOWUd4q3/Fsx
UHY50dihwuNXapfZTw27UokfftWF4epTvHsMS7QWOIN7KCyLwbcew/Ntjg0qoneY+wdB3KW1pySr
UsRcuWxWgmpvGYWhHCNL2VXUeKKBEGb2xckp3jIzmVa4E3l8X3k4SKjQh51boSjNaSulgA/UoehV
/7sBZ0MoSAZs+roByvfGhRbRZ1slvxyn+9GitpRJ2V21pz6W8hZv88NJOrNnw5x43k4sbDDgFD7Y
GwdZPjmqpyDP3DIIfuQFfcij2xxalG3+EqLdgl/wIXZDvC88qgsZdWNMkyNPjI4+ur7FQ/2ntpM2
86xtkYKUcMtQLgcc/SPyknvqfQ6OmJCbCDqicfvxSFSpBsnG2HdiANofVqyUKnYkav0IZ5/HNiIj
0l1/ugCpVfkLS4xAaFFd0IHpRcI8VFecbxOexJUm66CwrYZbpf6CEBh/M/Wq5/3ZKd3uOzZyeYTV
wGkHW2SfJOvwipw/NWJQLwALQAGVy6zDdlXjKLGNuUuCZ9x4v9Oi3lHnU9f/fiuSVwzTzOthmou4
M1oUt370VhhvzvhRdk6H+f/f7P77YYH+mjc6zfRXtmeGTlXk/kNnTsbH/SWV/kDGASnbs0SI/K9J
1yYm76+TXb9DdqfrIurdxDxPUXXb1sC7DglbaQTVb25Nw/ZebE2pmFd9VTDYOhtK46mnYlEDhMvg
jxXXoOfLJfbQDGAWOWusr++15kyjxzbSErgRzzxs9bXNHeTOyfn8+J3XZBk9H6olEvNfJcyEVVR+
mi8RfTROAc5l3b4UUWsR0ICazewGr6KjkDqgBuIs+qvb3Yf7iGVweSxuTRf1DGAfGNalVgipkgdO
1RlO4G1hASWDenlSkH8IVsijUSRGNrq1jLBt7wxoS78SiSycKkmZUEeBffo+ZQ0ZA8k0DSHFPoqT
OKfl+GA8S1IqyLNhkK6NXgpM0TlVyl8pjKEavBvvXjVdOc+SZtgQphuvQRisFwHu/NZQ0UlCisOc
8VBkaCUaM/PEvlKY5NecRgPCYmfYZ+62jSYN9u+WekZGJIYgdF3nGju/bR/QFgTkYAqkemoZSgG5
EWN3hK0/06t4ZAdE6JFkmVhOvmR6qJRWAkkLuzMClAesvnqW8qdhddhNchK/+g1HJjeZTgnk3LyY
cyxvuA4zJHriG5Y3/ShpdSUbBdHuhWcgSnZaR4C5XUWZgaD4aGDYcJxNjwaGtdtyrhz/oFm71zHx
SWSbhdD2B0ruVyP6H8jkv7/N6Wo6zvQoKaf9Hgvz6mgFyA89DFXAbVWJ33yk6Y9n0uaHTYZlQ59F
Fuhtbr8r3NjM224YAZvxIGQZvgN2jj0XagTlq/mQ22/WhEBlBOjoTYb0GIHqmsEGS7DsCjvVbegF
9M+oibkGvI5mcQRm0hLLco0a9gZ5AYk3GnSTheBThLbXAg/E1JoMv6i/Gta1Uihzk4ySI04eJLGS
0v2Tk+hrEZmts7PsLwGtDZ2cJRph+jds26UvGy0989sKfdaVvoIc92CiKi8uHvgVYVofEG8ntw1I
1eru91HFqonBLBfQvq28D20u19HPdC37yQgh7lV56/JA22RQXA6vBDlanh3kLYg1QWBmDCS6/MvO
HQH7N6GDPKt8ebZ15yRDs47Qsr/fV5DW0nQEP3t8PG/N5XW2Rj0KjW1ftLiClLVKn8UMXPh1DB82
J+Gu0vvrYBOt6w/yR5XDoRXsuI5bfuJyPhloIDViYn8IJ2vw2afU7JIoRvqtV9Le7Z7lGDGrqtBF
dBKw5oX/G/D+Mia+g1X7xBISXCwF9lQoFGncUAwDgGlLiwzSLpAFr3BseOyR/7CswQkLaoFSt7jf
2jmVWB0XD6hUI/jPr/HQJCCrsFrtfzgMSWJfK64LSHupPUzVwyUPVZfDlIh/rjwAeKm4T38kGb5s
a4RLT9COct+PFT7Qh6mq0o2NW/V8qwvDJeJT8a1JGGF7ZKUmMCB+d6rVkUxOLa1Sqr/snQc7oaLG
i78/x12uWd2Gao2ffzToW26emy8ex5+w9QNy1gVwZXUW/D9UJ/5XzbmoJhJ+j+NWjVPFlzZ3Qr+z
dW8gc7nxazplsLbh5HPL5MLiIjNrtzy4E7E2jTr5u7o8Uual0BkWw+wvcfVIleqxP98RVAO1oFUW
56IK8WC5ZS+i6w+GuzHfzMmFv5RMotjPUbzMzIESPdPBdtBEt7z7Nxp/RRRbZWKKONWdvxOB3FZ7
2vSkyQmf47BbjTTG/o04JJNFkSVNOF3LxBMmscDgcw2SghYkwFMvuEQ0wVNgyxIDerT9YWVB/+kG
10Hj8fQqTUFtChUjlyLf9p/dzhxO+KRn0vmyerINb8qmBmimLJbE027GOrTaWstsPDvkVydOLnqt
py+8VXCG4ugSPoJvMHcqRSd1Ek8vtNUQEiddzS9NRBEIhRguFZxwL4ZyvqIGBaxAG0KFZCyvM+vt
zWz9l3iJHvNLZuGX8yyhHnYaP293nZNuvcuql1WLf5YB5+7yx8hITxIKhq4a3rfTHw/c7UeIwqbi
K5OC+4hTpffPxBwDDDXHxrvJh6S3bfZn0Cp5Hglo8dT0UDj5BjCmr3ZB11QtD7raFRuu19zFRTZ4
anVZR54/voDYQhMCM/2u/pkm9etPCavVSiIdrUhfqByw42T19OTXBLqJp6raoEe/kHqiFSURkvfR
OwI8y1JsgIq8Hdh0QdWhUbTWpxU5uSr6uSpLV4YcCfBXC7wATHbmBuy7q4kybu2epvBKvwzkCa3H
P/LSwqtP59u7Q1mlf6bVadtqsq3lb/lD+0N0tNZ0YtsGbSzLELXLDbvJirP18za6/b+xJaHry9V5
tmwbz69zS3Xa2ISu0uiV5mWnKb3WIOj9ww8uAlQkgVk5gZYnTDNrc9v7RjJKWEp0VDnDTsjxPGOR
XfDDf7QiAtrYqKKbcTYudiDYKcD/yu1LIXC9khR4PiAlHRyLPbpAoz3fEwiH74W4KiP+fquJLQi0
e1fJvDdjUzqe7MTg4enwuDOFz5z5nJ8aPMbTErJKwEYVEB8vs7q6jNSiUsUo5HpSaYluX0tIQnCD
394zj4nj416EGSInGLnbrCW58EoX1KRCc/xKnnaGwaWNcNcXCxvof6nw4RgeYJKlwVkQJeNifWWH
B428izFiCOHTB/thSAikW1asq0W5NYpzh5HP5GszfT/0xFH2qFX8M+MjY3fbmgBjf7IJM7ZzM97r
sl3DKlvNc3f1rfGzfryWnrNp4jcu1sQpLWr15jxzNhiQwY4O6ZnXNCiHXa4f6jKTAs9ympkNLZtX
ehxN2l4fcANXVXgrn/OQjtHAP4ZOpoZslpCOIMHcLum01WLGp+B4i8xIA4zvbHvF2awG/y+dcNCz
KxJ0ggQPYGBJDbhgGWPLEp4H+eOUmVGsgbcOXW1c8KvaLkq4jPO+sXOZw4ohoaO0my5ScjrqXwhk
6TRLA/XVYpuq+MIPtJxEHMIQk2TsM9guwsnio9iYLTYhg7WxLofjzispSrC9hBhrduFXRqr85tUR
i1ADjKmz9oVBgRIOOrs63orNF0mxDErR19JC5V8AuBXJbVmjEojBme2h23Mw9cUhpZYq0hatCEfW
NzwGPrvbelo0BAop/mJuxh0LhBNyqUxAGqh4CIaI49BqV/oVlONS/GAS3XVSZr7Jtu6tBwLWK67J
GOJJZIRu1T12y2L2cwEuH0Pttv2PnBEUbuI4Yu+75qgKZ96UyFen3YjFhy7Rfx3WN1/eVk9phtgi
j203L9E/V0YVmtTL0ZtO0e0KaaGfXTBVf3NQuAlngea/v9fcTDV9fU38UPL1iMkav6MrwHHblJCs
JUpDFDGYVPHdcDGBXTT+hZsacWkNVZtFV0bc6+mZ5DlQ++FvSi5f2waUEOIzXioZ75kRMrRNxAYW
hi8TyGpTJIw3+cvrRhJiG/hzDnFEZt0MmZT97+lj45N18boNERRE2sE5v1vl1R86pdd45kl8Kx3Z
H1Td73Y9KShBBdkmVvqsyUrcvPCmqVLOdDLLWDvOLcA5d2/hLLRlY8D2PBhPv41bUTYscwokTuIe
kBrOVJ9PDy6Uo57YaEMu0rZ1KGZXenWVbszkySiJtRZMrR0N/u7+rBoGvpbyoYNBbVIN1iPq8ly8
RS8NTzlkkKNJ5iPvA2CWjasviVY5DAUUAtyL28lx0g5GZAwzEPRjhSaWlo9/c/bwplJ41xY5QlaZ
lWIScLW12uJ+UQkbuAiHuBxIdGOE+KN+w/i86sLyaCl3ZjyNbZxSGrCjlQQj7ruWQnZAZdT/GvlO
P/XdC24D05I/ac9LnL3o1Uc2QWelqOK8+i5fEpX7HTfoZyHj0hjlz+pJ7oE2Poib+stWltCM4fC2
SeUtMiSwWsxMWAd44cBSBQYAM76xHLERNWzVyXnVmQ0L1qa5XyPyy6pjsomhJItLzTa5wpbed5Yk
+hSLL/nZd28AfElS2AXFAX0JS/e+CeD3m8SbzyEuJH0afJSa7Unhy5DbDB+HEdcqdHlhQsYUwD87
LRpDo4zCvYJbl4w1myERsnEmjeExPQns53Qy5UDyIAjX6JlvwIPf9wQimwv5tIa+2FSqk7FNtj8A
lSyOYZhI03IE2AbFIJvIpjQxNHJmv5/W82cakcgzsWLVZgQHb3/1kxrt5rKq5g67wBGhUp/BZSKB
rc7/IZ16c0r+mQIlAr/5b6bSel4hKdf0mHma1rJx9wqfK9qU3ivp9pxXkp8xNbBXK0szXjKTKlQd
2VZl3qYtqQgSd4HgMbRPXCngAj1jhDl9qRo7Xuw3/fres+RxpykvOw6p1uVTgj+n+y1kVvSw3xBk
bRDkUci/bbt8PWFJhKz+MP9SX8R5rYjwT/NBuYDle+N/30lNg/eCcPi26WAReoHLXiIOdoYYjAda
5L74wpLUdzlP/IrKiFltRYLiiFPGI6EmTI39D48Kfp0fntFzerGmHsza1CxwM+qmzw7mPbD1yvLY
/phxrjJICNTaBdQqv2j35zv8hqEKt6wPqCT88dykvhAdZkOH5QvadaG9PZ++Gun14siGrNAj8ADn
4Y53UjGujHd/mpx/iTJCydUardXv5doQqvVsCeFmwrvkIbn+IohFjLeVgyNjlXvsIBhGtXWWeGIu
NDbCpuWlyvSqK2ctA3OFaVfavonlw9tlW7U3iShWxduvakg9F7bh9HqPetlIa4gd21jHPJcsbSJY
KiIBDZeMnzb7/oYVnCeRufXOjciTRW0eqJFwAN/MuSk13JOszHCZ6oByAHIFU0wVQaVo+XQEmLI0
9xzynrWeRbPQSzPYAMYUhbZVPFIqSF+DG0l6PRgHxtd9XMPA0ja/MeQ8uk6V0syu2S4Val1Bwk+N
JlButGNCD+JlgkfLW6l0JPvhKjoX2c3LECi1/ZMvZWSpj9eYYCVsz8XhhDaTFQ04bIG/xDXjgl2F
chNNSU5NNk51zEYB3kxYaC2XwPQ87jkPSHkMDXX00fOzE06+nxiFvbn3aeZWct0dZ5lZ39OZrpDE
Z5MkqWG4SfKvVKtiahMIkolgVgZeNrt0Wzgw5Aq1ZK17d6QaEOdC5+ataRyfhguESsbzBwj5eIgz
FUDGe8D/iQhntcm99K82VWyXnv672hxQc0mqWR8rWhfCONQq+SKz+/LjtTlvUJ1P3zdzDDgzkVzs
BGfoz6s4k8m8O3/DTTyklFcYts8+wReQZyce1Gu9DQUdsHDmtXiZaTAzrP+wz1fhm3eWl7MctuSC
OlovyihnG52tuk2sO2HOEwJm7P+z0mOi+2qvUwtZq9bNTAEhL4eFOxldXZf7fCau+Z2/sTweOSIH
oOWYVs6MZSdCf9xX0vFHB/g0QRKG+obFhKBIXkZ0XOzxNpRGTy5xnf3WrWpOZ0j1QHYVOsd8n12n
bq8aIA2uZ+Nd2oOQ/NOtgv0tH1TJg0tvL/j8ePrTQA4ddoiBIFBHd9qaC/pVZ7R3O86MCr326zDT
I69RH+J19F+94LwyMX7o20dFRk2qSNsGO/CqNzXdKXMNoOFwHpePC6GnKip86AsPczf2+p5yxlNq
2l5m7oIjXB3aAYVJD4qZeSE1dSlgvoWsX/ukNSefvmnEBuON4GyjPbflddZWdKfCgcTi9aDXnxtw
kA3dwubB8bBVTezuGFJJRbIHm6CBPp17ZESLZbW5zmxLoDHP+Gjtl7rzO+t6wZU3qvnadwTj6H+v
5uK/wQbu5z43co6e0xAVLxPczoLQu/mxslVNijxG3mrjyZTzJw75ucFZLg6TVADr2XyIFyglEDBn
DwI4B86oCO4hnM7j+0BghAS1m/HyLCHjHGRuHWVVsbmtMOKWvpesCYn7CXXqCvh8xXTcHFmGvk8e
DGnwtc+lgXg9rwZPUR2GZ3ux4tnVm46uBxAyRvrFnfmXxtbeMv6zuUD571i4qyVTHpY/kc75DyLr
kHYg+PZgY7Mi96JlqnPmLNbBEofNxt3BoZDGr3Jbj3wmyKj+GidHwUHBKMjmpttLoN/Dj1KNCcE3
Vt1ZmyHrhxmi/JH4g2SNWotVkrDhAofCjFCjUhVLLGrj+8NrBYuth7vybpFJwewyAi5ACGGGcQM/
pMNAwhmUDFys0gSlpn8xE8NevxUr1rfsEc71PQRbR9Hguiq3OB1zZnN5c7zNyvZQHOEB+ASEkTXT
frVZ9HF/bNZCiZCd7EtSA/cwMW9ZlydJSj8nOyBoRr625bpevt9+fjn7yUNTL1cngk+BJZF2ugMM
eNEeb89QiTLaK6BNRvYYQw6w7XgwcD+Jm2+ERQYtAFbQtVlRyTQVAnqTKbwrPea6wy6g+JZ960SP
WZU8I5O4kiE5zWwgkzHqwlk3b1mH2/UpVUe8wqndDOwM8/uDCFARZp5D7sUKgOOc/f8XOTOSIWjD
vaAkpAN2Xq/4MXb2TDifYPZv41iA+3daX9vjQlum06XGx8qaiZ5c89FxXcnLtjyNdOiJd48H8UaK
Aixxeev3TZ2pm9koCywY70PErvNBTr9lr+Qby9lCNBlb2Fv8hpHsPrI6XMnSBj+2fXwb4QMSwbt9
AY5bsmg0zYtprSZPwGQQVyGealNmadKLvHYXxpk2OaFIMfGmRT5AiNEXtH0Kz05URedWyGvW6mq+
4gWt5+Sc6sqeNmySVo917bhFHANY8M5LQMCD3jGG9Man7wO0mZj8GVOnOnt8Lpgar52Gmc+nYszM
wMnUXDsUBPDx1jXomWKQH/iQHMPT3FOzmZb78kaFG84GlKwy+2eiBaH6oEFd/1ST/8iOyZ3sEaS/
PNvaKXI1AR0Q4Y3IjvptwknLhPNQ8zpEA0RiabSLVFpCpRyRG/Ff1LqFVhy/QU6Z4t6Tooe1GDK0
ysX4RzmvrMTdgnA4ZfVLR59ptD0CBKxVFxgNze1faZ2yy5ha3UcST4GbTByyLBWvkChUFpn5yELO
Q8GraOufmZ+PirBpyLHhl0oaowhHXa8+AVc/DhAUbScqEYPAiFCXNiFqefR+YOdzVHG8KHRDa/Fi
wnRCJGEV9D2GMxFGy8NqzohodSpjm4G3IaU9l46QCFsq5tVEjLrgOF0upSVTNDkrWzxS22BtlwFU
3/YqI01v89uVxBTXnN0SMjPv41Bk6i6b+hnM7LR+92lAmCw/8QAX8Kn+TMwhcU7oSPbs/Sm3r9MC
PezWcDlUTo7GHKTW16L7mDsM3HyOXv97zWlMyHqo18R5d2SFDYhkRSwlxX3Axhw1Vq8uYfVeIcSt
3Wn2krgi8d46ECJEsRYjDpe96PHPrDkpylbmrB88RumjCllT/B2lmsvtsed85SIxfKT9yasjPQxR
jzdGMZTbgaYe54owI+zi2aZuSPp6DiYh2fqCYv+LF3Haz+hPrXtoVUwW/+ZChQGUf3cwJ063yRlb
B6BzzmVZ7loHmWMhiwyoNiYlVCq6Ara2rEkm//I3HgJsgEu7NPUhS0+RUu6aITbizB2A2JOOiZ+E
vXrVMtz0nOx8ss76wOnXGjNM2Je+L7FRw8PUuwyUNUdPdzgLaBS3J6Ps5kFaMLKlujOB3tLrIP/z
E+jNoqoCuU35H0JMI4nu8qcM4IhMNqEVHsS47NvdwHE9oHkuIIG7mXHCCmgelaYwXDt+1WTL01mY
h+MNRDzelOK/c0kr8ZNZEF9J8LXWYIhHLtZrTZ+VFYSDMGVH/KaEGKd25n58sarI28DMNia1hXOE
IxJv3d5AfHD8l7ZQTmCuCf+44/U94u7njwCi/a9i8P1u0XaXbzU8tsAWMrAXtKzZJcIQgIV4j9P/
gB6qeqGUGO8VxiE+WF0kS7UHRoDN2K8cFgZhu41osChM5sI/JJJWWGUp8cuhWJt4hraxdXdBvdSv
FIjaD6eFAvlE1svrGsC19x7ODNtMO3xrCXy8G7t8pKaqVMGIGPBUpDpJwGK7YGw2V2qw60RfK9T6
w18bngoiDmIwxcBrEioey02THfVeIbv5YVFDenAmLOOcY0H634orctjGftBOljqt6tCapCkXj9Kt
QsHFZfnP++XgvSKydIRzJDRg0SoQmvggNO7TFYxC923BFBTeXWjtCcB4R4ye+Npsxv+B4hyMEI76
zZ+nvTpzhchznkTLAdMxmhdDUw/3VQXQUhZVfOQIzggYUlwTH+mKNO/2jv4ol1I0r75EpRQVGHP1
cFLkSRFyEEVe8yvw8WBanHBK3pPH4B7CVQy/aaPNdIlIenN/EvIe2hKOSndpKm3X4lCv+xMsB2kD
URuNQv2Cdy1uotfiLyh8X1NtzWwxSiEf+ICBrggBoEIAq1XDopXTK5qYiSMjkcB3tonZ67DLb5eW
VKggAjkpmPWyctIM+gO77pmsuOmVGdYu18TVrRB/C9sFLYmnmwgox2pgQ/YgKGMUT5eURLVJvN2G
YHMCOfGLVirz6WnW50pNXs6SpZ0tWkTn/zr5rnwUgdcEAYqcb9PCFp2GWzQ7AJFVoFlkWbC8MCRp
dTgQdPcaHKf8cVlrKRcVJ/mcqP3J4MKjrwBsELTIHIzfgrml7L7Fu6+bVWi8FNvwf90IQ3vM4aJi
IIDp/Wn0rioSKizyrv7xXRD04b/z+m/Y0/mv/kTrK9NhA0akHA4k6rVjVU6edZIoCrk9eS8BwiXB
j7duXaMd81hc5zPU0E+HCKKL67Wlz+uOg08oORw1z3X5ycEiHJmCTsWfvJqgwhG1BfbrHGIjEM5E
A3f35j771p8yigbbg0RkXns+UP80vKJgNIRu7gMs4zm3D5wQtMUk39gHDpTtCWfrAGEg+JjzNNBb
OGsII7StgsiS8abLRYoGz6LD47io/r+XwwK9vMNeRfHlS4eD0eNuHZTgLN4jZUSrdRS1YKKBIfeC
o7n5c7mqMKb9NQGtsKSfV206fiB0KKniK1npmYkDjTyWvmOg7Kih3OBWGyyAcfXuX434h3d0K12W
xrzpFrr6svGny0G5GipqIvkTNJ2aLzebkblWec231fOG/wAeXOkzYvu/RpTwlbvkCFxBGyTHb15+
/05d/uPv+l2f9bEYY7E+H6aoQPjriZDrnEBZVmRgxSfyqIRsZMV0nQ3eOVSrdpfHQTnua3tGErpk
MJn8W5DqQ7GH9TUnERj1WoXhpR+jrJriy4GlJfRVla8bD3jmtGk0Ltn32TOfRvtRcxYoybr2JR3U
qQq3pWTMDkBQsb2i6wcK36eSIBPgc1QV/G7kYfezb9f21Tuy66Dv8RrUtABIzIkW9b1/DGcGAuHd
O/URv4xVfEN5tZRDYBsahI0uZlKJ3GteQ935cminH7823BRVLyrrfHnZvpueAig1QcfgCRTzsEHE
eMvJzIBps4YXxHh9ZwfB3zJmGcdkaXUpqph3UAFQaRNoY/dhPrPflRQZpHAEd0T8qU6i93AUkNmj
saOpM2NGKPDA1E8k+rLMr8ac27psGZfkIH2LAjTp6TlMULZcbBUmUPLAiIosEnWOsdvfd3aRL3is
mSnn/QkhgmI9VsMCD6GU1w2j0/ZyXc6bLjM9v+29xT0syFkmG2jSBftS/mFXK/4NVYck9J6jm/q8
QrNfEqoxReuu1aWwmHauSdbXRiM/aAwJPUeGmtMBT06YM/P+NIPSpzkaP/2XBn5bAoj0AMTyuQ2c
5czclrtKKuu1hidjWQL/o1wd1634KvLmcGV4fO+5WMS/q/ZSfUKx5tUvDol63h/gRzxIprLoEQlo
iEt0T6IrQSI6Oqa/KchmBnVjsO/4m56/zbWFzx5ASp1WOwJcyy/P2meiY0Cye3un5AZHSOYkc1gM
G+dBuJPhc8ib3sjs5gsQbJR5SzOekqY3Ym9DyAFTiovFua9zh7fwgV4ZKdX7cA7Fg4oSALYiwsAM
6+KQ24edMUUPaXZhW447bY75hYYe6A3opNe2iqbvIapHj7Z4DzlIPei6YpoTfhUxlm6UTVxhdied
cENFwRV7bC4AOEHhSlUEcbBuC45iQVHGdUSZNRdaQNWXP/NRVJnFNIIOUwPxn1mN9yo+r9HBjR1Y
fUrAeV2vOLWUW2QWBDVoaJ1neCTxaMHjdkNa1q4bHjpXrf3yKZP1v5tASA1keTRH7xrWP41tIrXX
7F55pFRs58dA5xE6+qUIb5PkJAifOjEfMxK6p+E4Au6vfu73zQP4ZcRc3qFsd0J7zJeS+P2/+FOy
zTwYC2Kd+m9GbK+8v+qAirrG+sBPo8e/vNy5gUuogKhEkrSWvXV7l0aHrhpYbrGYWNDMgwRD8uO6
A3q052RiIV66V8P87z+o8pacTltUBTwrvcSR8zPSOm+0btltOQWbLSymExyhNDZqA81VIbCmOy34
I5qudmAJDWVMBeJ598fySe3bY4TsZOss52yqklneB0sEOW1JpJnNEeeapq2SSCsrL3sVGo0LLcNz
pufuXChNOT68if2Ex+QM1ch9HfJdPTFl47NtTqMVhPjR3vgKbI/KuU9zLkrPFZH/fiDZ+ruxn9Hq
JovRAJ9lagRZyd0cjNoQUpt2nsMtiBx+im3h/3cFM1yJfZUiI5BPdJBGtM9Zg/nNkbWqNCh4vMa7
SXU3tqkB7+JLiiIVW9Z9e6pFG2DDrWce0ykuWGZ5+FJ5qHQiOYzVXuo3ByeeXe1y1+bYf4a9xO5L
/NDzHebzfTEnrXxDRphrLui0Pq9OOizT2Xb4VIJCrf5WP3oOkoYk6UK3vMC5k1a1T4mpX5H2O7AF
97h2uOzypBnPtF69od8zmL/FiFtfHSFNwyFXIrMUqVbjSy7QImtC0rTpPkINSd2BCihJtKVFfpF+
tlG8iQt8G+vT/ymTikLWqnn3J575mq2V0QwNSDJcwGnKgfr3lzBpAyKtaex2tVbeChOXzZjYW0gK
Nib8JDzDPpUBE4V4prEoFVPF8qufEbL3eYFEoM6CNBFs6QKhzLaVyAZlqbg0za45bL/O+Qfc9Tf7
ZAc49K1Q4k2uwJ6TGEPj/K+kClVf6uZqoZif/aVXtZk5rnWmVhBYPS0vtKIoj9AooELwv1Ep++X/
UJMpmgXO3ie/livNiy5epOk/Psdld/yTSQJO2glPkqWarfMLOGgdtf4NsDDpneV+DiUWOH39UWXx
4Uwqhc5NS+Ic+HLC55llVaaDV7Ev3hXWSOmwKs/VwJlpJLctwFRgDqZ1O6xiXyuBpbJcXZ5fhlVP
9OCE0AzgrAqBRApMOuim7ylevo3IMT/6TEZLxAeztjw2bXYjfme5jQd/Mh2F2taDcmG6vyKeKsMi
NrpZD0sg4cNX0/Gy/FmjGsK1Ef2Y6jDGh0pHUXpqYaYYWBJZsiOnvCZH+Afg87s4JW9iVMx/pYLL
wXBgI/5tcDLR9rSyheIFyx6JZLAf11jrz6GexHJZPoSV9kilBKw0eRYQM+ZSfroRWoHnX86JtLnK
PYFBEuWGaeL4/b+ofnCgkaKFha8gN7TKQtwt+7gCsAkvRN9x4LPcYkPRdBLfQPRECIJtWR3OiVWP
ZyvuM9pmP8NRjAO8gT779cpcgLxuxMMnD5MJCqGXr2BynlFnAxRARL+ZT2zLxZWqWGgbE6kL6gBb
qHAKlMJh8kLWNDcf3VCyRO1k3zxYqNYxUFpU+I/pWejrO5a6qIRoI06YBOLmLPWqpRbu1Lt8p3wu
rubYqzLqEU9Zo8/yiAfREVW9z05Gc9xudEGMa/ENP6m+Pq1TJOo5g+MNtEhOtNKxA1sA2+cSEufo
KiizhL5h1hGi/xpiwDD8oGSDLUo2WMIkkSVO0NoDDXFuWV5hzawLur78rsApViMTKAB6ex5LZfjX
3Z5C4A3u4cbK92pCVqy3xevemUE5yrMBM3+ciWJcI4oA/T/1mahzTTXt5/imCIWkZzSa8fd6ZCnp
Tfwt/uZYj+/rErgmFDqj9AKDApD67SArt8zizgsSvD+8tqQN3Z0Plm5as8MA4s63DRgGldTjA978
T5s/dJDVoue8NfjEHco//o+GMIFOwqgD0NMG/NOxrKoySv9etsm3mzJyGXhdFzNMP3xecIs6kem1
C010uTnvn/rZFec/PseNuOCdQsTgbQwWxylybJyqRusHLjX363B6f7ejbys5D1eIV+RANdM8GKLK
jyecmlx/wv7JVhOqkrVmVB2tqw7AbKpxUvoACrhweZgdZ1D2k2TT7mJDVGE0irFTS9QRdde2vAt9
AwlK1rgHDA/+0TZbBZiK7XQSO2Nfw15ZRCWPlzoeEf37zd0EpFdcsqcJs4Hup4u1QehJtARjqprl
QoEJ+/URc7ZwoU5pC+F5vmfakFiIN9m89WOLFg41VVeKSdmMW2+EfaDdQ0s9Kgzb8hmlCQ611txs
Y7f8K2tcVzsdumrTlmcSqj3Hqp+trPCPvZaovqlWnKenWFKoFI1TFbYYe01oViYaveJQwXTYX8+t
kmHu10AeR8V07XIeKN5W8o+h6YC1sLTqUoDu40LZpeEYklZPUGj780wFD3M8QXyGdeLy61tz8ITd
RgiN4z83TGAx1+cmYBwXfIg4tRqzp7RY1Vx6JyuapqyaHqHJLoFtjcxtHFG/6xkWkXib4kqPBinf
Qr4dC7IsirACU6b85P/+LIZpHwYj62a50YZHsmfsrZ9qpwWqrzfwd/ed0GhIUiNaKAVTbFp7ghki
HXphWfwRdomcyCWrQJE0UW9BckfNOuJ4hgxrpnZ5mu5L3Vhd/52omqyBplKrWGRDjvoFrRHFCN6u
WQCseVROOv51BbbSO8RM8qwWYyApqdufHT6J9SVnf7hyFz3Ec27+Y7vioAIWn/3jCTDFXfe8SY8N
b6UwyeoldQmSumH3XywoAVYZLnrn+uvikgK1uJWLtM7yJcerlGCD7LPMI3exsQ+kAwmwmnVBh8QQ
GGxL9NW6Lk4PwmGj/xpK0Xdd5Z9uvpxh2n92oRz4RNdnqi3ohne+1yjxnop/Bx8C/ImdKPqRkwCd
G41+/4vT7CIgUNMjvBRdN8tTWoGQvZ3wn6Md/JJXT5APfiQd03AXpxqKUWOCvMSuq3Hy25S9H+U/
bOinShFAtBVkz0I82LkAq2WBTHaLXuTc+OHx8mfH8zuIEdHRxyljrQvhKCZAbatIFs40kOTcCJJ6
sx8QV1rz7DvcKUNm8jbcdVLQqiKI9eFB5t4D5JZdEUXoNFK4tm53Qclq0e1k/mYHBvAepKADD3Mr
hxGkPWkqSyWtN5ymr2a8kSDjR7vwl2TjqeRESXQC7xIWQMQlD1tMm551CjNNToURlXPbM7IBDFAV
ZA+Zc1Dcxsuiib00KPnwZQj6Ippu5HOwb96KhwiBh5Q0ajcSzfIGilnpis84bkgjHAC1TYVLLNd5
k83zCZmIiWalv4/An9V1bdDuHn/sfZAlND7voWXLDo9hf9zN6V2kRkqdPjc2zYHpUvz8HUUja6ll
Xkpr/mnFH3IQfgcO1qiaETJEytgwX1FiCWLn7doF+a5MW2cEfzs8M7cNdmJEc35jGOsKCN+isOJ5
a39evfRrFrQ4xeRQ3nhRhC7vsjEIDdLe8qbfyRKiJ66S384/xa8r1ID1nmvK0mgC8xtrcI78brZp
QooEOFlbQ3CE9gJ3VuufT1aA+/59pdHd0E7Xo42+g85aP7OAGzW/pgvhom1Vgm6pWrYfYiG2uWJ9
8GI48OsPD+sMBcxHmU1A5XttxPzSTGwkVrfFZ0bfN0Ekcz+QhrWQvDLih7eVmcUMFGHAaVCDxVms
K0463LZLccupsp1ppeJW4L9GP4kUmmi+jCXovAP4VdIcuudRoesoxGMG61m7m2E5WW+vZqwRUDZZ
tlSUE03K2vjpN2JiL0OfKYF607wwo5QXfGCTmE4PjFcnlBe0JPrutrzMVpjcP8TSfdqU59QIsOQR
hhL+inUcNU8ZfNEW/GGXgkw8y6kJpn2OpxwjfYFjr9LZOT89kn0aQbhVEpb0/FtSbDPDRCAoDAf0
ehv2k3NTc+pL380SQLRfxMCx0SrmEWZI5De/xrwrn0gHHEy1LDwFSH+hkp7fhnGuqQUdENPqeorS
aTtvlebg/DSm3oIdp40okpdTU/uFMEfFyYgiWiMOptWVNoG1lW6ciKwrQ+5pCDfT9SYg024Y34E5
vPBsvbPVRdnsoCMpec9XdE4wDY38Um33ZO2R4eY4bJcM04KfnE6DD0CF+eG8xFBmrO60Hiv4kUUw
y6CWflWGTwr9hJudhGvwPN+UgkEy5wAsAL/SYzqGcJLVcdxaBdt3+hbcg5ul/ldjcy6vadhgoVrf
G90l0GN3Cu5SlYUI0bacvJ/z6gB/kpVbfvFCtAu7PU9bfEDGSKDnL7+T605OEIdbyYnALjDsey9d
c4V3RpN1p93/eIYAt69R0mRiSBy37EtW5zi+jv91e83i8jHfCCXR0kx+CPv+6TGTiaC/84rrdvgI
55Qj2el5eM+bWWiG6lOAUlpjSwXQbMi8LwlKyMLMraX3LUbuwSUvImkwYa7bh0bqDO3lopDKR07m
V4M5tbtM6gtyUdq8ZOyCfJP8ZSUr2arrarJs/t0Eh05vocYaFBcJEkGnb6si32rwCXdWvXj2J9dq
ECvuALGHRdgD6j8KHYSDgZ7CwsBR7f2OxIXzTmwO2kU4CVRXXJJm8vlaN8XZWu8GuDc2kJeXNynH
VorleRkoGCg1JpThSwix1tCCtKli3RAkfIN1lLyYIVM5ggAPA/7Pl0YTnqoRV/MyFLLM2ReugnER
4Hv7jBeSJp5cvkWUkB49Y3GIIjhUpF8rk6Hn/w0yNc6w7BYHAaZYpwgsUnA2RTcp06g958JKQd0N
YgZurhQD+3kPBXFCnFbpRplp8NvJlJ61Jw13TfQvfT9cVNuThPJfSxJBqj0gJuYPMd0B/P/FzjXm
ZTa05eWRaLbioI3Wroqi1Cwr7EyOaJxmL3x5lUE5nq4KhjHIihywAlG2iKDQV0OKFczqEvErvZQw
949n3WmTejUJCpm+EAkf9DENZhGIQM/KqBCKV7mq4uPfI64GsmkTrZKHOizuiz01YQ0kkdtZPNid
7pQT47vFIXuy6JoWfj64sTtUX82uISkd84tNr415bDWggRNWpW0pM6eCTfIIchhI/5+wqPNEUiWc
sJfRhmAnzhEhA/8XVBHPPbjCUt39D0YncXqFeOVFuwqZqod7ikl9QrjZIu2t/Ktcb1TtXqXLlUEt
C7ObbMIvJGxqco27Yp2zvTLD19wLNDkuvwed9Cs/+bfVa6GZ4SkTKl8LuIftQzLPXriBLMoMYSnI
q5KtlSjRVhM5GfA0rEP4krgp+G6qZilAzHbczmfX9e0oFQPwpEQPwCpBz8kt+1ga7OKhHt6UD+aO
NHEDAbO0qYwQViHXj29i/pItYB1onfHQLX7SYbqvIEPWWaZRHBSsJYHOndWEC8alkByKfKyYIfZ6
DQQci3rF0VKDzDVS6se06B/7otJw4HDhX6r7vr3mb19Q5P8nJTkBNgz7xRVhhisuMOSDs5YlRXZW
E+b1p9YFtDhnXrmWXaHOIu9rprMHyQZnrsQK7s8QCt5rbvgutUcFBrea2Ss0ThRUa2rcuTyImHSZ
efVS61nNXp+gWkzmlC3t0g/fJVWdsylcFLqPZXoTiFt6O9AQrOmKORmdtnGBApCxOcCqRucDNG+f
5bBZGJ2Vno4mAH/+iwWguEMdFKx1OYy/Rmjtxi51t3pKIjsnD6iioGHY7OlobYhllrZHdGY/khFy
Iz09Yn/QwK0P7mQ8gsTE4QwWy7jdRgKwnEicATAMcEkyLtjn4xunAgMS4FNtHqOXCNe1wKMeJA6O
Q9xH/nHsq4T8t0r2Yfw1DLrXqSP6DU2o0L3b2CAhTf49/ujSis+knkkzwhwdqydXTAab/jbMqhDk
vD5oWlohYH+JMIt27hOLWTiDd/EepQ6pu4kTMC9LeEe5xFpImEe9ipeQZMQ081PNdZfBmNl83HKR
e4gbllT7TA6Zfvsm0zGBSCazlkeZR654McChAPFhqDePtqTT5uu2QyZo/ZNn/DQsocOYpV0zAYR8
dbJZtizXHtU8bMBVIPbzTYRM5tOdFeXSTywc7Jg9BGbs1A3Bx3pfsze3YqyzfvKQOs9fkRqRr2Kn
34JSCTxjiQxaX+ZjSOOjpQZlL0H36kAemLVuDch479bqYnWXLoK0Ob9Eal4NfCwq+g8ChKD2em6K
FZIbG/y08EAF/QOvTR//vocp7fDdezkg2nCgUrN36+jxMxEkqtryxJsao1Uks77mq8bZrnPTW/2u
frkjUVJ21utTNf5bnrkk3JM7Z01VR/vlM0yLIN+ezXzEG/lQAqjJH13U5LASJfcyRmBzIuwsu8Dq
FlMfEmG0nijVWDAh9CkZTxfIsmFz+grmUwOWCqsDuZiKE/n3LQkEBAQrlD4O74ciWMjYVUdcA/Ml
rwSupmSdvbQM2mgB6GFVdZTDh1GzuLE51GjLT4jk+PtjAKmOOXxHynQysmL+ZrziU2LNvAe3Lwg4
hfGIMGFA6PK3riWGZJFNVI338lqbTPQZ0iNhqPXgwU/l5Tg5sQSnxJI643EmsHWDlLnM/6nhhj9P
LL30mG+aDx9SqtUM+Ucap2zTzqAQW+dWFHwFshv84A7o4wZhBemO5XeB+AGaavt8E1Rpap9A40eY
kPiKWt/yURvlucUcmUZvs4RZ0wi7Ddc3hLDgKCHf6Vgh3JoJtNliaYIF1gAWDaj5eFdiJ3EpW1gv
k66+tesRnJU7aOX0yYCONM9lEDVZn3u+zfw1BeqAf6aqJSGKtyC0JwkAL9qJMl54fEr5BH7q/391
AFZw/6NmuoVwfDEUhjmXTbhUQmmbK7/IpRuBeE2bRkpZGTZaZmCmHHUjUwwHK0vEAhiyhTqnBpes
fq7Ws2SCaANvghuRTgKglCmk0k+EbUvcmFRPan7h3Z9eBiMrAzyq1RrjjO608SQOfb77BGY8u98b
DexmVg/d1uy4UOoYVAXFpuXesyCKbZvYV9DDJ2vO1T7gARdCyOtm2dOPHPl2qsxkMi4aoV/j8o72
rQMQzeKzEQQ6JVML1yixdtJS53aI3fszygIFTSUt15t4YFhzPnvpySP/Q2giv1qzAOAGj1KalYFu
WnxD9trvTgtT/lpGr5cj7fixstwpN+1iL045Iq7boBpJk9tWKpyutmVbe4eTuTnPN90VXrUWZMjO
+kX3G01+W+YIcdqwy/wdOf/AaTmN+JeDoNzhzCZEu0j1BVryBrnMVBEWVURinzL539L6PvNovgBr
45a6VSF+wAK2BIkv8opnKcwnGGzgrKmNd/UcrbcF0fceKDOnhJS06SEySWrY4RgmTLvKFiixfSWB
DhNEs833S78VIASrCRznGOStaW4tkOS2HRWluV/qE0exJ3UWNY/cQu2XBa3MYNwxjauBlGkzUAfj
h8C4qJYvYynA90hR4yUrp0FguUTnhNRKl5Ynbwj2qEXniM9cRZ1rxeitUsIdUtCm1As6z0ntlqR+
gyhIXcm9mrQZ5/hpU8T4RUM1qaZq2i8vd71ynXmdRdl025Equ7zyUJ2uQTH9W9mmHpvFyRd9FNKO
qzpulG6nDW/hlleCc2BHKAqtdo+WkB5N1BOQd+2Ue3YhYkvzRHpxrj0L9yPmrDUmKPtwMkGrFBSW
VNfVdHdTP2hMq+kf7aQRLtFcyjx3a6lqc+06u2R+vYcBAhJ5TTa2WWSIFFQy+UJPTMU4iBPN0QUS
w7wxSYt5yuqhHW2lZTTg7fV207I3TY7oO0Jdzf538NXpPBtZvI8Io+HUtzZBIXdb94clCNQd81RJ
8xrCbYdr169AuI4sg7nTDKXAMHXOSiYW6ERg/kAog5uwbS2OVrYEs61pvmlDnmIq2dyfule18bzW
lqYYUgZ6vuESxjPDEqTgX5sdQ0phH28P8QuAmJRDa4OobE1V/hZVpezKxIdMnbX1Dq+JIPRCbC1g
prfCHs1Dd+RKacHn1cLg17mrED/u1VGJlRqt9R8vsTBKZVItmaQ5SfBBC+ztMezcBEdEu5Wfz1IA
l7bZFjr5DsAhI4RQB9BWvG90V169CBqHSxS/xLZCHSfL6o+Fe/i52qyIX88O80G3ikfS/WRki6iX
NKeeIw+4Q2IwlPpmMwdW89dXusr17RSi6jXae9KNJBYB4lZby2vyLEaXjSikak5Ym4MDdoboplje
i8T9oBeLZL7rSN+l49UGz2ArUkTnUZQ75cHTxw9MOws2xOKG2Jo/hiGYBHY46xPTxPNB3AOtP0RE
HGrm8OK1jIYnhShs5Pl+OvsIV+WngjImWi2r2iEWCcVVYR1Sah0ALVsuaShRjlOpXUQm9Z2ptl5/
Vp9EBlbfXLposF0othUSWUHFo5euCjg/rCwptSUPlpgDBcispqNccCvjT0fnOucIiaxf3ZID31XN
hNnOhcPI8eMK5fiqSgJ1LEE2gBqXAQvVr8/l+9J49HP7PR92Ep28xaWAGC33C70yOKdZ6dtaJDUM
A78gpJ2yYqBAjz2inaqz2vqCuJEqD2UcGxvNTObIM8uAPzQI2ph/IzyYi/39xXDVwCFbC4tCpDf7
BjfvVmJeLl/4EmKF+Xa95cc6v0fIiHAGe0DVS2gWR3a9vT894qT14qQRgO9JhqpDH4QeyB87enDh
gKMn+VAR+blRNmie1db6cEmX0RNAfzqkULLy7NqNKSVj8hJhd03/Jnyo4MzHfRtJ7gWICSsnKnFC
UsuKmbi2nNin42nbWWrMcsl/yNbFUThIWl7mzxYPmzLIc7FKDkT9r0+4yAC3uAg5qin5XjtV4Q6N
ErJwGwoOXC62l4DhkK3P6dnQXRBjJycZxKb7SBW8u35AkXlJJ33guDmAJxZgQMsBR6h5x8eB8hqY
06OTjN6ae2koa3XNcQIEAIMtimFZlaoPbqTBNpAX07me2qpmxlQuw0ChQbfvOGqwUq+62EvmcL6g
PPaNvugE1gpjCCg1W0rns4ahgjByrXQoxxK9Bwmyba9UUDxFoVUGlu3uqh89Uc9QHX4pKEoW5BWj
xh1GUD9/bIvHe3oKWgV4fAGRor/ogbx6y9+yH6uAOf4bbeMHVYnr4yXTVvXT3dTPLH3Mdm0twOPl
Hp4IHHap4JaPlnldtVQT/VMOgHz4SDxuq4ZMQhLM69TCkbnBjHLa6uwD+M+4K/9QavxEO50VbI4z
72cZC2GZzmXiBSWoqgwrHpppSJCSYttY9lvIHZ42wO9KusBD5Ike+baRD0a20w9e63gFK1tbn8rw
JRuoakFpFmptiwegN+yHNb44eXNXMufdTc9TcxDafkNFFOKKTm2XHGb8iwD5CgKgd8RNc24lBB9Z
ngfmbrOHSsQchU7TN5X2PLY+lHiqzW08NVA/wNVLgUuV9MUqdJJiw60Yg5UmQMzkJ8FDcP3U/dXa
yws+KBfllR5RYOc59jK2BPJJgE1KHrKi4q7gf5YUEqlG2ILjFjXQm1qO1ZagDL9iSuMYiUancL5L
IJu+QlDraHEL2ErsdTWWVjN+LxQorPL8Bzj/YfhmfZYu+rdCntgqkia5QW+oS3qVpaqhwvFiEUp9
O2w0T5+r5bEJS+aU26oF7IOYTgCG+X15oC6qWjUzD/yYjkibTCrtqgqDeJW9Tk1CZEJRvp0Fw3i2
ei2Wj6nI1I5c4RbO83KBbOOou3XK4YvG7eXLOtV1yEMgxL8EIdTanQlZ4fF7lr2NydMXzJEYDBe3
FaMHVwfJv2OD6d2FtaEC5HNBdJVHcpAHkNXdA9LnzYIe0OZEWisMHs//9hc9OoVsTVUpHpc42BEl
xGjcIA4ALh7LKa3b/GQfDMZ/0yjWzVoMdiCH5j070821medcfERQS6wF9QhkB3gD6X4EuzupnEFJ
fPKFanBkT+I8PtMrjfWwwzM1vlIw/dfifT9VSKiBbRCJWoNvsTUqjk2kEuoB+V26ZHvmqGacDxT7
fSFWhqe5W1asHucCMU6EcIl2zOxDjlaPsYRL+zU6HTUnk+sJRRjcIIXXGy93maMznLQmoCyue7jV
sP5U/3A/x9iehIISUlUfnt2haaNQ8XWv0G1YXy7GCtRxKO34ZbEz1sCrR4XsXN6NVF1siCrnjWvN
AwvX6+5GyWEOErNa2F3tpb3ovaXoNPx/I0j1/TasDbDLi7WhhFzaesjy9wyQE2iKpLtVMSHku3/2
hsgsOVe18YPeBwXbRmyjdJbRyA48KWtMntdeg99vNfwg6EyuypfE20UINh/BVNZjtynmN9R5MY2Z
MIeGvfFN3m7CxoRSsF+fcveJY0gNIBPzhxLVC0iDqO+6FDJaF7RxUHm8VxTzYSnk2Yf9gmZjArQt
79DXA6PhnEI4+13ynE2c8azv8YpUOaLU5SB0NwWkPFlHWsnq8lyn1Im+7rbqUyxJSkOAhn0AVP6q
GYx3i/XTbRNzh7apn5RJB6CBD/GlA3GXZTOTEPmhsnkTWfu/o8qwvNUod/iQMVVLWBXpvwstXz/V
IbAnXvj2Q66ZbFI11wGMs/q/7K6IjFksAiPOZ6l+zZPzpDzZaACVa1DM8kNTOGM2AVpNOXRNitDx
Mv6/WTXoyoBcryVueJy9/OWjsC6+1FD6Scxnf+V/ECxURzVDl5RKXXYvi6gjlyIh+orwLtOh2amx
34+5ynVJ8NJlHVyd52KzIeA/jsM3ZTrUbms3Z+pDcrc0RzCuDbPlPZ4imZTMbNwjEPH+LPwDMxHL
WEN4+kKzWQCTltH5rzt0GTLsPXVtkhjRfyzKnrrQy5DRJQWweyGLn+dsp30X+BO4jsMk0LEIKkSs
KD4CN7C4u4y5fcOpvLsGfLY9YInnChUuu3Mldt4dZAdwPV9SV5ocb3bkguDU2sKQ3lr/aYP2KU7X
HCodUZdkZY2YRUXQFYDHOwIpCQb829ksvbTCMNU5Rrcw01M2aIrZKK630QOsznQfUQKTMi32hv6T
U2FMJM9ndTkz7EvLyLR6wqiWnLHRIWSi8Tos+BFqTwDXBOG31HKPdh39HYQ3OF5OgePgmYDapnVV
gxYQ1j2CN1NEidvdRwucZdY/toVi9LhvADjfmVE2M/0O/LywHQ1+5hJJBrmGWcEd/7ZGD9xw7vGw
fGAveKiVNi1+a2jLSEdhs/pgJSijbf83fMN/E8a2RiHftXtw2p3KLqXrD/zoFfkSJpuN24N3HABg
QS3riAQz+zathO/KfHCMNADJfSwSd/Bb/e46Os5OSIMnlfIBddAx7PMmkwTCSB1u14AFvF5C+azJ
FoJIkFH0bQyZbDitAP3bauUMqsRK2ZfGhilWuetn3OHu14zpkkkfcYHlw3pfmHuSmnpiu+E1XKve
YlF2kEjEmJpi/Sc18wxhUV2zccBIvWpwaqMcLhFhohJAey81CKH9ZIK43ge3lInyIzwh0xzvlZzO
ysCZlYtTgm3S06vyzVKpswaxlQVRNI/Y+XoWd5T43j/hA2ctPoH1K530IuwB98ysx+yBNlkP1/P6
bGasaVyM1e2akg1BA6hxoyiAw0B0y7SM+nrf/h9J4nl1pKMhN6k/gIUJ0sGu4YPMnKAADx1U4lYt
Zg1W13ZvfyW1pp+++Qq9GFfdaiv5Zv4TfrXWis7SQ9Wp2faLO4tWPHilUGlD9OfuwoDNbp6+VVaC
1O8DYBQ6XGXhSR51kxmtBBMuDjZCx12eN3YqZLtIChgVpWnzY4/3VDxry6lvCxJCY5RiQRHFrJGv
Azqb4Qh+2oA8Hp/ehGFiH7zyEUUgo+tYPhx6D9Y7F/OxUf/y59YcliNXtg8CaiRcUiSD0UBzW2yS
XO/fm560dWBLd8CU8iqrIQmwXUPRvFQludTIt/SYSKwXGgHsk5I/I9lP9mXB+QnjqZMU1ROHz6NT
LFjEBSf6oOaoBXPVRckT6fnaZMxlIk2URQfQjml68ymK/b1qL4spv60jb2vQfGIK0Tdg+vUwHuFJ
88hSA6Ocna7PnZa4p2iV4oZmBxB+Tl2grLSkBbuiyaIPfgaoHfcJG7VQl86XWZ5XkkyEUx7t/Uu/
AddCETYGpkWd9O+4OTZiqqtDksEpyfXWaYmyNLV5WIj74JKFwsyk0lPS7KFQhE5eQOOCKHqmcWpS
XNwjZ+lqSjZdFnJroDL79Vq7j003kgFvdRB/d4+WYs5Dkrmw4ytc3h+jiWkqWxTsBbrFRMdycZN5
8W0hPsS0K5+Hw/RHWtychFYtQTr44KCq4ed6E4fLDuoLs0qK0awztm0vmNKzm3/GsmxZUyHc3FRl
wj0zkVm7oMGllYsI9uAfkX/ldYGeQFKXiA146G8nOCBJ4emisZKuUHIILqWlVTCRd5yhslfJuvEt
naTLi/cPo2riKH/vulLAOjbBPgsfeq1Lu5mdLuj6LIiXjbf3dlgh5aUqSVs5oN3M9xUotGOz4E1v
gMAf5SrPvObPfdjtqtR8rK/wcBNBP5I9zkWUj4OpRP9O26QL4FB+BI/u+B47VghOVD5nh6LvQ0EQ
llzIcwIUBpk+/Mc5yx5zFB1ztRf8pXRLUl6ISuLmiikWD+3VDAsvQmuVjNXxt0RpxUW//z14nTxF
ry6GHfu6lh2J9gPPpBLslWhLLbQcDVjymZgpdkdnphODAa9BxWUmGSoDCZwr1e1qi8QM6OOL/rQh
Kh6EQ9r6wgz+YtPHBx3DCDXQL0pg73TqKr41p/g58c67G+ZPKfkmcfNyVMg32amxiz1Ig84bwVRh
QvYveUdZIcOCkMICUN5uj1ZExrtC7gRzhtaWDaDBOsuoO0a2SqWlBXTXt/5Dg5m6+uwuv4HAY+o5
uoLImzUS2wUym4W7G3t857HSdib+nmHy6QeIAeJhCb1RFQAqnIzKsSPrqV35loGObXfcBGX2bZg2
pRg7jNci5hMuMA7n9oYpPhQJbJvUJNBERxyy3xyMgMzxH2gNsTaeHtT79HWV9qEPndv6qRwb2Onz
2oP0k5KRrLx1NrrIAhG0H+CnqAHcQbrpvCb369Zgt46k9+5LdZYpG6u01rA0agwX59k9VYAqbSqr
zqGX3obn3oxdLrbM64/5O3c1k3GpjGVfYff1Fl5G6XD2JfIJHchtG9KvRn1NO3myYUUExIgdWlyG
M5TFlz8AUkK9/11VFVjpqnm6kA/o4eOZfLeqVBue3Miej7/HJLVxuzXwx4D1rhBxGlC8z/QiwrYE
LZ2wIDwlQc9bUc6ZguTq6u6i4vzuVc2HM2MkJNaH2ZfsowpGmpyAc3a0D4lP37kyHbI2CauuOl+m
QN6dkQ10WHYE4Vo8CKxHdqBLZl0mbFh39whztV9/LM4SRCKz5ySdiHiiEHOK7ZD5SF8zSgzATEQU
Nbpe930gIp/R1kbzHjufytf7keNwTeeEZ1pkHqUNAv+465eW7/dyyrs5D6BiTvngqs/+oAmxTOlj
0S/ElR8NBIsQiCCLGUPWolm6XnjsksM7qAHt8v28sUZgOh6q4GYsGSEiybdeL5zoFDVlV5Emle6U
rVa6nWymRoFzxCQNoadmhgqq1BTmWW6npEjY1D81/PJNs6ov6lZnS2Oeyx3+SJPv923U0KKJ32Xi
ZUmd4LaLb0M/FCgkAKmdF2+DIkEP90F8enUOibuzpUAUAr+8w6DikAGh43S+RcsHl5/4KD7hNHi1
tIYHM/tsl3cZH13/QcLoNS7T1tefKX9mGO3Kc423pe8DpCYdrEGmN8+Rq+KsSxPJDJWQF7w7ToBr
x9mXAnBneTH2wXd0T/CtLMZOrvguyryLj7fTs1X8fdGRhTzcu3s61ieY14w+OqV7V1pkmDryM+S2
zyFRLqDcbPy32+zgmbv1OP0OQS/X7WIllqEZ5DVLG3/4OPiYEMh1FjDwyOR83jde2J2/AyfnECFZ
1Jh/OsonUflzjF/yglsHqKthV8QMm3f2PPaaSKiKKnJc12pu8qmUqr2himqvqpivKmEeR9i4FIlU
fOforcN4314iboGrOCAfS2dNaExo/+bGzugQyS7i5NNlReF6JTqByZE1oKfzFQNdJOvv2YmTlqvW
96d3RW+IzxWm79bq8ZkZLBWALzksnHqWTd5s0HtcuZ2za5+iUU5A+qDMPfBtPBR48/utKqhdEziA
AEng79/zpMZjClNaOIUOWGG/mOLqt9UWa/MVamCr3QCHCoLr05V0qjZaWr4mKDkZLL1cS2oD3mFs
mNXcrT/GXm25PeSHwvGO1wjzRCfsO1ny5G0yD3lLYkttsOoA6DsSyI++iMA0xl5TfOyr4hR7d7b3
ZAio+X3KcfZs+mjeCqlo18ZWPS0/kvzY66q3s3aGcZf07zNIDuTqZl83fyVp0Quw5dQe0ybopume
n2Q1wsOCIC5yknxuRtTEhRlmMnXk3oIKo183WPD71nNGkS19882kBybHtN+jOl7OGxpVXhaayJZF
k60vyXntew8i+XA49OGfwnEPCsA5rdGx9IVMFkHPJdK3OHrvgPxg1ayHXaQwez8pYXmXTk7Jy6e2
DrwiC2jkokbf0C6GuVAY15oCrLVues8zr3XjqF6PXktDjYwxjcB3IMuWUz1mW5OSUmsDapgh6tan
tFzkioUxVc65jTMgK6PvtVAea2D/XydQRdL4yOb3H8DMQVj4AbxzIXb4AFeD0q3B7STJaFQGxNwp
7mjAePnyqqvvn3lnd4Zgbir7DHdxJ22tcN28RdekoloP5Ef6xEicP8/rSxKzXhWo91Ay2n5LOWqV
28PEJbC6DstrCEVvrVL3FKQLsyGjGMNJgNOzVzuNsxnJUuFIxl8JyK+CIBv/Bx8Co7C41pjrirpe
atYvbPH7TA25PVUzEcFVqKIiAwp6zqX7W1p22TQVPim4kBsgyF3rld3rXV/rr9jWEnA3zWE/vQeU
fPnYUGI/LDXHiJBw2hGlhK34zzy8xZRomT69t7s4yrtO5F1yd56C+azAoxr4irJMC2K42kCIHqOM
oyfFTDOFlvHmH1dUlawLlkQI2syUDpiauMA0roSI1iNv1aObO1f974CN18bZAgYUgGW0bXOlPx3g
BrT739qMjAxELs8ZRu0LtO6MtHQnODgkkx55rLyhit3S7BhyuaKvBcrOkHKjzjWfsDV1Fn7kYxbM
t2wIOmus4CBgl6vQUbTRIkz7W0Sm6IxC1Nl4e++sA8WqNwbLJ7DhPjE7tubO+m5Z8W7nJq00cc2M
8llTE+POH/8D4KPtDeW6GXBkFBSoqmpSIPZw3L1M4eexbG8RGcHW4L/GWkE3j8CAq65S9oDFA7ji
LOiEco0g0LkczlI0XrJWPWAPiqoqFRQJ+KdYOqZ5YdyWzNRuqPkLRJLLBCwPLTQFHrxH8H+x/rmK
ynDqUXIbQyHNATMZNJvMh9S8aybdidpXZopPHLUcfz+v9+aPCRxSbOUOuVnhvDH6Vwd5uTqKxcof
4v6JTw77lR7VglJKXa6f/7prAhjkUCtrt3aS+Lbu5P/Rj+ZUbI7qqAHicLOdgPkfN1hjpNjwGRHR
5PqfVbHm7D/8aRWlUDNLReruDsPAO7J6V45eJeW3BNAnQxroWSW2M+SOLLIagemtDSk0dSNdtu8q
3VjDHmdszIksJ5os3Le12DtfPvt74b44v/Vp31J3Tq03ABWEKJV5sB5ztJx4bgnhvaSTgeZ52amR
4VOgj1F+PuYTf7ThgiKKW3WxwWO+EKEFjJoN5/K/2NUMxNvChseC4ONRQE+BnwakQ2a7EOJ8UMrP
2VPKdN0wJ0PsvVdI5PzUAQmNRP/g8I21NJf81IC0WhJrYcGbFdofm8JpDNa6ZbYGVBK5Axmydp4k
5gtC+DyTydCLTNvtVP92U0MqCWHhdAnUlBHkBBYjttTuvGDGUJOpHpo7bRmR1k6amr5kUGmn+L0E
jzWeGYl2H9ArnzLS12SksfWJNpC3R4pSIYnS3zB3yFDl+Vj/F8RElRDafWnXIdGwHFFvyhavVLZ3
jLeSl31ImtmKgyN9PUNQrzcsjhhzoZLXEbjr6Ubegqx0CqJl2QNWGYYYgVpdbXaF7O6wXzr0FVI1
EAlbvxs3kV3ErBNinq3EhYietUCuTxyTMPHH6llWgXqIGvJnRW4r+6BOTDaaADQK5DcCCZF1V+1q
NulvWJ6y8dRzd+2wWaFbqYccu9rLgPLFmtYfISJn5qxC69Is1gIfpgkcKo1cileGr52uQfO3hKMs
K9lLQHmoE5OWqkiPdmZyuFiRGPRY/L1nccCpq2bELgBI7b6t3IYCfkscoaMxDkgUTx7iLvoLr1TB
fgGyhPwrPrGPmVbIdOeWHeLMavMv9dNLmISX4qXesUjbYm0HKcs7yQ9H0ai9nJ6AXxGloWr/PeQK
K9fXa7pO0aX4p6TGeFe90524Z6h8sxq8BzBkShs6G0RQJNpK0OK1CHRY24R7F3M+EGgxt64FsO/O
rP1rrZ4ysaikiUm9Pmgqmu2L+jdKiyanqTxlKNY9ecNfvHSKqh0xOq4cFCcsVPyNsJwqepNcMSIF
pgrRxIXVt6/pksDQDdULLETLUvDeAYiOmdLTrbVwjPrJ4g7rUdUW1LdKeFlES4d5nqF4UUxSAvFv
kXMV/iQdVtJJWTdumdOy39JT7wqbDpLYzrZ3Izdo57idWuboFKxDyQaxdhFbINIkhjX8L3sKbnkr
H3vLPPeaeKetbDtvu2Tw87cf0xJfDDY9w+C+WH1C2qhzd6s6YPEks6JIr3tXBNz3hAcNcrtkKdxP
FQYeToWLBntzo81FOvD/qP0PjAN5WJtEnJyCLQYrOpM28j7pIumsc6wEE5JXN0GYuRQGvCI+q0yy
dD0bzeDpTFpZ6DfxoZ3yLKPYqd21u5VRfWz7RjTZ2GAkbv7prSyCqTXcaRL1/X/VqLdhA004wkp/
Yp2zdw+4lLlFSL0W1BK1yTr81CxrHpoyP8W23jy2fBxbbH2+WWK4qDERRwTSuzdRzEjK0j7uQH1/
PvSDPOqtDJmwhQ9zPTobBoVd8qdIsR6HmYWdaPOhUTbslpXb6UVwUJch6VVMXOs/H1eEHpJUcobP
tnuir7hmNweNh/G2t2X+L8PS5IxunakBpHy+3d8oGUJVLuRfWn3Q12RjxLJUNiFiAvvt1Pc9MzpM
u6Bk1JQlUWoPOrXydeEigBWWaKzN4HChGjHLAvuR1LX8JWCtLuJavh8OvXGVCpPt45K8B3c1XxC7
2+75tOUeqW8AflAjmDELPGlSnRU7l6WmuIHke//0DqcdI9Af1BJVi6AiBhMxYpekwd/K8bsO1x7d
1v54SHsHvmJbCP13b/YSsZDT0oaPRch9s/4n5nBptFbC4k7McxAf5xsUp5RVwHwYEdpNrbE/+SAH
j3FBv6wtx/ImSp4XaCoUFM4Imovze/5cbMsWfChzXveklZtyIHrP5Ga271BoA3iqlOycSzyLKlt+
NuWGDL7MehG4MPk19h9c4YlePa2a7Rz8DasfqoOp8Vci3/+wO5uP2LJzxc6cgfkbBJKVQKgfc0i1
VgVxLMEEvMKIeno7j4q2ulfSv5o1PaikJoFhK4v/L1xmDAqWk9ccCPK2Bj2uHHHa8RRy+L19QUYA
KfL7TwKOR3npd4r3xsoqoqyOvqcNKCVhn9Hf3mjyIVIjaWN8kv1gi12FTOHt+pWzPdv6yDz+Au7h
tCAOUKg3SkITKk22wRNfiQY5TStNot9aGr59arSAPnl4EILNd+eJJq8d0J/pwpPrUnooDyTRTyae
h5fnVspM077wUTJONBcBREBE51p8pdI7P3ht0Cj5pCUcfid0q8DVoUDVsCxvEvuK18fytCH4wHPy
MxIQdwQeAh7+H8peOycnZOh0KZ9tsa9zdS+vmU+nNShy1nogUJ+/VfQ1Joo4rLipXlqrfhEYI14p
MeB1IrJ1syZmNSlYYYunLJ+fr8Ao/gkN4yEW8PXy+oKAghJrK6//g+dPQfa+mgM+123OmzHtv8X9
rz39i0FS3ENwJ/KTI1zdHwjU/mOOzou5nQrHtKFjLF8igcpQ/jeORL/PzZdRUnjwYGRWH63qEtna
fkn7wa0MDudzn80WF+1HGSmYiKmpEe295Xuu4kfvkCB7KtlG1zmHZdi/7qch6HRlYcUlO5XL6MqQ
z9zPxnbBeB1aTJpXOuCzFDBm4c+S54yaVbZyuqTByRkfKMAQEt46u8R1bI3eE5sOONV6lsnXJUeG
HQHtcTo35ODDKWsX5hiq/iSyHUkEVe2OHD8L6Hu3Nq7CI4xY6HTeKjqBllyLlw1wBWpFIWd98EQn
qxWJRIzNUL56ZAzyCVl6ulmVf3xZStDRpH5h/4OCqJreeP+cv6BTOpV1UNh5DhXQweCEJMXg4u+9
/x8g7nbJkAasAf/d3F7N0qnrXw6IBRXujpNyYIT6Z9n8GP1dReTSkERe0DYd9+a52AS5Hfpnwl6s
FKkgVSwHC87JY9fNebraQQf1VZ2wn7ht+n8j4OV5vzZna6FGAAOXUTgf8a4sCiEPsib1Ccj7/JSU
+TO0LFFugd0mQuoLFKgq7xSHRsa/ewAZAsfVxp3U4ny+8cg6DKSmuQIQulBRR/Yld0yFnKAr09Zh
Qz5I7Od8WwUOHPWFTo7oGPVC/M+Fabm9nICBkIMxK7662I4h6LmQWd/07g3I1/PDNjF/QLyenk6K
1pQWII+Uho8PgQ0CW5SWyEFivAh2rVDRulGNtSu5l2VZ5B7BQyd21CO75igrhR6WI7+HA8HFV1eh
xiM+UGxlJ3sQpKNLjzjVxEaEOcs94WuJe7R6wjMWsbVGJRWHDJLV4UsPE0+dusDjm1tRYXnbHw6r
CTSyhgcPvy4MEsocIgRAA1xPGpV0WOzkayQEfAZDdPzpKhfcvh7NjoB8q3hk54G+B66Ei0MKBG40
Ov29WwFTQovwNOmLOZCGz2futf+J8DPmmzcKhO17wyKgSZghoyuwfgJ2MdGM5YO3ymEOuCuF7shq
nEHH5DxcHw2f37JBbHG67cKH3waE7kYWzUNN8EqPeN6s7BDmLFDdGvGrr+figqj9Reu9TrBYA8dC
YNaY1HDv1MI7JJ+3unA8qlUzjPR3UF7RcnjrStUjZoUVRkyX67F4N9OSS2GY6Ir/niNhiRiMEgp3
/Ea46IvkLODAo/AeusI5YTbBA9/lOgtTfPD9sqSctZ9mVfvXwm9Nt3jEWPpjly70E2+30HF0IBM0
lQiuk5EPJAi96hlBI/u6saHsC3heZw04VESFY2b3no9QJTSJRhzJ++CpzeREj6lwMR1RaPRyJ9I/
08Q+Ek64fBntaTGT/QMrB9lZEcjdzvAcEnEERjAx/ueNXS9sRpuAW5JZgG7CwXMuSdLwk13HKPEK
1UyV3c3XBqkfDlIw8a+LWMQSrcygelnnYtdK1tkkMCxZSByfDDmMs9BdkYbPmmVFyM41rosTVmnL
8QMGLikwfMfbhbEOaLodhSJTsRkFiQh9FO1g8QaBWL7+unk32iL4kdJhusbwhnnyjdkHgYg8Iaza
Qm8J1nOos7iFmNIv50iH/11Sndhy+eX5U3OOvsgOx+blBvj6xyW3r90/VV3teGtHDWMOynw2/er8
Hu3Iq20TpO1ueTQRZHpsqo6Nf6FtaQad6J6E736amTnaZabw2jVwmRgc5N64ieXvJx4AmAFKWSVt
LfSPHamkn0eRMxOQkrldoLAUDqZArqqI9v4CyMKBQ6fWbgM8KQJtCxTW5rs0FT02uq8wD1Mq/699
cuDyLrt/xlEyJv4UzkeNApv3wF/dc0IWMqbghv1f6lUchS8RJyP6iJXBrwfXlZrMvy3s1cCeHsBR
5AKcnGn9t/Cju9rc7zIx6a1sbADbXXLPFSRGQ3+qEfkPv+UGU/CdYnzQBQRlmkdqrNJNPdwQcBl8
l2Rvfrs6mUI+sbpgFwrlFuR+PC040NHFiIHmhy/z9GPOwyYjS8h9LmWbXP1sY8TOVg+VpxOz25aM
wgFe2E9LDmXINPr0x7OAgEhkhIDQTjR3LKJmtCS5EV2wI9m8Ng6TJcJLbEm7oWwclDQPFT6HHQ8w
yebVYUDaZUM8c/kKgDw3g0qBdDlawB/seQs1Uxd11VS2vvhbKgwYXtE3qDLnUEqjREs/lBykhE6N
j6FjUqLX5gK9W4FHRcaSTOdVBMz9DNhDbPGZPlPV0mSHLVIPu5JJ4ht+VJQxKKUxx5DRVRTiVWmy
m/9EHVXddswJGP95FkQCl67uGVTxS+Dc0vx/ppeLj3FBRioX64BsfJ9Ard0Dd6iJs/loYFpg3qyk
lQ/vanke5Tpt9cVylvPNAJMthzYODBS0fGS9XlklOhDMvqgW4gjnVLzrL5pjCgkA6c60qvFNYF/6
lNwXwIMIPn1zevDVSS+CBdh+iEg5sIpznzj1QMkoik/aeRjb+7hdVSd2q+ldKNCBqB1apiW7dxqI
3tHFAGfOqXZ3HemUfmsfJDlALMC0W2tJEnKAk6SmT/ES6Q6PMcT6463MCWQroLBC5PnuuEuSRj5z
gkJ8PiNcSE9Q7ySiAGDKl4TwyYWOWYP8YG9YKpV45/XYZbYkbfgdgMNqpZmuCq64iayjeib+fD6o
Ouo7f54M128eE3c7NaoXq5zyDRd83Kn1cwJJymwC4e4uC3nh6VsCg0dZNzRmnIBKS6v3V1DYKpzv
6Kcqu1abb3a+/8bYFdphLILSe9ZSDVk+84xHNCGSPpJtLy/0KJ2AjNjUuNlG4GWl4lJ7GI3w1d3n
eqE+zzslKsqxzGl7vX71O/G8W/74+Bha6qIT/3aIbuvIBqh8rovclPO+pCGEItgeH7JLJb2pjZiI
PyskWyBhahL0qBmD1BMinNExi6GtFxrTa5PK/PlIErdfO8AYjlL3DdEEZT40EeKYznEEX5qf9r21
6p5QOkRLRyua66hnnVsKzXgU5Smd2RgfJp/dBrSVo/5l1Rwk4GLhDp2FXmu7ccQR/vP+spaP+Q4c
mgp6oMq+zbIVl0l1F9yGHpp8jFysUKHVAYflqdUDh2e6qUC4eFkxBS8AHI1sdn8OMBCM8m/3spQm
p8I9gIKc6Tp5NDl+mmdJyWYFQmWsFghqbGMrofOj8h3h3nZxLnmlKYQMSejYQdead8v93k6stIhq
VD1jWyPe6FAG5t24k6f34DgjYhgbjLq1BXi/+ustt9+fh8usjJjboiR4zaO3n342FPrXnn9neCby
PeTvAR0hCFVux9O8vW74JfimTLU2Bkiz8s0kggBI5BfZqxbXT8poUCMDVYCLfR0JzavVYDQtNWdW
lhn7JuQ8M685Ec1lEVxM6YbjBI0efEsWdhyyOnkflaYvMjzGQCuyH+4LMDUD+FQnRZkUCdzByhUT
yqou6dB07iYnSoxOBZXqhhNzjEqYkddmHV2SN51MYU3ip2aBNN10jU0PUjlShcuX1jDjoO8uH3tL
ISYe+Bjk2dHDdtfu/RSB9k/QEiHAraUQbuX008FXs5WYFeZ4IClLqp/bjxfGT0uR4uu4GC49uWsu
sWX4PGfj9K5+bQQ8uVJ3SoY1wOmVCjj0iQtgcFG7+pnxKSIwSZozF3A6XAqLJ6GkEacZNS3jTTLM
rEMZ2xU+zwvWapl9nN55wZv3V15l47Lzjl3ykIcJvcBVfkPSmZMt7iH3XyY0haG3+pPIZvF7ANZD
Pfjo/dqlCTxicmKv2cAkXQii+Vjy6dUiyXgUH9HyS6BEVlTHvfIE232N64wjo9FION1Jb2fjRuBh
DTjGp7FJiWiowws5Z5T4VTiw751QXuB6PkAdqTES8VnM+cVjHdTttlIRccOLNHU1pmFcp8LdFm+4
AYFQcjOzk1slVGOn3cvV2H/oAsU+KLh7R3i0cr6dkhhJAwoCWrf0PMRo2pHSM+nKTPRv/G3QZ6Tl
ogeTX6TL36duQwzWN0TIIeEpfKRYLFvrygJUp0R6O0wevYQFDa58MbOLZbgve36VO7rA7PMygm3Y
tz1TJ0yaZ9TLXDxINUcf9CYvrs4vFimiUso7c9kZuFuG2HNq2yqwhHgG5Pu4t2vcKhwnE1xmqBOW
cPo7eBX9f+0raWiPkGjaIZxkACy+ThC9WEKeWaoPaWyTxksFUuYt12gV2DF7WMQ0oPMXfPP//BJY
FAw11I0U+cT9wY+VJV24Csc/GP3TaxFIT0fd+tgI/v7evDA9l9qmqCWRu363GVXY/6Waw62TNqkC
zVvWgtVznedI2s3FCYlJf0hvbeuOnC6H+raX3OsnbKR+DXCkZIl4/c9Vgn4ALF20ZGvlY1sxIRUK
Vxx5QZdw55PHQh7Uov40iDyl2Ewjo61uE/kXI4ETTuY5UiNKaEVExxVVgUveSlu6WVwKP6fPJoRt
gnqGPL58ZDNTNafzAUoaDeIk/1oBJGL//j+q+5shRF/7VUk9CwwbHE2w7vH0gCwqTY/A4jW+dHdd
B5grz0xLpAfgPP8HYyLKvuiklTFqTS4XadDiKPz1qg/D9Fml3CEJYLXAu6+2shMI81mpnyK+JbkI
VCeDSFD9NfCqmnFfWgVCy1RnA+Pg219oPVogiuMYJPACn4DkexBbM+nUFe6qLdFO3oBSXj6PhZml
A7tPtEhqC4nyHTAerSeTjt8pFvubdRc9jAVkV7xvO9vfA26Npnxqx8MRso/tOG9C8Pzf9FEcljcm
csMNb/oF8bRSqEz3lkesT1wHdYFIifVqtZLJjyWNoiuIuchTSolLJ+UemUMqz9SZ8KLdtjZr0tYd
5edjHwD7Wh2uww7gVbvAg9RTza64fCQ8S6sD5wXL7i0KRqIacVJxDcZWC1YyaHdNHcHn/ccrblSu
ZFwORSL3CBcKopaWq0sD4Yy/rwDdE0UcqZtSZ22+SmL8KU3BsTryJbqSRUiKVsawT0maWM0uDdbd
+qBZwTugedWuD95DtvITtIoLV9aPYiglk7h4vLsAYLNOX5DzjbpfmbXpv4Y4uBM0+eE7VN9pu5iB
WnQHYImxKL1LnUMFG8Ya4KM1Ke4DxSyE3I16nXw/czf0KtgZ7Nwm15EoP9bbeXVHK6ePYBDwrFx9
Gz22JD09/oUv7qg2CBWgogwrS3oPhUfyyiiap/q2uUD6V3yNlE3zXoXpDVKkIcP/jsim+zIim0hG
HNIuiKav2VWIiUedPvIpbq8zZ73YhAxGWA82bQ7B/XpcQk1Ppi3KmMPbadSSrxaIoMejq1sSsUs6
vIvMWOE8ZrSvP4O4ul6I2ekCxa7SaLuyZAe3CttL/b4Bt9jhX94he0w0IDviuDxOHm8ZA6q6DIbX
xxz/yIJe9QWPeBITNjBOpo7KFZW7yqcvTvEdsUatEwsnJPLFqdu2tV6PPBg2wTamI/V0sO+LRCcu
NUxGTPfvF9hBjefmOVx9ITEqNTBuXSUyRAoOI0e0uZSL4agr8ZnrHeHFGESAo7a3Ktk6I7hEYPtU
cNQ/39jQoxsgz7RdZUI0dsVBHtrppmOsdFptJFzP71VXAkKCNu0axgyVbjZXxCGxFRedqvN91jrf
b9JY2E+ju47f0gbCNExckntJXSot6qEB7yMAO/LCvqoN/H1suTuj7maYM5RS9i6ZJm6N5A996i/x
IH/nO+ay3liTUn9W6Xvjs09ByGCORPDGsX1oHd5zbTA5zQHOYgf/nD0hk9rh23Vk+Ftx2RKcZ/XV
zWbkEOy8BseADxV+B1jvpVRbZDLXJyrNUxcWKTeZaIGx3hlEOEiS/Bx4EGRB2z0r59Mb+ATDexfF
z8b9i+J2jMKm4GTVJ/9zbO1X82OQBmlULtBM00A2H2Tr7mRUoES/Dr22MUiWJyfdzI4W+iN/aWBc
axWzBIGUMCRz9CphVo5L86ssB38k1zZtRHa/UP3M/ZCS5tEeBrQ4qVSE0JjfGOt3lVvrvT1Dc8eZ
sgD8a/oI3xlPGcxA2TF9O1UmMyg4/poSpSd+NVISqhdZL4xZKhGalsOkzq49R4OVQBUTPLr91d5c
8M91k/l7o8a5NHUNgJLy6r9jgD7XHNU+HeBEww+ZTAlNBOdnhQ41GSVcJCXFbAHqqkK5TG2xwuZy
e5Hn5AOfyuab1DY7Jt1XcL4Ejcc7BiT5OBOqIR1R3tkwiy0xWGRigRUai3K/P0ZvAdC0KlTTmlEs
ynroBqaHiNGpYSOecPgCsnqHCVASkSmuThDtmweDvGUfF84TYjTuD6VDN3hbB1idXeGKq5A//LmF
EBDmWiKOTOZNPck+0cf76d9yfHMUkxXqH36VIO9rTguPy7nwq0rE4YPdJbxbPKC7CyzhkzV6DTiz
cICDy6xnFLbKgsUPB13zB2jV+sHoCasIBpV53PmrXQ6vQesJgAN3SukLncZNJ/PKp8KaB3ziRs1C
nkSzClHy1dk+SNQULJIAEfCW2YztW28H867YkwnNZ6aUB6gf3jMNnOdbPpFwsWGWeYueLIm0dxcD
o912TtPVC/Lz44+Zt9YbsA23g2k47sMWlle+UuLhdrRPO4zuCYpM/AVoI2yTXMeg9EpQ1xiUbFU6
gDqu0DwyKcbu/fwioPPMob0CLud0DfOVefZCpsNdnywb8WuDQk2HUIZtje+GwKBDiyrFM9lstWxJ
F8No1Ay3LXWZza2TVhb2Njt1fJ8DxKOtREM7gM5mlV8xnOj6igqYBqkRpCLd64XTVSqxb5OXt75x
WBZlJk+EMza0BcO813wyFPfPU72mO2zahUBQgihyaik3VLS5y/S9ub6LN2L+32jcyarFCkoxI8yF
A1H5PJRWTzOHZt607H3QWNHAvAFWT3mz9563yZS0VBORxsGkjDNIipLImjGU/+h88qBeAPk2SzVE
D/UaWbDruY1fV9mDSJXi8hYEwRFTZAuasyRpVZewknwWImY+eFJR0WmP8SOAt0kmJUOjre9cjeKD
2dRhQalShYNOu3kQL/r90nErU2cf7Vs9xv2ejkkk435qgtxlsc5l3d6mNaYb6yY8Vekc0te/UmF0
nXOxLgJfLmPjHzbFX5acPZYKYNKKxf9wrZ5fKAhoWPO04q5Gnh6JGJFXFEh3aLnXz8SY5k5BO1DR
pr0R7rMh5ZbDowgdnL2FnY/AgPgyeu5CsXYiB/blZHSvSb4UdmHghQuQxySeoeek1oT3S4XaSfAv
OV5sse3X/+IMZHhbb+3lI3at/PpYYuWtcDfrBJYdLi3KuNlt+6u9tfMjE+jEs1SdD+E2ZXwS4DQu
nEpsMUkhyysfsvxaJaqZ1n6xNJuplurXBW+rMgi76qsWSoAMrE7BUdeER84SfBIxZMB+h3yZ9Nsa
ucNDnrG3MTq9lSNmuLOVHbEtr7CuwCMCS1sauhm+BgbxYEfVHcqV79InN6Bj+snlA/GskUYG6SpU
CQW0pKVxVFc7hFqpZTLxhWy9aCCVcuOyuwwETjBJupV9lI6OTXia8MC44wuky868Kk2hbjyR6Mrn
G7NIJGx03XrwINwtth/KTr0odeHYTcHTdf/i7KVDqgUbK4jv7cdm/kiNFkh+GuII6h5C51CWGq1y
6ctgGUmy5LiwfJqFN5HbjDcjUDka5km1kHL3sLNMCkJkblac8tTk/8mJhxGydIIfAs/yNYKbvl4J
a/zyk+qM88Rl/Ylvz/mGQ3JGOaq+AYpJvcA8LOeFVTkIy33XranwU0oMG6c9c4+FKpvByFDoeC9s
2qWUP3DoX6Hk2FAuWaIgvimFkIgjToT52WZMd0gk3/pbrQLOHi+8tMkSVU/V4E89LLJVaKj2jBvz
+4u8L3XZs9g8hpYB4ciPJK64XRO1v1uaHYnXcxK0PSddQhY0VFUrw6Ndk4NFDJJqj0CiXj3zwBxp
TuJK1kF+2qSe++QZmPws2pXXRgnfrbmadDx6utzRRdS4Z6xcJ61yuqRBAPDquRlAUbvrn0WQqDIM
mjPJ1Oya+kFawrBjM06E0Z292hbgTxLS7zWBWcxNx0nyiKruO9GBPT/kMTZ3Mva9AMWgauW07GS4
AhwtC5L0TA1j3mj50+be94I0htKNid7vPqdEljXa/zun86IoEhd8gdnrGwTCvupbQUTZIrJxw2EU
9E97Ls3o/sRA8DTcpwU+KRI7nHAgifEj4/Fq2UVP/iCLRToiUrfPVCKVzd4j/dLFmy+e7npB0NEH
eb6a2GxTF/Q/1btXG83GSoINB/sXXglh1cwmr8ZwYxUtajY89VVdFHwWwqlh6QE2hDJz518eakuL
8fc48QcP16wF13+pDZRwEmg1LjAHaef1TzVaRp2DI8duH/bfE7S1N58VbBitY9ez8yFDJNu3sTZ2
ummIl3PLfcdp3yW7s3qgeaxAJS9SBgPwYhczQp/vb2JSTigJ55lUXboILRcT7mgrJVh+qcvTVzxt
ceMwnfYkcJelqMOI0efg4FftusihNYccBsWp99nKLi6slwvcfMBgQ7IL0V2Q1cSLC8QLppmqzkfj
tGgGtTbBvok1PixgznKlHB8+EccQ2khqXTHugl5DaZ1Jvqo2DrR46bdBfeh6H8Lb52Fllj+BAqJD
+PaOC3ogPsyvIkugSmHKo/aWnSLJkRLMEN0jAL5j1eJMZXLLh2lFQNNrVd1Dr/9dvWZ7Th/ZGT5Z
awafDyzIWNi428pRY1UoHY8GU3G+gDb5cOdKLOlNpNbmk/rPRCxR7ol++Gi4Se1aM1ZKE7h1CZW2
FB1DJY8mRXbHQWBA3RAVssyd8y2sQPvqFJYCYuXqx9tUcToBwEfdfcDFSOEJ7B5YXU2seHFtWieV
ZnSiXEuceRHDVM4vEHamvBWNkPGIvSuAIJrxlfbQY05KEkTmSztQFupK8eDa8ZwgAX3HewYR7oPq
PKSayBXVJ4k/UyTwdj/h6IOlvy3Dk6Xd5eCCkYng26M//zvM0FXQMKQNwlYuoY4TATAG6yIVjgz9
K3Tlvt5XeqnrjeActD8W5eS2iAk5bPs+6VNidBdvM4l/DHArEDjlysiyz5PKumV2Mzw1CLGsQ64+
LoI3Pf595BvcKOoPzOv17FbDPa6K88eRvaRZSqEifwH/5FQfgadTwG5VXN09c2/8jLUD4nQwdeC7
kFsWnFNCes3xIpJviiIcqMXHnKs8vdU7Wn8E1rfHL+uZ/bDoXBoI3aCljfL4jXAwOxwRdNE1AZXP
R38oiz01zwXyJyfTEa34jodIIZe+Cw+W6vdfsDMWncwOTJmRFBd+WimCRPNOPGiwf8KjWAg9tsnm
bDLVfUZzqmb0dMVhizg7rPfh7TXUrcigI5bM2Q9lqKAOoaw6u2l5mIlqCW91RHyCiZs6sxuCAH5g
7EiU3cbvIKckf5jlWg0LFX2UaeQGiP7MMMQuCS0YtILLgjhBwbTI0TZjLrLF9vxH/Mq6rTDZZnbZ
9XK4W+p1gtHhWNuAMzgTRQ5jVGpvXxtICUdPOh5VzugzXvdQjlM7iZSTLnpgEhRLa64osypvRDYf
G5hdbxGSfiJa33NRUtCVUUn+oXXrKu2EtdgcRTSHm0q1C17hPeXmhq4ahdnePWqoRU/+6Ywub5lq
qJtwsBN4AKlYmmACEfCS+ETwrpNhS1jcqWxbh+uk8apRptfdOHZcufjsIY8j8yCEFHRmDWkctQj/
iEj8o/9L2L/S6WQnJ671j811ziouqRqc4whHNdRQxpvrwuJbqbpzbNduawPVAlbcUGRdWB9B4sWy
Gh0C7xhCg6jMD8WS4ITcyIz0ngPBufhFelkqKjUihL4ZFpVrYWhMA8lTlqxAHBIgQcYXdLWHHU3X
ZI7QJReAwX/YG1eTKc8KptljuM3ES+fXaHgO64hpOjFF970/v+rfikfOvOy3h0Fn4OEXVbw/p+Pz
C36T4jq0CqWPhISjedxjld4KjC0j5PTpu6uB59p/hvcCzCUb/VrW6TE9dOd8iokECRDEKkoIUcB8
oNYARMmIncmfVtfh2ttWhKqX4LeG3X/+rB+8W0CpZ7sbkGytDI1JripTHHaVHnQGOhwaLDcgC3QA
ZY6A/7GTaVeHB6lxY0tDaezQ1fx4QWrKqqt6z2dZu3AvHK/sjuiYYEENE5INSlFubKGXofn1+3qX
vCbhbLh36G2jivyUWDVNdVt2VrF73oum3rpMx3cAWWsApNO69ehtyccoxS3XLzeKfLWPI5u/fzvg
skZRa23BjYbfLnNQbfFKGZ9udtKquLFJc3lWGYbNpOpe90VMam9eV7ErjIDmxo8+TwkiGLsVnI0T
CvMrhntChQvJyJCgWwLR/viSW+MwL+xm0cZLFfi0vyiq1aJD3nT11mpgzFbtyYroYCF0nopQUx05
ecv3rQH9zYDZD+7hODjU5jWkX0yliovA0thDb3S6WPv/Sp6mlB/WsAn+phdkBTVf4DFKZaU9XgGJ
gVoPpPUOQSe3zxFnI2E3xYOahA3G0sSX+X1x6eAkeDjynsv8teo6ND295bIwGcRdZBhQcXdQ9Zb3
HZ8ywINFIuyYYeNwzfntctC7x+coSo5JwYZgLavfJQOuibFATwmsoWdNy9j5Px7NMBocwBLjNH5N
D77enxsdn9wahyTeDLmaFEHxaT/BJgcX544iaWoaPDUYHpJhp2Azrl/bFuT2pvf6Mm6ZN4MYcz0q
KcFbrgSLvXX+Yn4QH6uUKna5jVkEC22prFWGN8QrE+G3gdNdgvvw64NoiETXnG5NsMlx28qviOlg
jpKnO5Too6dzSpoZoSXD99FKfwRZq8MwpqI+8kkxfyMGq8JUzTLdSuJhpYso37qXEq5B5EbP1qhJ
vyUQOTBxzyMl1GriTncq7yo58Vo3D2W8aM/xhBkiTgEzHaAKr1/ByAy9khD22lyIzDpb0yH6KN8B
eXvUQ/GU4Zlldp2te19osLuNkQ3GP9vSXRhZLKbdacNqii+a7NWdpNLTWma7gQMe9HBAWH4IDomo
OE0+zHEctrbgOFo1Gfb/f/qU+vkXgPEyLQkXqM1zixwiqG5jGRTB5EWgLskvVKbZHteWKYu1FOa/
s1TMvvmGZsSLh6rDgYVyXfDvEVJXjUXG6dOQ6xDfiARhNhQ3MaWP4liVuS90fr0tEGaiQLGwsQUy
1lD5wVf+E5h4k0dJn0UfZpspf4ctb7SzuGC1CkSMvkuI4bl4HmHbTid3gyOoK91Bkw8wSTQLPLWf
x5bpRpdc2x/df/HB38VYFnWDr24D/fbh6P8crpXoLFs/n7KJYnoKrkC0Z2uqOVg1uCo9XJ2tKdms
rEf/U+A6TzA89C0ssW6XytqQxoWFwZolaF4ZAqOo7xbQQqysWs8AVv0YFYEWoP80bZP5CzwoTlAL
4U4vFWvRSaLURRxkdc2iJVM6L2qDipGY3CDWe015WYACWgvPv2ZSs2X39w3vm9yw3V4prHUsaLGU
5HWeqFg3W2T+wG+a/YdqNwVZ5A3P7vBsYW952pTP2tn7RXy3Fiwr1RS68WBMFlP3py1gc+YqTbTZ
JDqCEkl+GsJuK+jNf7np02xajGg/kRkuiMWdSbzkT4koPjfW9pS6brrv9hRNHI/Z+moOdgbaSG/G
vREpEiiYsbx4f7VCoupxxJqiEKw2omwTn46J4JJzhKjbAtUlbSDgT4Nxz8GZ4yDSZWcjP4tf88I2
soq30eJfST3tJn9CBHRiJ1pm3TIXBpgZRrDTbNmPTI+W31jcIhIXoDsNrV3SCQFVyGVMxCM9zIiY
wCdF4A4dFn2YkBYvyt4QO86ToToaWLS9nC//uo1IgAz1RnC8EIZkJppgxHhB4YjJ+zzpidAo2cER
JqLaPZL6eOl737+C7FFJ5cQdLfAYGcFzqA9NVYDSRGmMLALu0eCSVGG7njfKMpRViAVYIiMLdvO7
UyyTbnH39HWl4QWcoc70UjAwArm5OKzweOBzYmgoEApVGGrJ6ZjbtZUkFfYuQyUZFq+RINP8nGOY
LzOgMtVurlZjQHJIMGI1llnEoN28IrPTzSMHFzdglqLqaXGF87IgCxm1HOdp2AaJGQ03689vjd/Q
gjnsl4WRqZ3XP/H9CD54O2be0s8rMzRbQoHw+SLd6GbpWBtPkrou2mQFH+YoMrhIyIkskMijIkCM
3r8zc+EHvcoQMY2frT9XNanKvGLDnAQamtzDZKXXAvtolYMR+e2Gji3IeRWUcxvl+HCgUZSDEwKb
aTX+qKNrtzK9jFa8FX8XGZ78fytKN8Tr3q+xSgVsgDH06QVJ8u37/zCicpzBMCpBn+38i23k88gW
PadDpGpurOGOAv8tQneF4/+ErSaD7UOgXzi4CNCf+2ftXScvSewW/+yAJBFcJdc1KjET3mxTfLF9
O26ojdoPZ2OihenyZWEPwmJIACSWfJzV5+Y4GxOjo/Hv0nOz/JfewHIxJj1Xvcd8haqRC4ByJ2xo
d/25LWr67ZlWMc8KOMFlMz7FXpcQ4gOfDK9JTHuDYoDCFBRg2qCnx4XAq1tJS+iWb6u5+E4bm7fx
oY/55AUU4AzWW/KeaBd/bCcEEDM/7VwOeguTZw6Ino/fkNRJE9ox5LqNcyfDQ3WDZoPWL3C75kjG
TG860YJbb/Ndw25MadpphUJEqMcpb5x7sWbZkXr0o80H/+iytHKoMpYW8alLIgAP4LhmUf8eUJK2
pxkqd9SMkeCaqDPgwIAVDPjIIWj2/7BlK+4xT565Hp6Coi1Nv2km7Wb4TTyJYYDyF/Er3ySIA5BM
oPxt0RwlfeYT8BxDdVM23VjNlOJdWSJXMauETjJqa+UxV7oc9b8TinSVO8Wg7Mh+o2dKNXs7tH8Z
bQhBk8dR6HbuWGe8ZHaDr8YdP7pkuPCZL7yzuLVp0OpbLdC5TwI5gYvC0tJevJ27F91jLJM1rAV9
wbFQhf9U6DoSJSKGrjOsCdHVc1G0DggdfOHI9RCMs2Makqk11jQ+aRUt5borZJsgaoElcMH0OtdU
H0kSZXyXh8CHmJByR9m+WrUT4koC+Tw8Fzm+sKPjWuSPkY5DbTogyBxi6kpRhN2Xul0l4ltpZH7E
Y4RjIA29agSkCebhLVpp2z6YcOEE4e3KUKVvIQzCdTL8cg7yhyvNdjNDP+Blp2lc2HCUMRGkiulL
60ama+KtqnZJyq8eGlR4JfmBT8Uzj2EDPUa1aEstQnXRdyjUPIVL9GqgJD9CFXNRfroJoO2FhT6L
7lt1H7HLIcsE4+zWwFT3BafB7y4yJRYL3Iu0lhp3JePMP246mhKm5ujimXrpRR06cjel6ZskLkhU
G3nk1E8J1xmr96OfeBY3hDQ5ldlLdwpu+829ZvP5aNW4ct40VEbLuBBxeODFLmmWagalBfnBFoGF
gDD/Qcx4fDAzcwKDuSIgpTHQI1eQnDLjVP2AJz8P/Y8ikidkpkIYxh93pMJ0PxpK1tW2XIikdIwJ
/T8L+8UjZM/y/azTghwra8MkXIAs31OztBNr+Ah6FniXh1m4AswmgqlGYeOk8LFK2/VWLD9L+5V4
U/HmdPQ9dEfRzsmrcLafqAP5K8GSkkfcXKYI2qjHLNhCpabVxTSgjpuRsRBexzu0F4aNsQHOn/zU
cr4Yg1P7kMt0mIWK1tSpKxg2fO1KfgxD2ddB7AtSCOnnVtvAytKhURHVci5xhg+RMCZzG530f9j8
XOmACyMK7YOqNuW2z98/AL0agLTRc0dTwFeZvSELKi3k6KJDKP0QjsCC9Eo82bevMvnbUC43uv6/
QT8xnGhgBHyeAbzLYx83HFEHkt/C8V+Av5f5GCaG+ro0Nz3fHr6oXv6seqcaeIGa+V/sAfP9qiaJ
xbkRr/Z/b2SD6Vg+A9+TZaxuGVYhujK9DxQxoYTXly96eHMZsp6Z+fo3PjH4elp0Rr80lOWtz7L6
jzIznsY9hwNv9tVTZAneIBIXo/yOyrqaRYj2eHDzkcGWdsaZvUDxMuvG91v/kzrsfg56w0S5EqEo
jZ2ML4iQgWTt85BjYxnfNiBPZxoYtSz4sQxIVbNO0hePCwHVM2BtkMVeRIzjA9c0kF5tw1Nv/Qe5
z+5hnjel2WdkcfWuiPR8t3foPe6BFdQeViHVyMJUwMnKjm1nDMstMLxSTztDc0iCyZ7HdKl/11Yx
CD7bz91NUH2Z4G5hP/i6McL88kHbF9GkrWC657cZjnCrkgyNZRwfLEpKAJ+Aj7hSLRbzLEyX7ddo
ffe4fOmfL1qIYuXUwLPsP0Ll+Q3wzmqfKno+kblFTYRfyygpyckB0GTYlcqNRyJ4eaTPvoBbGNsY
AQLXHQDdZf0rDUcKYisytJnW029K8MvvGaphxNxbBUW8GPCLiEcQHo1tYMTGi3JnH6vcRxEICg3i
M0X4qB27VPA1ZPABDgUNCY/nA2XDQ1+04u0ht4dmKpXDyH2IqgzzabLozjRqJsUue189oYZ/seeb
yX1KsMfLgaHdI1TW7sIT307XYH5EnkwtER3i63NVythBCxUFy963buplj9EttOrYGRVqZQMJ4+XH
OwRH3kCkLZjmW+4/5THIdxAbLvlUnxsLP1XOKVB+T7vwn7b8ktE3pO/CmWKH5PbYHlI2Ezk3utU7
drSpvtqyFoUS30osRwHlDQ1H+XO9QfDCPU/ylINRNbKp0Goh3pRrZdt87863AtXM/zyCkmNO7vaO
yYuMVizhcAJE1fVBwXOuBrpBUk9fn51Rn3pwDv6IHmtnXKolPc4HVrMLIQHrGTww6eZMP/ST1C6U
4AuBlQyKrKnh0CuBjYyV5yQJlxs0C1CqPfudreFAr0bKsKvU2XzcjAy+Gn9wjcRXnOYnuJAtbwlY
2a6TTe4ciQYGDCI9veCNiQgBKEk6MaIQ1e39GDoxKN+GUJXBDzNbfUSJ1YKIiSj/mZvKGjKNRQYT
a2HBhmvXsBzAJNCvEVnsNTHnQ1ooL7tTen+xRKFL/o9gOGLYOIsQPdGFPlOo1AvswjOHwRIhVf7B
4hzilWwNBUCnWEK4VgM2rqoI0NoKOfW8y4PfJd3oHwa7IEZadoIdVibpKw6twWyXBNa0VW0XrCFq
KVM8ChSMArQuh8hIRC9ZhuVsps3ntt/OPbj6axNmk0qJB5yUbmRs5Td8j2Ql08rJQ5c2mv/m4NJF
2HdIjWpjiixgCsmLtSupQ6Mvhcbx2QfFOlcQIU5Gxa5/LYAj6husZ3YWgPhT/6tVNzljuwR8MBg+
z7h7LPBgkebHkg+w7PalMzq0cdnLa3SS+cL7cvHRAz4j2ut1ozUIAF0Dq51TbLVBkNVcdjf59MSD
sIcSFvqBBQ5vj5/CYjX3jBA+exxXImflTT4eVeOHHMt9t/0lJcmAOyTMxIQ/ES+UEDDaIGTDdPdR
Lpe0YwlJqhhZwpOFeItJeuPSqWXVB2uJZvO7APT5zVnxANEXEo8emHDo0BENSZquDE/Pd7AWxnOJ
8wlnRJ9brYX9MiRVmf2+0whTnCGbSYoPweYFbigG6l8Q97e7krUWLoyCJ5Iu088nIyf0Td8mVPfH
1ML0M6izoFxxrhADxiRqpPxfD+PqvABfa4hR9msjrgv62ipyMhOdR46u6r4PXYnbMYbLASs5CU/1
z/ZxYxTgRPM46hEVyKRGfkWMnXTtE6Gh6I2TnGZ4JmcgHm8HFTksdVasABBjSHYvi2tn2VGuXUyw
zzrYl8YTDC+USU06IIKRjlgNgPKYSrKglUny1KYQq8cSKurbPynEjAaYj9jL26xN/X3e73T1igMJ
UUqGTQrekualtgqfvjIe1ptA23QCKqExn4Sm3IJmbS1mcVXPhycQ+DncN14XL4q/tPkYejuYrurR
hjsTtzZkib9jN0IBBF2hBFBzmW0CIlGU6W0w5n054v5d7qiagIrnC1oEPM7isq+BJZ6r6BFBY/zS
AY2kbQ7g8r+Bce444AIkp5SsZbnO9cd9/fNuRRL0Gsu31LBkAiJlKd2Pk0U7CVkPfSWOnbA4R9v1
hH0zkcwnWc524MmXXyG+7U5N21k1oyEdJPg/Fac/9WRKLBW2Qp9jMA48pKbAUKxEAtwqI4sbKMmx
HsmnGpmB+79N0mSS0Ik1Mf58XIZymI+zHuh9xDOFz0YN5X33UNMg0RmQNCIdin/ACLXK/MKj05Xn
O4leAjYhsnD3qvVWh7YpSvS7Hz8tLYfWPI56Pr2LdXz1S2S0xEVyMgrAwyUjDUby9Y/PxE+ocHVB
Og5ylfQusuEPAcXXYUXHB7V/E3z875upViVbo+jkN2ArbYoLTTb4HTymqcVtBaeExRi+7beGc5D8
ZDBPVI/rQFK5YFRPl85TJz8a+NOAT7j5ok2MSW6itE9E3qfv5YCaDoa5Mq92hrRsukx9h/dAlDAt
53G16tWOsDZr0d1KWiKR2D0X54JA5tVsmQSS53hztOy0guVQ7jHZgsFmaSuk/EO0FEunkTPfJWAZ
DwdqHw2ND83hh0yAVei8UuPenAGrIaxPM10ELmyv0bpvci7x4Z1aHzSspGB2kmwrE79De2AVihTe
qEcXDQv9jHfuahV+RMChflx8F06EJo5ZCuuikaO510LH9NrqpJ8hNF4M43DCwYIRw6fWGL2YKrr5
UxFjMUBOig9Kd3+i3+n8UbO2Lnrjqy3HJ9mmpImf4/mWGn9VbnTy7XMoVjIXIMvQpnzZs7otOChj
bc2xOx1Y0LbJRNZlQIwT711KdtdZNe1pgs90Ae0AlKROQ9y4iMwYoFY5EnniQrkHdeFlF56sAwO3
u8e5kZhifMjeuTKKiJFVyGmikweKlhf0seT72fkmRdDMIcXzO1UQJgHAmiX/ScKAkgUnOSW3DeV+
Jvyrog9cUvdmCm0GXYnAwRSrzCV5vwLXifhyfMl62llM610GfdK33HLdVEINQcpeeU01uGjzOvlp
zMZOfRoPnsyn0xSAhtHk3SGuoFY5IEhLx6OiZFyFM52S8PxG0IUUhZ/Dls/qM0gZ409jd9RA+Mdl
B5PcTdXfRRNzx65UHfHWMSFw2nQGLmtQvra1uFUr1CHffOJOTrzEl6zu7pOHE6w6oc9DGrBx+Ik3
JTl56fLGwGO71feVJl1Eb78tgeSjWREoNuavwXiFejbzdCSF3K1GLo+5xXILcbuvFXAMo+dJvMg+
RwBFuMZmgG3zG5yX6eILqndEFjqrpUj2/n8pMth8ceh34kKJgBPPI9Hyy+F8EpbIwGsn/6thbU/o
+xCz8vg8+YPgaCnNgOtEPkN17BuiKcASOFRZTKXeOVYMTqIJmVpWbvteorBwUczgP2bHQiw3vptn
n+hEkJlHOpItnyHABadXqYZ8Ubyk8MPq8G3wPpIc5Nk5ny35NFxMxlcmjLmcBfxhM4ESXfoKh8vm
AmR9qDSi2H7HhyuZAu5mu7V3/Gfo2eVODZPSL+HON3M/BZip35zjPgFlDuoaG96+8zIry+fAp+kD
wm23cnWFMcbl/P/mH1hM2aVo9JzDg1WimprVd1dQ4Q85A1G3JU3VWEDuIwzREkHXGbxMpHnNKH9m
JsiFk5fFV+FJX20OjYHUyz0AhAsTP0cfnzDUSY4YYOkAnANeeUKJo115qXy88pg0BHlyekdsTJkb
bUM9+Ajhm05mK2z4v6vyjoZV+6sScOPZIn8lc8xqrhTGZzXlbIA/o9BVwKeeOZR/nNCgN7fEcq1Q
V4vEOP8i0uP1zceAxkU6TvEWTTiDAlNgxTlVz3f0DzXwBkzquwx94k8aAo8YNMJtMKP/REIVzBA9
2t17R64faweaU1rVbEjzdPtXb9UamjnViBdQkUrhkW2XHxEcTsktJSlH87nPlXFHl2Pwtwla4J5t
dsHR1FCoG8cGDoTgKMHkUZtnzxacb+WyKcMDOlFwp3n4mkkKOu0SHuag08LQnxQj+GK3IHsKwyy0
rAX+cZIOWeq0g9OvCB9y8UKMttcXXpXnKqUh5nD9UTGLBH/dL8asyNKb7cMUcRXIv0w9P3kuCvf9
ndph3rJjPItd0Uz7hOw4pFNxb8ZAVRKEGG3uLe+w6hsoXI8zTnW/8S9BudtF/C5K33qqYpnMgav5
b8pgAKswjExuYZnqOwQN9HH6w1yz7ipmoEdHKxar5YbZ1ipcR2e0krmlmvEAgY2yCNGCx33ZdA25
6eiUEKmLHBQZX/XvGQ8MLelvVHwfQxuWlbTzfhSBInDEV66YUge8EPDXzMEC0Fz/bOtc8MoiKwct
PTi5F+VAUWMXJae5JKGNTRpWXUxe8Ak03HnidDYmcBqtLHmxChyAeMGfhZTCmU3k+ukMX92RDLXE
YK7xTi3K4zMr8D6C4i5HGo7wY37fK6NbQgO9a5UMVJQDG7ZBJNaAXdli/AufOKxvt7vFBrXhbfyc
wQBVkw2c7iRCAfPH6oR2s90vJJ4fEBX+8jt19rhLNv3o86/hOqitj5NMEgA/CQNtrxnyylg3wbnL
t4DQAwSNqMwJlOboJ/Dz5ZJIfmbfjqATXoiku0F1LPejjgwg/nT89Etw3kjJkWIAiftCeCB9sjP5
E71NX2y9xERZZixzfQo98lT5XlwwDrmQ0406habwF8fF4RpnNCB4H2h8/8HxCLHIpFeXr0HDjA4o
NYPXitwShVpK2n3VLGXqnqbJ/QdFx0w8XbPc0dzr6CQCrYF/LtdEjXKAmmzq/q5sXMESFoa9jMhp
fkb5KtvJzHaEmEs6+lhLrq+J/jrMIK75E9jjzkkCGPShTig8G0FhNStaFEd25xJzU4WocV7Cgnrq
II0aazbgwZPMviXVv5hNfSmka3FwETzZHIJ+udKAaCH7abD+Uqmeg3Us0v817h6pn1OUSN6k/0m0
S6O5DUP3CrEqZEE0likFwl3u0GBIw15WDr6cTk0jFU3RUJper8BU0VLj9+6prjZ2x4AMyes/fV2t
nWx3/8ns9CAnJqMNIxbk+/kIAhB640caHkooqHCKb3opOL02AwwwG9BOEWSj8iWFtxCEFR3HroL/
EvC87qs2ybpZJx9dIZBUXFLjDJy/7s3RWqOqwg2kTcA8Yz7WgD19+V3fivqV2ppLbVCxvTvlOkuq
dIjM2WglIaQiNf3LLWVOGYmJy/e4Rafuzg0HEN3DwSX064Y0QJIoB2ZfI1vqj1EqSUnsSRS7Nq93
EwS1sbww70W+N7Ts2SgKYLTm3VYdtl5hYaukVbTve06O323T7ARS3DqHR1F1WysI4kjNfA+pf10t
oKVW8xXBZirHjXbYAAg4v9NCC69PKZpRrRDzmameAZcRl+L+mqwXkK3AvsoNgQrgD0vrgRMGnSiW
ZDfHG3JUKHbAymrgGi4cXtQ2GJZF4NqJsc/ocCvFnYiZa+wLKQVVDgmcd+grsp2kKlsAPejKVcDG
brNOxwNLymNjsdkevXXN3M9+fQ6Y3AoUc0gnvHC3m1FoGMCKbWjDkl+6oDEzEpTOc01ftatnGWTG
igu0VcdPHMffIxnZMYTGRQVtMEHY7sc2ifKdvo4z6+E0b9eJ2/Vga66j/GoRZSOE0/eMWkVpFbJG
YG9/6utmFtm05mMexSL4shqTEYCuyz2WvYbKVwWJZb71fMwPBMgCcIMOfj0I2BX6zufrcK4BAFdM
zLFT17RW+Pu7VsuDlc3Q/MgpRuR1JPdCiX60+0J8TmGhbZXnBAnfqThiMyNn6mGe1xbEGECNG3Fj
Ylns361KZFkeCjaF1VPc81ZYyZfaG/BZRhRiu6FtBWntvmHeSFhFFkqClOJl3xU16itE4nDxkaOz
c9pG6NlXFr4pwv3To2020cRtwvsHmflh0W3d5XfTbrAvLl50B65jNlMhfC3hhAvWRUwVhg9T6OH+
8lS4ZejfG24aaH8xo9xZulXIQk/viOlOTLc57S+QnOyqFLqmuBr8xmjOafpY3vQeJlE+DSn4UkgK
Nsxjy1+pYSobPKNjR8QJRBqRYG+wO3TG5s7MYi2D9nRNZoPKaWxEpUwytqDGhd/O4flRVTMtzZJl
hIb56O8xmwRqzwXUVolilGRPLG9IRD1hKIzjuuxuyzouUu87arT2VMfoKnu6rqnGNHGgIFrGvNQa
OhcDBG7MXbFGgpIoyG0xXjC5I0ywU++AGVJWLWC4+ACF5ru9p+dU8tJvmtyBr71zj+1V5p4prL9K
9u9AvlHUIB++HR2/AQy+pND0ie1bspEcY87WEPguiHx/zygFLdVbTutgjXzYj0ZS7mJcmzBVjcQM
83Jk+zRGj+Jn9pZg2UlGJbPfQhdjLgrABu0JebpGjZsDodZGzFC6I43iKBqQUsKgOXPzLuuMfDi2
XiWGuxok3wQkWBZrhuMCS8Fw6Wr4J+6atcQ9lw4jp7i1zEHG472SejVbJieiBU1pNdCR0+2WfHa7
9wPRmwxch/RE1zYOfb0+/5eX3x6RQzzcEeL2HfQfOJV89wj9Q+K2eZeLqZa61nmE2OeT74zpYqMc
jsr+vJrvnBJpEJtvcWd18/XCTQJpUEnzudaahUpVz6D8wKlQoLNEukW2P1RyrOt1/r7vEls1agSE
nMRws4YdQBy0DXeeSW9FWkuq5xhPa3ue8vR8Kie+kTdMe5hw6Uc90jJsBW/WORahCDoKIjKC1rG9
WchQs0kUxJA8ndns1MbkCIKm3wsslpnKpSvoxrvNsYJ2VMqy9bkNEraAPLHgq0XqHaWccQiALMWj
atHGdeAPtZ0ksZ0XPxtQrTrjqz1ACr44cb4tm6kC0ZyMFsAF6nin6Ttq6um9LGD7G4daT5+mHw0W
yxN0rkhIT1ENNhSoBC85kix35pEiZR9au1mxb+8gnbjOnnKMOmdLDXhOh/j1n4WqY3RfMriqNIFn
yESgX6RnLG/q11Rdn30jOD/vJU2G0/BPWYXugK+ioCe0o4BXERGLtHca2RiF+Q34EPiwtJGBm3DP
BcsYNVSYGa8r8kSETUaJEAIo8bf15eCbPd2LbfT+QdIjEeM+GlU43bowdNAREn/xiEGpwHkru1Ej
k0QJA75bmS+PmOohoUTmqPR4ZC48rRon48PDWMVt6wJVb2EIZ40zqFdW9wlRBF2a12p5e2lJkFrT
OVt66aDF6uhDt13ucKTboQA4JDht/wVafBfx8FUNmvKyJ5bkw6P4+0DnlPPfkNuRUkSHH31XBnNs
WnSJBfMoQOCUSYMIdSjXkHhmPkQz78MzBF/UcTyiMhmEdAelSkXdLWLVNIZL6y454l1OexgupOcc
tv7okgnIkhtoMf1VM+/BFnM9YbtSzQW8RpTzTGoHahW6oo8ahz/cXqd4CwSmfXDC+SHpXiaFfD8C
KYUl4VSbq/WDuP3ed3ef2YQA1DeXz9G99Q81O49EHasRbK1Jq7q02VJH7345PyJq9Idfotjd973v
h0YrBenHuiAaHDJW5V9QXzTEPHEw8khxcckRfWOFoKNne234EwBzj60HjHWBB194tLnnqEUaMJFq
jJ4eNTPf408K7ot7EhdarPbLhailNVxjQUftYMYgfo8UQrFV/Sl60UXJnjsnJzAiO1JcQevO4Yuv
mCnb7x/fSEjxiTMsYgGqqc+T0X126iPYZ6JgMv+FR1NHpivwwpP9GmxyabbLp681FIjEj4xzg+CO
2OX8H/QjdO0udOZkOeF2VxXt6HCWiR1dHXCrYD0pcUc9AMOCF+eILM1shPZ7+pC24gGQz/D242E5
X6dlpvtoxAjxF9wzGc63RI33og5vZyW5J9akNzVVBriVu/gNOC2MZ9hG45Eds9xtCBwNjh2Zyyfe
3ZgIhLoicUflQ0XyAOshe7ng4de0dmAK7ltNc7ZsQTBjGjTibMwE6XqtpUlhp0bZtRBnU6gXAEfm
o0v0X9NkwYRYPRNAcpIavDnGdNuk5RbxGyPwcG9awvzavTRGH5FO64BKprd/nTqtE5g+z3tOgSOn
VlS8DQ8ftax0IJEXkVGPBTFUxeA3TYwrLkdWaI4YJ9+vCFKEqhBMzlIE0pq9g3uAlO+KN4AxAnfD
BqtTu1zModjG702HWFtONFmx8W2xGWd4EUsyDSDgSaGU3IMWOZWeOflXoN2DQpr5gaD6j4Uc3R8Q
0r9ehOIFo7wK3DCm/0mLuyfuXR+uCjGvzSiBy12TtBsskwtMXT1hPmyZHhHlm/gWECQ3A4eR80cR
tUt56HNcacYm5B2K8IW5DBYg8qNmUX3pQUi5a08B+Y6m/gZIyv0JePkTK5i27GivKKdJrGoI27nY
bQ+5R5dhjjrX+yYzOMW+DMsNFJAVwNlZmRrpx7vKzX/YnLmh9Kbwj9ppgnGPvLlPlYu1JkDeSzGN
/oAYpj9vKpV4bmT2yYvz5+3LUkYn/KBeR4r7T2rOlJBidx2TnbpAGbJvxz8UhJdqu+Q39m9V6TLr
NvJsq6Ag+ef2zrDBMsiv6V02YYqvRX9pjDlpL1lmsM3h0yvCNn4Dz5ac/JcXfrweSxenWOCY5kk2
pso4//5bYwo4OBRaTrTpWIr6TTe1Ckkxwa0Y14qu84kHWJXdYr5cQiaDS+86TNsctQXqbCdg2y3S
c6C0weBAmpmo9BNTnmVLklZr70L3TK2YATOKXWVs8LI/2nMah0MNJ7E8C1oiUcbI9/Q1ps8GhdWY
fgHf2mWcLoZACIwLI+xZStv3+apJj0BNZs46mUtmqy3YEfnwu2AhqyQzh8YbVWyBHtgVV9HnCp/F
8gAtf7a8Hsd9hdzKa+MejAFAWPQoTTnxFUC5KfotD6aBGkEh+YnjVjQZLXZnj7JSKMNMJ/LdxXFZ
C2VXyWFTnT4U2bUWpP7Gx+A8k9+M2qmkiOGJ/iRFQju8p1HnoX7LfHk2sQ9gdmsvD6gCmSmoumd6
Cn9/AX5JAzQtgn8bfgbbSpy8PJS5INJGFZzQetS+O8/AdZAHDrbUs+cYi5nK84gib/369RAu843Z
bLjte4fHcQeF3vmdBfFggUhqmks9L3oBIxPHH8GWRw4jifKAvCvql+HjFZnZ1hY1hen1H4Y19Sp2
hGz2emScY87HWGflI/xq1x2r2P5TR49nOepv6xlpLQfqrZPLsnT2xyl4AFlStWykdOtZwA4mSCjP
ryn6iqJJF63jr+kCI3LyyVdh153tDNsfKW9tuu13RaaYPCrahU9o0qChVMDpRhnTXUCnk40NJ6YO
6PwoAPGI7sJYGmiFQYdQKK53UAE5473cYDDlgAtGtIQfS+EOtZw0v0bI2uINUsRndenZxK8Psu4Q
G4RwmHpYxxd2DxP0yOCuKc+NlzQMFzyVFCoibPMUqB544QcXRBpACiqKlE5AlZFoVEuOtKfEKVm4
mGgIcpb/7xVIIHFeeLhBZe6VXB4Is4UOK8j1YZBxPnkP5wUgjKTPI3QDVr2UuLGd5EgvYD22kJbC
daU9191K9ep7FgW0tzyYpsGzMWCSSqS2+DSdUPGuq/cR2qaEl3IdbMk0NxDi0lRSCAM6Hx2xXUKp
o88uHN3chWGV7SLOdPvw9lDCv4TIrcA+wSRh8OQlAow/5jjfYEw82EEBnoK5BR0uTqt17z6YFph4
RgHI2MGYP2Muvvq39dWkQxiw0CUyMZBLSCBwHSbXmRMUcbEDI+WDMIyb5+J3qyQz0gJpYR+7tSJ/
MM3hWi+mkINudfrSe/3u3ajiQaty54JUFL2TRGxKapW6Z2gNUfvz3ZPbmiEnbmV8J9XHk0NLJgKA
1GbZgKFzFQBhd/ucubvm8c/ofhXbcWSpZk9Cd1G4yqoQ6ZTJMsj2P7KBgoyAtnzopxTAbzcZTfmh
wtT3GyJmXzIyrFhRpfy2FuEuhogJ8fWYHJHnOboHiCBtBOsJEczDaMeVOhB1p7NlTT1sXlptjv11
oz5gN7kWvUipLqUf365WYdGQHh5iYmX4LIxkMG4oOAOP0VQiNuMWpboYG89aSFLRKeNwWw9kCxNi
8KpMFOxJ8VCMTH0dOmhlm6apN1Gf3UXXqUX2lfVVg6a5VFLcnK49/anlli3+4PCDHkBz9i73Y6f4
qVoThnkiQLENlJPjqmqZsujExnLRj34qvutjgz+AhwCK1xuUkmpVVHy8O8YCEvcy/l5jICoxDjIt
UhIs3KWbW+jfVkdBECgdMrN78owC+um3xgbDBltMou9wc2g3+/+SXpEYZbtsQ+9oMuWo4kewS+7e
t0HFkY+VQffwP0nje96+/Ck1Z+TedX1HKsrgiIStkdjRLttkqqoXXRUXQmcIXl7/4/Q/bg47/28i
CeVZEMPFqRopNOEV+fAYmIH/tFHUNJCdxIuOvOlFKSTrKgqzHJEXeqQtUhLyed0F3zeTNAyynHRq
Mib/p2mX6qtxhi495O97rb6w/V0DxCiXXlXQoEKeEGFMnPHI1Rt30Tl453T0g52m7LpDo0eXrFqV
59bAhxnqkajb5wilaDNEAA9RgUl6gF6JHNzu20hThTBtORYCX9Fu8ZXob79s0ATEepItpU5jTNzg
QCai6PmuCWs65vKnYJZA4lD10Iyi1Uz5zV6Ha2pApS58PXZB/8EvbzYcv66PKZ1eWcR8b7WywCeJ
FsmPgc2fO/PGr1sf/Lw2qMFPsxWEGg/+sFV++UeSKNV2VoOoqZGjrlaw4FypHvguSy0wpy3nfPx3
7xa/zADmwkLXYBv7zo7MxTbHiKMW8wy72HRknnouKJouJ+dxo+w+JqjzxupUiztnDl3ovMCEOL0o
bVZPaJgGuPPKb9CYLVRkFXrLbAfQO4/GCsFVuHtd0ApGAcOSIi9DbKcgsSHhnvYTGN88gK5nxCx9
9lg4dgpDalf1oJKDs6Px/YHVFfA8+so9itMYcvlABOWsoVca+4qeMbz2KgdyUyAQyz99c2oKH5c/
9DcJFlDKXLyPf1vrUG0t3AMCWdb/SUvEuFioXxoun8RAw7l+lQInugqH8vulVp5XYacz4u2vPEZf
BnnJgZuQ0PR3oonJQ0VvpZTiFCXEgu60CbwIWoZ+bURADUnUpHT+cekzQB9oC8CUTaCktKqBDkoS
u5Vnx/TAYY1jrE/SOjxXiD8iwuy4SL1Ko7TDlWpEdemJJf/L/myijKdLiCDaiwDEJoQX94pqgOls
gd1DknTbjI3132Q0UJL0BdnTEptbZxBtNAFieAVqbWX3OJF1TYRJ9bA4yJ9eO4jJKICMR6Lv+zSa
uA8zmjKqU87I7mP8FJwucISvyy45VQhYEg6GYpbSbFxebrBM3kYKBtN+y0/GDeZGXBU3GAWpD6qQ
o2XQ5ZPwq5QhdLJdryqJW6akYJADLCqKq5jqjgVUHc/OVMhmbeAozQIV67ji2ZInMKticl1o41IV
uAbm76fQwm35R49hzkzytvPapI6AQoC6Tviq4Xxqn38M2n9jl9CSr82EPzljjWxmSPpgDACWUfZo
i/NFcK1aAeTMacu3MEMm9k6rfNKw1XOWylYgod8yAclIkjnTWb9P8bI6CpNACth7sn+cWBKgNMXA
cbQ8Z+ql+dDaXMLaE7caLPx8Ik6INHGn6uu/jIkPOpRLc2pVJ52TCa1DBlEtc8Ft2I+lY98LH6UL
dxNOu98mCXnPmtRBLJjRvHYQlcpEZ8SEGSYKwoLyuC6uidUaQA4V5NY0SJ2fOVRBc9IHTpPHT90K
E3pYpcv+o/ZqFs8zakpBAgXzZE2dKajUPzFLUaS6gFDmOHvzbAV9tQNH/yybBSjtDpQfiIY+DMCi
0ykIlQEthbf6hrpbzqbHKRJDUz150+SkXzMl91Oy10naL5gFBRRBwZKZGSjCFouaG1UPIyLEdLd5
47J+sahAy2iQXyIGeUyZ2RW9xHtYyJA74vwashnf8l1ZVBUNL/t3/ERF6Osn72g+m7VxpPFsNyIt
Fn8iQIvZga9vo/XPE1ZDW0YmHo8NMsETWy8TuD2MqEYF76unhxTb6jDtX2urxgMMTKg/ShgSU8jK
Fv4+vN5vSkLpE/7SekWTbSLZpDZeGGadUv9Or9PUeAacyWlubcQ3YDgxs5QdkmGbCHj6CqnwkQPU
oaeYJLi843g7LwSFLpcQnXdiBsx0ir6mq2N97oFfbevZ4LRqOUkSW9tgr6Zznrc7cG3mK74tlgAM
aNdqwBp7Qx6Wwk5yyW+0Hcm70MzFtflDgNAJQJNbwhYjV1evK0mh6GUaEa/QnSuYoQqshZ0FHFKL
ZYLDleInuB3yrxVmdDEGGzgpshPU4q7vJQQNPdkr42v4iDKRP2krSuMMyxqIM7qT2Urc+JBZ5eV8
xHqL1XpMEZtKWBVI8CvrcV4EVCGZRgU+S65pPXk8fgVPbZaSRknYqp38N4Sb5zKTpxTOl219ukpL
KwDMAau6azD1tlgH2ghKmid0uL3/LnLj9WUdi1NrFR/EhNiDPakOEjvA2LcrcmvPlUmPOfi3CSF/
lFERT+Rg5MVNSk4NxhMoThFz/z9ufSvCyOQ7eU6qp4LINK30MIANRE4VaI0wg7owbyHGyMUuweZF
q7jCft3uHw8rMvQpTx8qwQ/3FQEpRKC+qbDf1c55jh966t8ObKBZ2UWZF8MYUuZbQMtST850xFjG
Zl1DBVwHDm/9DUpDa5WLGmNBtyZK2FJwkoZs6a2MbLOHp+Hd+lonh6J512poZ/vt+nSdKi/zYKCh
FRDTnQwJGXmTDKwby2nCG35zjcLJ0ICAAHjP411B2veGuFFxnxFtRPUhYmgpYBe1hIxG69R/y2rx
F1/H0ENEoN04yUwYtSnrLxD75D00HYDWei0EXlFk4uVAMY1xTUj9GY+e/qu0Dq5HHyupevlNwNGp
SDVFcLRofv8Gxn8trIWCopZEuuaiGuSFIPmUZRkadhT+PqNjt04ad6LN7OPVm2WxpaBST5UGxu/+
kfMRIS/exI4aJ4gEf+g0W5VdDOF4zVx2R+nYlm587k9aa8EgrqpjOe2jnnmbODhmDCOsbt72pjjD
YT2KzlIoH50oMy2IFs9WbXYr2wzFMvfPBslkCqs7jN2zHEVU4w9bQJhsSv+4nexosNgbQwvATQLj
c9hMg97/YdwLtJ54tf/iPI4UxjBZLaaRj7qkXtWWYHZ/e4PRP9kyQtHZ1m88Wf7EpFxki09/MUBr
JPKz/+M27s+YukkeK9/ktHcwnLv0hrFsfkqEJtqgyDxp7llSsuA6X5fVk3y6iL8E+7Rbz0TNMnQ5
cUy67OY20p1WmVh9hpU6wOWLbIgu8qR3CV216KBJOZ/TbVPMjeVDTluafJrjeKaunT2bESOuBfuW
7leLMEGzE38gQZl4NIbx2HOq9rShGNxKwiNz2T0dLPeFBPP32YQUNpSBVEYS+gQoPiACxuYT56uy
NoIggrl1dV1uW1MTHObGuFtiH5SBka8hEhk5snG9RGLaLhHZYrUpUjbD3KvAnwiFua5JusE9+sd5
sRS9HsAtVjgabNdoZI039FY3Kutu/P5yxg2Um+whJcHcbEYj6jqFFfSLtKneS1HrrC8XIGPl89h+
6Itp6cBuvmqbUscXW4xfqlhVtv/77mqBKIdFt5OAW6vAK68SdpmZJHmnyUXumlVBhZ8yGrxsYlfG
o1MgIjDP/f8rshcGM4k9DUoby7Fk1NGF/zYX31/s5QNPree0+vE1GbzTlC9lIXHufGYV881GiPHO
hZSTegcX1MvFkwNsgbpyiMrkxafdQHxV1QCFeBzdU/EN4tRte7/B6kROEuqMI1CNS6TO8UPjZ7Wj
SNYLJsv7bRJJa3PLS3PQfNTS4O/cf5evgIZ496fLjyMkaGHd88xpbgPLvsAHRyLKATH5uHT7t925
JGU6+lwdzMx3mNhugHV+FUfQ7PkLtTnhibCZhekiUi5+d13Rtkwl2Vyebceus3/foi99ZU/++V3I
HQFO+zCIiU0Mm8LwDZamFExUfYlbgiJUHdiS9P7VicINNeaw7AZ1puaAvK2Km/KwPK6eIUPORJ2k
tAN2L288U5a39BW9BEh865kNZovP0iOk8jIQMmgV3iYHdVxfmKGh6LqP6cukkTEy0TC1sfhYCCD6
z2ZaNwszNKVxS9hwfe6LyIfoGf9odSs6axnKqw2NBU3i9JbTKGEyUG4SyLtdVLpeU3HKYbQ8Lfj9
17D0VsTMDRu2yj8Mxp7ImLl+DI4dvUYfeektswsAwtvFED81gzRJRq/pgl7rVD2oZF9NCyFOUNy9
jmq9KSi0zPyjmR0OI4QAqog0cXwN2Dp0C3fVoeoc0pCGdasPKMAX91jkwZl+IfMIMwaRxbRdrPIk
UjQ4YKNfbvs2a03CRidw2KGsmXcDwh/y/OX/ipHr/l7v2aTSb6qUiMZ1dPDA2uNFSz5IZRHEJ7u8
jqw6ADjlkAoU9QUZH/OzUZFfDiwUkGDVnl2VdeAfKVUox0MYIhZWgOSXw5Q3tppcW8HH0wRcDGvi
1h/M/KXF8qhYUjjuZJu24qxuhb5WopcVP6HQ1ynKc7IDP+RbIanYAcu7brATeX1rWt9qOe2fVMIO
WfUJRDFVQkRacWS0YM9z1uCbGZpCq/xxMZXynHfG6cKxsG7K+xLWOCmcIWSprQ5KD8eO7u3cn5FM
SxrBMm+zMzHEtuasv9aXeU2aW8b2Q1jnHIhkxL3a9v64ZzaFXum264PEdUdnmzTCt6mBid09N/Xj
Ojw+SBNM6N/sRdCYQf/LDbMC7Wkyeush1HfrbvIxMopsFCv7B4wF37J/q8/8XIxZe8uPe1bVNY7s
E4E1IFY2NFutXWqc3i3leH4X/gwxoJVP7psaExk/7K9eINp13ZludrGgravPTYsbXEBOQwsdTdrw
KhZl6nwyq2/hOt51d70V/sYMgmyonX28RcKFnx11c3i2H2F1QHBVae7tAi28gj+bPBYslael4lNI
Gs5yaEbS2TI6/Pw2juCBirFObjw5h5C5v7dZPVMPojqJcJ7AWF6Ycikz4QE0Q8wktMyEYt4IG7EI
9KUuPwrrT+lntUEFH6RJlPyls5WsR5eunai1mEc9Jtv+Xv/ZyvvViyxUayV2jgeE4BSVM59EMKcE
TbPTWLGuAL80ersmNkgTNreAWG9+XsUwPBqc2uA5yuO92vBezzXVF5S7wKOZhmh+I3/Z7IE3U7fe
OiqbE/2ZVlgrx6h/216oSfUGC16RzueQny9zjpU0K3ZusoO5F/a0gu0lrQQ4ArnWqe8ncoZQdAfO
vuwc5YsqxMi4w7eNViM5D1S2SBDY38Gwq2rwxZ8sNGMW0Q3AftA5ZaeDX4vcgop3cIRsKoNsghOa
7Yg7pZxzDcfu7DUiSzPxUBzGjkdvev4ZEUZNq4Kpol4jvjP/mUfI8nq81ag/iZcvfQoIzrp1QgWl
n4enEmnM+4+GnCbQE+KfmD0Gc67ER81wD7h6WuvUhuVFKhdjnqZmNKM1onWgmqmW3SIJw/5Hfg76
GwAcB8AQF+nTJ9XDFvVW+gNvmZVX//Z1X4CGEg64+32hdj0rttouwGUbRwIa0yl+IV3OOKVft1+l
xbCwhwmZbh06o/6sYeYSSlPj+HAwpTvKKKZ0oxZkWaOFZG+hRnIwPdN63nH+sQXmIJPHIE5er5ya
UFhrApr/RWNhmcMuQtTufD6Y4Ub8FwmC9ipQezNNyhjDAW/AKJrD+IJPrempP3cKGVF5RtULFJLp
9ksXtuU8n0158U/sAz8aX3CVzV8ZrCjfQbsWcidLsAoBA7PyO5f2Dqe9wWhTX+DS9qARayNc60+4
d3/fL4rg3SvCsZeWFpcJjMxTpIeqLhkK3DwldoQa4tma/jGtnwpGiocAfOcXnTS2w7nvj3N5J36y
C9WgGFOoVGfUUtpyLmZBfYxxNAOL2blK9+95jiVe5SIXbctviWgh8vk823Bnrvb0YYK9whv+i+T9
ZKU53bKG63Tq+8jsSqgETvnpzwAlx9zkIdadLi49r/ZblANuy0zl8kcJL3kW/pgXhkCHKCdxfPKU
J4Fj0ovO2DCbNcVuGreI0otAr6bqKKNOzUbcbxYfWACKM8Ri6j1sSqvIF0KIwVbVAiGvxVhx/VbL
6woYHn3r5/8ZsVG4+rifH9kDjNthZ8I3lf9C7Y4huYzAvuma7duHciawWHF+T90JcgbZgw5HMEbI
dmffWv+HhpjI+ncdXUfReGPS7Si0SfkfPURlb5HGDc/b1G4O4IfGwsi7lEmZ92X6lYXQv5FvGVRw
utoMFGNQQ/wb2tK/j180485PO0xxtDrx25cwqBS+tArFIfg9hP20ofptCCbBkiVRYQ6U4BoOHRMr
TsWvxFxoj1DB3h12ahJMx105sM1mrYXj9AYK8CsazdUJMnzMhfQcQggrxyGEIQ7j4d/fnd4SMZv/
vSnSqwf9bmj9CeFnXScWCmTBl2vNfHDgRuVVfkGUuVV5DOXsvXyZVt0c/SVVpVkpWRLdA+5hf4wV
NAT1Yt4PcSerBs7SuVLV8PZqrmQokwnjKnYUF1ybT9HE5Nj+rfCBPu61cYXLG2hgvcckItdsfs1M
ShATl/1jk/4pAFPjH+pwRSO04Qh/H+/Goqa2uy8NZYswpUCCyNRVoM3+zf1drnBsQjkC7nAiMYQp
QQmAS13oD4mJvpZBShacGa2EYhmMN7onHz0bflt2Z8SkyC4reIehc6HV0g06t36SuiECVo4gRL3s
GU54kYMFCZFvrru2v0Z+3Man8wFfsyEhCPhccG5B+Kv+sZvllP0+KeFmt9dI3qnFTHFDmrSsAueH
iSE5FWDipeWNBBWTKRBBCuSIbPf2Wzif5LoB6KaCP+42HwCgqOJv98wD/A/Zc0F5ZI06VIqkwADl
qBQIQw8WxUD+NToRcrkPd9HZsYs6cg35c0+9Nr6RQhO3YE/2Ds+5otjvmNGK6Ab8HO0rjKpyYXSY
gEhRdM2CoynE7neK33PzEKtY6JJfMH8zPcET7YvvQpDfk/ihGuxf4qF7KY0+GAa1KIa5vrfG1QvZ
XbezEGQCddKMm3JZrgcD0nWVh+8EEPo4KTDwUPafD8dnTDD85yJh0vpnkujh9y/s5jKbBZa/OWha
fWgnIdYNRPNTYJBOpLt/QNoNPdRob5w+H3H5r+egj9L4aOVEuhTITpmvYbgzpzFeBXvCBVhJn5jv
Z6IJ8/mPHMj4t28z96/tXZ5zaxllUFuaeggNnFlkN4yyqYF5L4ttHZcAO2f/lHYOs5mK0Kk0c6RG
QVeezzUmFr/ZapbWPhist6kDDLQ+QML2ZcNXPw/IcKrWxf3o4OY/R1RFfc16ci6b4A63x+F3K1Zd
Cn7CT9krMy+sdUxx8Ccgv7hRolEVGdr57uTmQA26JZtOI3OvyDAMW70B5k2NbYBvC3/mlfmXJLQF
RHI7YeVu+PjK1gKeU+901tZMBShTK1BKk5ygBWIMjErXxPwALxbShv+czXjQEr3ZcZKLlJynO+AC
hAxXJubbOPrpYslz6ToP6iVypWZ0P1LvvZFIbr1RpGect/q8EBbvpJrWUljXe4rzrSb2tQ+SWtDd
eBj20FAycd5CX8tecsNRDZQMB6SA5dCAsjIgvkiqaHBEmOJO+/B4fJbuqBCb7xN65K4AWRz05TyL
AYRg93rC4xvuZMGWpa/Nsg9FV32aVdZq2ifAmrRFK8dnqZbe0cS8H8qp1KOB20q8UW5Nj2MkmNBF
EV/kGh4IwKVaI7DvkP0RxQZOJsc8whDE/Kpp+CieBZ9cEVtT35JB+NtkLCW+aU7u3TuNaOcv9vKR
DpLIZF/tVIa5h/OU9u0WWJx7jxxxweMGETaYzIWK5ACNaAYQBf0ocZlZj97lrbEXTiESm1I6+urf
YHhncp8DvZjcdqf+yjIlYE6UuOUNSoql7NZl909Ui2k3GxB2kDAwdHmBp2dbv1Sn/+c9EXlnu9te
KMfT8KeSNh7YJehZIV+DtKJrbB1p0wb2rqUB2ib/OIc48YPDzWZnUFKFFJ680kv/ODTPbo3VRP/l
2U63gHpzjPAvFU9gh1LWLVkzO/FPxrcCcut5Jp474CyFuLFn3A8SRcl/KWmyGvRTJCttFEaXZyGs
sAuVtLBNaxE5DjmUr6k6oH91FY5HMR0kh5fnOEQYiGYta2za4e5j9Uq00aQjpyWbT5GZ6PX+aZsZ
bEM54ymObmlgBF0jgrAWJjddX6+OFxxJ0opn0KgUG1IRG+4Bugp84foIX8RbaHwLnLXWUtMoIfp/
z/xl73A0CxrFPsAIgJfQCiZEGUA9mAZ1CQybkNCbjXfgRWqH3p1/AZk7ybStcXGd6f6rLEBXJSMR
1MI7DeFrzmPfWG/JgWHKnBVLwAjpn8fSEMDfYHD8tmEHWSgg/jVvZYwsNLmJ2EH6vt4wIs/oAcQv
nUGtJAImsf4xD2JGnqcr/3OPqi3xb+brlzTyx5hS1XqEnMTI9BH75NLYkBeNC3KcfkR3vi66fDGh
7so7baYq4yWyaIbvkfhTeDA47W+PgjnA+dZUeeHW4gbMcalJSQ7wwyb17+hX2jQgLVbzRVe0O/Mq
A8wGRjhIFFoLDxgYcojIWq2gxy6BMKLyctRHZYtyDuE+HhcaFDDIFBH2ebLaW4+s4oczC4Rnnnsm
WyymcXxndiLi2DiApaaWiTNajmyQsdQUFOYpFgHtNTyn0oOo9+fPNDeBKBxbVnUN2+yrriaDYD74
UGRZPnT00zskAAhM0fM7+HTaz1FrkBqb1Js2QPLOrpw/q0HE6uLhYrSVBC3wkQHgWBb9HkZo5Cw7
eTZGcyzkTz6vl0JwsQdqXJ7AqZcfMceMCvRRrBNM1gSJBmQf8fu6lyKrycd2bFQ67CQjH2/yWeJ3
HFq6oGZEvl0qMMEt2qGaovLC0C1fuKdnKqtOiE8rcZb814DDPRlLkOty4Dafki8EzLYzeM6PZjn2
I2Z8JzLqkc8kgGEnrZMeM3taxfeQGzJl3AW8EFmZ18hCpdEciI5sOkYk1lACLc0zTarLjuc6r4nq
cWM0WZN0KggZAHrC2QWepF4JftL4GTVSVnIJutBI6O1Pf/MXwNI9s6ZXESJs/IfbSIX+huLwnljk
HD+hdQY+bvBHGtDrvIWD+29CZVa2D8R/GeLkOmlZAmxSnmUvq7SbpXGJJyAt0W6jQpnSM0S0r/8b
tlJbFcw9RLwtQvAv/TKZkOdPVU5Q1msWvVDMcmI4iaRi7sun+tVt1BdsWs0+ZWg76MWFP5IwP/Nd
aQyUGbTiVrDJgomcb7ykuV3vxDFwdo10KgUd+tk/aXcfZh/+7n3ZI2msEyg8gS5UX1mRhe5+bT1V
evVzW/EjHootuUdaAQENZOuSKm1n+L041jJJ6BUu0EyAyfY9ALAR7NVldZrOdJtMf0t/YoN7b9zk
7W+aVS2dQNH/Y6G/DZfGkEkJiu4q5nFyTeAO0gdT929ipFKTFI6tccxJmsKKMKKqmItFvt82r5mf
scF1BPhkDYr/rrUO/GCqFqyXPt2Rba5py4ifBR3sgrdoeYzrX0rMZv/gJe/O/RdsmyoP05nrdrV+
TpGS0cdistqwoUqivkmRhKsDiomowpNv65DZMwSz2E5RgLKIb2xa86xJGF6Ha3iuFXrA1XzM1q27
fZNV5YEcTUimJcWv5AcIbfmV+cVWMwRNnXIlXVO59vB02smKe/D+PrYGEYxuige1Nn7nK7EiAM7J
pv5JJcEHhDx3wuJWYlYCKDai1S9U8cZ6bxH3e/8QzO70amMKIm+2E+bPiUkw6dcaI57hdgV+p98+
kL95p/Bxe1qIDkMp04ma5Sjn4Sd42Iu73IuIViG6f0fxonwuc2v+Vz68FJ7H9hZL45AK8GgS/ODe
w011y3MUPuJI219vPTFszNcBAF8ljpmLlwepUzmkdaJPXiqsGqqrYo6iyl/zj5dRrYb/7FcWwA0E
OYa4hytnQLJBAPf5fVg9Q/+aXVUakAK1cktbpZwUqdluhmuds82JII3GMaTFWpXQoUIyBEjNYY0d
L5kLt74p3+29/dkpuq8TDkgDvpPCMJZzZKGOjaI//VltL/wukj7l5nI8Lqq45ZASPg4K7GJIutjq
8z7guTuxBV24yqvmrSYVF9NsltB/kbnRctytcXXWuz3D7LrLwyEDqXUpsAzpoyEDVb55UZr8oVQa
YAikAXr5c6YkWzIN5EANBlOBFGv22gRhSjk2gcXXCTqydF7dMtQG4jTIlaNnOqRzdSLd+2c49Na8
ZF2b5nd45Fzx5mbSvAakbwn+3pS+tR3pt3NA88J5hUVnQoswoPQeoXRBDeiBCxM1HV/E+udYwm47
IkmPLlTgdpmlkA42xOGXkDyeOJ4qFcFkwiW/u4xm5MV4LZz+NhLsHSDb9X1eXrPMtbzkhCjMd1m4
pUIKeVb2GZjjgeGC1oN7uheZnHtoKnY1VFCxmpLwhqI8T8IloP1II3Atd7XAgq8EKpjJvHpstzHy
aG0mqBFh/OECBYvY/8w74gN3y9LAXJMdhA3xpl0/fc9krdxPxlv6dWPqiCBxKjAmbITtdNRrFPpy
a7pRrrRZE+HbQc4vjIP/L0i+2QTVc+PSFWjUdKGL/gugPwi+8H376jaQTFaTv4wLX3KtxPClhpyS
DPM1K5Dbj7FsMWg3Bk+wDBK1VtjcTZ5nQv42N3UqYY2YE/CS3YK+frV8S6afxAEDjPopEjCIN+ma
a6fS2jpR8u4UubvdrZ5biDuyUFg1FxNLJHSFnSAuom1AHj/pLPRKPBrDvBVH9IkVbkj1xNXePQuY
2IwlrWYX/Xyd50ikOlbmCdn8rvXAXoR2ImufS8KSlSCE+qLfTmTV0sW4hxO8fuBsOUcYjWWGe0FK
aWgc0ot4DBOed8jm5fXtDJb1Yn57/WfX/Xfcyv4MOPQY0J5PFIuZY8umuQQjjNzHRmgby0US1d/t
rFmoAjQLZaLSYh94WPJT+0FOIq4I4IdN/YOb+u4+IdpfIKgS3PeXFuDDjBeGz3lD1/U0iTvkO8yj
zbBMFeCBZe5MCYgNI3ZGHQXd9CDZqbrl12H+LH/dwAHWQYYS/j53dNB5mUDpqltrNUCcqpcdIPeD
p/o/tW+mC67UsPuUK8pa1WYzHQIcJRmlSU4IkGUspNG+pJRbjtPCjkeao61ZNdA7FzX99SoPCYQV
EsuR30XedUeIlmv5rrc3fZWvYvDpapPV3R3ED9U3NgwzPCs8WF8H30/SxnpzGIjsP2+VaeEDX01p
t1y4pW4luBF7je68VhZ/Bxsfwsub2a/zIZYHqUUZ1sQhsedfWd1ofee6LCCR/0eFa9iFal8iCpTk
s6BTJp0SrIH/LtmpDxz9KiiSATrbWnv4VduNttWgC939GelpHijXsFhAFe00l0GkwpAaVruGWEjF
XqlJlaHzC1n0OWbfPpBJxRACRBf4obqyvvvIB0dGjuu+O/R8BghfqKHAmynZdsKZukQKQ6ANmD2Y
z6GK5xEHxvM8B5NX/2yZBKZsA2dbWDdxAFh41VvtsKVduay8XjGp6nqIUDWM+goBTiTAvbO+LHEI
jZPXxKzvq9mdyUUTVjozirYVCIm3G1vVTILEKC8cDSZztGyLR00AeCkoRt9zPzEg8+PrWOQKp0Im
qT0yiWPP5GUEidS6Al7N6ZKh7AcwgF1NxETenhBDsX7swZ9Wx9lTSNVtidWlIhDZ2vaYdkKxXct8
ZDsISZr1CfjcMsf0ApGIuo5a+PP3VCO7C8oi+90nszo3HyKfR0UddROoj4kMvDysE9hFO0m5Sihi
0FvqAc1kBWEdjEcFWaS8X/EGZu2SpJVqx+yjWrcFrdwjUJg4+KUjLp/TG5XBFv1iRyAmoVFkFzuX
ZTlfEN4o+yYJ5dewSZZogQj3CZMn6k+VsvuAQmXfHBPs6calA2wNNwOrau+XUPdzOOOm6MH488vZ
URZlUV4bh3f8RqISeyd0hROLimN8bAFybs4+22jy+iZ/RrKjI0U0Y27wIJ+8hYeIlLbxHiY3ixek
PxH1fYT1zFJ1j1G+8Z6hG+mH3YjopJWmUujTmqTMx0zsjySwx8fKQ+D6RC7IXkHBwZ8zC7buMVHM
eu5f/2sB4rTYoqHix/rsWrbn2nDlGB+rND03XaIUsZK14uU8d+/g9u/wNsF9AuRMzwsMBlVTnUvV
YqWyZOCkcZYYFlJPB/sONlYuPvmvWm0s+b+LmCI+f2ZscmhHxW8SurMiLqdsF1XOZJx3XvB6zr3l
y34Ojn7nOqaajApscENUXKWQTwe43CZu3p10dz0YtVjAVnxAqIqSJvhVV5Cs9BJ5HcWzTNd3GoSa
3mekxxiaKYuskdh2marM9fO0FHIpSPiihkUpd3MHcRCV7ARx8YnENR2+4a9Am4f5NekbhSXM9dG8
AtT1MJvl8oSNdOQZ7PXWYBXZnEfrDjvI4TH6qYhTaLdXusDDIleohTcnkL55g+Jp/0aVRQ1OIOkX
6ulgGhfFBERfIWzUkT9m0Vs9wBw5++y8Z+7qAFXvAZ0ViIiD/549FLs/oufZ5eCyckVd58eYF8dH
hYQsgiEyxltkRop2EXH9PhRcTBU5KBsXOUwjX2DRo4J9riERCf79JjBDRuG39izevAKaZwGNdwG6
UMMpwwnzC1uFjXpl7kldBA605wl28vrPdv/ue12megTr2YWfD4w89scd+YmHHI8aEmbYvfDs2+9E
yA4dNVF2uY0aCSoiRkLLvFdFpjF1adA49+UkNYAxvUjCoO/hL7g5x29kTFWRNwTTbl11QnmKPvzL
2z5njLSGOO8mbZ3/Zwy8U74OJqmUuwd8u/d4DXUW8cJJ/XiMwSlMKfd8fMCBBia7gFLX3w/ClOuw
mJwC36U80ZFLVWgd6cr+H678hZdVlBsM7dZq5rsyA/qNcjxXzjCSc6G0muuwTJtzOy9pc0wGsP9H
AKqucWt2AU7PcMSvBhgQr4gfUCOYMKZQJXG1fCSqn26uit9Id6L3u7HYDtXwqXYL4cLM79J6U9k9
lJKQUAO29W6kWpMZujJdagzgXKdgAPR6Vzcp+NWmrudBG6y3tK9slpRUv0rlNO1lbICVzoONJcvF
NFFakq6j5NaW20QpoQMa4PiN6LsXE8dH5Qojek8YT8CMJln6D71DKocVHh9Mhj8tQk1NUczlvE9P
f5bUec8nMt/Smh72yQxIt8QL6AydiB2Mm8tGZoR5r5svLhqNq9dl7w0wpibwNqBzKIQbc7IkN6M1
b/FKWIouDptjjNW9QbduSf/lHpEYqofi+uAWEm2T/XnRlKwYUmCXTx6ATY+IrRS2yxz5zPpNeGnQ
cms1ds23DIqBLbsYQgvojSeBNboig19rnFHHizA8tGbyL3aL+5pQLxjijJzcOeTEugE+qJm2lx0R
VOhzCWsIvfRh1LUPVwcBlkKPi7WzF0zbDe7tkXou06W6G7yghxMLYbyRRVCT5RLOv9gItk01EptG
wWp5YBR8g13aNZEvWPZ40lGGFTqmvg4ps9e/6rJS3dvqIcdATNaFes8sR+NuEA7Yw2BlN1fT0rfN
chsuehwa0/gnsh3n52ekoE5q4o+tdPqsvRZYBKAigrGLxVcPb49VDPooQ9Qwkvf3omgtjpPG+MdB
JyZCHSpcfGhFGVIzx2d6ak89Xo47zkQb0KmqNKM6kvqFxZFhtnd6A2tlg+oYoI2RZBwjUX98p9D0
fuIzsJ0QPXP65v5hKO5i08tYdObQPTXlFmjJaoa3p6k2RuM+XoMZG883dlLaUXf3c4aSR5BcYSBb
1l/ZOCiaBt/lx0cwfTholhhV/n+LhecuCiR/zmEaj0qvD7e5IAYfb4nHV95MfpnRN1Ursr3woKkH
4KXB8Ou/5o3GzzqbJrGnAGejC/2mhs+OLfPpFfw+WmJ+mNvjvAqkeWkmKlSvUH8YbCjrDhveVQML
P3fFAB1+Qpezlw23vULVbC9xys0+0/9l3/znoAh3MBMLHkF7/NDr8151qouTDF9Ysrk57N1NgRME
F3tXDyjN9n67usYXRhmp+mNSf/UQnYjStVw8wwaNNavvC+G90kSx1zw3b5n+JMVRQ2i5qSGxkbEP
TZWj7WBpof0uUzfzfU2QoKG8p0A/8pyQlaXmDBnRcNs07ZOr+Z+/4xC69orjUl9l828n1a3uWluZ
mvQ0qul0tD/Y7OIXRJCkhZEAHnFfZq6bdZScZu9NsKXv3KaC14aSM/X+6GBxFlZDfu1jB/kgzpg+
mT3Y1HhT4xiZ6NiI63r5PUJ/4KTsGPPdw3eGv9vynYMOkOitniJSyp94nePmzIRPKs56rZE0C9/8
x3a0jHzaLd9H6Mp7iaqvN5d7LbAu2NRAahvHLlblo/fwVe9TRpwKTNwURBIInYvljXDnz2frWBwq
7s2S2YhOiCFSUzACQI4EBB7hMM6p1RUwvu55ADggHwkvpXWIdHluj8gtW1Ev5aN8UKLJjBBRxuxG
g/Eiqga6hGm4LOZhVK614w2QUR9n7XzxvnwsfgN/oqhSjCGehXZ55QTlqvUlGyifEjfP8SdkKQa1
kmRwXw9j7Id+gosAGGMP/lsVtv4XPXhYcur1SmEU7KkaoQcpsrJMX5RR7Xr5Ib8QjCN/GqCMUHlX
G3P6pBPfCun3JQF9QvmHV6PoNCxbonWD7KYieKkunxeVue8PirIt3Cyg0Q9ayXUJuN5ALeLpz6Sm
xafnOBj+U/7duZ+zpqK2Acv3YohzN9333N6SksX4K+DZrlgyG+TkYll6RQziumBTIU7/EWxY2KET
OUx3cVkaAcB2Iqd4xTm2nc7i+a356R6I0X9z19jcKiyOelmSqcDBsxe/wRzaxzRNhjtR6OpsVI6B
XsVk0FxGix6kE+sjdhbvg16bLJRqzApU+dFo0nGt/IYEW2pMk8KSD2/Wuo3HJQ507Eq+yAoKAUtT
itk8i72EINPuKEc/EAnk6lRcmtT+9f3r+uP1tcuFhGuIdU3f0px1/Jj5OqHVGmk81XAAkZeYPCxI
Gjiu9G4tBij47EstB1b5fDpAbSlN9hlhF0LZe68pvMnI1qiAd7k2BbmQKXPWiQCXHdapgvxAoaQN
V0XUNTTWUkn0VdFUe+WLBp7OtemEF9p7yNCUUioFaHlkVA/mXbMfXbUKNJzV063yXoPQrzbnjgvG
KAmAao3XT9+vM4vMOlcPUCKFpArfYdfhE2UREbqYUdAeXPBPrO0kCRwV33ugwrxZtSNVPxIJCqvH
0HyWlr8fuiIqrVWGLL5Y1zx+Olby2tveFYuI3Ieawx/Iny755dp1/VuLWYzxM53Kh7c2xSGEEVo9
7j8uOfp9jLK1HYXEiE+DiK/E7xw/Yckft+fVhZa/hYL4kQHA0OACvuQiHcND1WFOmz8DuS4BBYsZ
weQI9FsDfe4YVkBqB81R7oolAAycK/ZsNc3B5ym6aMm64fY2u14+o4z8pjNF3K40uRno8PAp5ukq
wE1Pu5E7ptUrtch1ASSALVM8gPTBV1WGnew2OXdjrm1WBw7ePQ2k7M1s4FlUzERVjeOzIACtwjMd
k3Z3ypOPJgjcpu+t5IeiTFXWcWoWWW8zajmw8G/9059A6YC8w6snJNly0yhZ1PKudTe5kbHKD4sK
fRSWI7UnX6IKye408ki47mITO2kLA0Tta/XhQrqDryeXezioZL2xPxq2yFHqXl42E1dqshPKCI7i
4WKDVyfWOMtw6sX2ewz7VpgjJmBkQqh6b/rGaF9bk7b8mrBpMbNPXtMol/Yy8RstXU2lcqH4wyz0
OEeqk9IsNwDyXD1IqDcgho36S5HG24WyYXBwqFtDV340ay/HsC8RvRnJKHOxEf0PMYKwEiBQCfDU
8REi6AK6Pp7g2SQaQp3xnH1mobohLKvlwF/lbL3oxGCUc5nTxVAkCR/kJxcLvdJaN4U0Am5KL6md
8KnXyRCw/GIYiK/MnrX1eMxoABP7yc2dTLHikmVMNJ8pH2D40Nmn5yotvONjiWhbAVTji5xPvnwK
ZEWPY7tjwnRVYUZL2SV7rzTBfNDhL6NTz33KtolMEV0AtlubwJ37oyI9uYzv5gFHeG5ueHssleyq
Og4hEioj8dA2nlieIqN/7SIlOh6usVQouRAbDwico/cVyWWq1ZlvmGZvQJEzhBiE02A6CJ29ByLq
FtjmcBjvFnuieG1EQpr2aQ0tBlYxkDTCmW2UPn9fblu8lLH0+waRL51yjDy4EXxrquMPgYqyZ8Oq
Le91hdlhRLpp9HFBcFbygH4jkeilwrg7tQL1Ae8gBAc/tGLVQdF1zekpG84B5ByOLjO/tPz3IfxG
jDHKzVhNaSQ/ENDsy0wp/nSMwGdbHa2UjpFYewP39Sxg4XiuHOfgn0xTAeA+3rvwQ5OuiAR1M/go
EZkzAqHY+wHWsBAGhj7WtvCO1U9BYoHIZB5llUn3PTEit7A86tNKPT+PPIBzrNQb7+MgNBsxvaJa
ScQN2oXUWxYwPG9HozHcWgzHV63sGqYy00q8XP8mk+SL0GkbWhVSUfUQ0bxO8S3WRU6xfRD6QsuS
zE2dkcS9wm40im2NuKygsCKNCebq0u7VNCOO4TYiEK0UA1iAb6r9HxxxQsGGojYpP3zgr0WBa/BO
xkSvayJ9aWOXS7u9AWiHvqoOka/4UUjVpNCYHAEm3aqc1WefNgi8z65oznsA32HyZy4ZyiZFZiw2
Trt3jTMKQq3Sq1eje9MmbBcH17Kq4Vxp3jh1Dmg9DgXGjY9BMlr/kPC8SEjGfcD2ojV2NbdwuFH2
rpdgsyIf0BvF0TR6/8QZrqfWCTvKeiWnfJX7drCJMMDNBk4c7KFEIQQpdDorohbtVPxVmFNdQbBv
zs1HJzUUj3pLwKfBy9tEH1OuO5JvRCcuQ2leOb+7p012vLohAynzYya4aDgiwq6xRUMkfHxvDlQ6
ER/syL8VlnRjTy44k3wa9qFewpYcJlXUiIy2gigTpLnuMrRPUA1FykhfpBU2R+lU3FZyfGPPeORU
LKpfrjscXrFxBZ8P+yUBg+mnn/Uv09AUBvLD+27h1hgwAKZF1K5G/lydhJ+XtRoYHE2KAxaiALpR
A9kmTsh8wBDt6+y2LazfMy+SuMkjAPeKLJ5O98yGKZhXF0etEznkKXe3nEJEx1kRe08LACqDnjMS
Yx418IhSG5cK5MuRiU1DMU9HzeGXGaUQLpggrGkU0RLdliNTMh0yCjYaSMrrM4TSn3fvr9jIxW+X
Doutpv5YNRH6E4obXxH1IA2LxwfP6XvAoOO1KQmmENwZ+enDqjHk7NlHDXsiKYtbWye4LSUKp227
7yngkeukWx32URJ6xcIj2IKgnF3jXv9f4vyr73wogr6jmBBlxbg4n6NuejiEaa0XfpbbsMbS9aN1
D4eudw+Wx+3nAiZFx4eqzDPrA2cb5TUP9I/uVV2QVhI4+lXqVnaJCaMq+FBmKrd3XdraFlq20DMQ
7vig2iVd1mmFIwbQFoC5ojoOraKhmZZ6IJmttXm51AXecwa4SOuRGOX/G4Feh4fC3X3DLT/KpNw+
oA974ibBHXErbU0IDMScYE+Bysdsz1Otn9S7TJz1d2W4dywdk9VoCWtIZLlPP5Jc9JQCOtsQDpSH
ygv4k6iq7AIWNxz3MpBHs6N/IySxVElotiI0M9rELdvwboTJ7GknxoAFMZ2C3HB7V0RGNw/3HY6q
MGZFSVecipvdbT4bSsxQqK53pIBWlpOi9psfkLcpjw/4I6Oo28fx1oB3FNC1SwrouIjQzFCPafiu
apj3HGyeRn7vl0zB4lsmxSsWKmOfgd3XfHzwgDqWmVVmXKa3ercd1hAFBm0u9bisI2muFc/WgOJB
xMVpdI0VcTXKkHVTWRtoHoYAGKwzF8aWoSegTn0WwaSsjrxN65pCBXxHV8LyUR5p560LPG3Z6+I/
B5KVLVk/cZ/HhZTbbX/r+Q6S8orxbPqVSIk7itMI86VxDN/uc/vu0/exXSjs83JvjRAM/KgN9Z+1
gZadxc+dKFzKtwr/mIInjVO2GhI9/zJB39rAzOX09Uq55bsBcKIjwQb9DPRsT/Y4f9BBHDTJwjYy
wp8SS3QYpdjpUTX77a+jRE7gOkNr62+rWkFL1EqZ1WGTD2Hynq4EBr2UNcXUlmLO2Ks6r5AgUIHz
h5A072QWdZfzIgIsDqCLAyJedx0DI6kAYpXJFhIn7+dnFRCX6Kh+UeNNkvLucL4goFOSwaLj4lem
BWU/Cs/sbVikt28fDoazYwz7sUzHMMSfcPOwkT404d/9E9kp2vLdsIdPNYb9Wvx8wQDhb1AIJZlX
Fte4nCBgHxhWt5TFtSutaUP5qQChXZcMkp6y2lkueFdAmq/U4jrMMWnyqeMZVKchhlp3Bs9Lcmty
2NkvWy8R+gxF8Wv9K/77GJVD0W8jdGw86er0SZbtZ8hUdK9ltTllUe4TEYkFRyTdXYedvJNnBnsd
wIVvkyJbxic14ydyC7FfxjEdrzAmiKEMe2URuysn3weyu2Ck/T0PkZp5nR4MTTu1HRexq5I8uodd
SrkJsbF4CZYboJ2/9pdocS/2T1Ojzmgz5NJm2+gYxYfb3vlR1KqZYDxDTWOBTs1axQjZhC3IhhaG
sZV09Gx860iHSTRskbfJcl8Bx9fjHFvAQoSRhzJnZ2LgbVTkeBQPoIuGODm6dsslan/aeaIRmJl5
/tBqZ+zjvQ8/6kVtSzAbNTMs/au8RXVKMjl/nsLNPcn2rmIqXkZ+M8GBM5Qbh3LzxkkAUupHG4Sw
nVyPeJ3rDpyUUp9wEBCRPG5IWkW2VM21vFySYOdcxnXZVu5vUWBX3SYPt/AmwOIpjMKjt2LJRSe1
i9fzpYzvVTILz4dr+CeUPtkP3ugMNsK258MqPLKaHkrsBbSjXbzj3vHmFUl5RTmclT3sh7k4fFc/
XScDxNXZbZ65XjHdea5ppMUrWWrDOlklkYykiJDnNVMnx7YxPg3zliJ6WLiSzbm8ex68Gdk13lsH
ZWeKp6cEb3T9cP5Yqa+1moquZ1Jr+nTb+dPdngddnkCZ5a6eRsT298FgfVDRTwYLZGPPaSohSnr9
FzF8T5CN6WSipLMiVoqN31CQjaJdgqvAShywBfgqweri1yqjMHvytkhTHgvPe/hmN8h8Byd02so4
sHIpj6ta2nRkbmI5bpwOJEgYx+ZuObYRkkDdCabaBEMODucfZfEM9Vcltl0DGKrFdcaNRyPeuM6c
1MiX6IWs8gtRit72ZOjH1vq9lL0vcv2asPcKcBmkzN5tjBOHsRHRV3IfDm3wmrDrVJdYQC33v1at
G82ixxt6YUqL+VAcsnFlibT0zneL+jDbuegIA1Vx0z5UWdqoyKHTcuL5RKSYVwukHXDxV5UYZyle
f0yXnJFxsbx07XD5uZsrrMwSYCW+Mu2Sc6yAfOKda/m6ECv2/0dNtOeb/RY8ICyr85qObaoPT4yF
tnbNIK6k5KY8tjX21uMIB7T7mbSiZ/i+gg0vluaLWrn8fTi+r05Q7RUv/c3TvvlDvf8GtGeZ0vEo
rZ5zj9vpV+Tb+UhhR78ZRJhgH0oWvpZLheFl8Mvy0ZgGYlEkBAYHFapObSnAOx67jG9UPU4IBTJM
cnE4YTkwqiTAZ2WUXj9PHHdfCgVujdCLGeF2p5VDBDp3Zjz3bQkxayMrE8YnpHf0iqzmF+MEcrsr
wTOjuqQa6Tv19C44XFWirwKfmin890HgtbYnwyvii2eP66VnK5bH2oA6QXsuKxlKdn36hEnJbJo/
JmYKyEJfqLTxJNbd41Ap2JeizxeacVqZoqt+kugA442b02CEdw0z656DzJPWbDIJZL5JHhzq31rR
r2z8HR8E574/dCUZDNnOEnlxyZ5MBydx7yMFoyeE+uZetFk67rYbzSglszqv4mrZ9TySo5+rnXuT
rvsPfIHWGupfHF1IcMZCjG5HKjkhampIgKSJqc8bfSzQdiQMQrD64Uj0D2FVcV7b1Fz5SvgYsjtV
y7GBXLWdPLujj2vX4Q0JOsSIlL5m8iYifll1WX8zzIebubEWWWEznep+oa3hQBM3q6/ay/QnDRwe
DN+hcLylnHsxsPITaHXJ06TVrFGQZtPzWU6at0DSSHyv+C6O3QiDu9IbfCZuB02b58eqeLjaMEU5
BpFNp2J7HKPkGRSwcyHhO8ll8MJPS9QWKm49pSjz56gpW4CT1+gj0v8/dbnH9JTpwXDgtxgcj+0g
cHySHnbmpduKLT/fjyr8TV7FsGnhRk9uxFcEncCRISx0GRx7+hddicc8KGCYHKFJStcCq/NlXBpA
zOx2Q1Fc0y57LlKqlyOKl5xx+Z+e/RqA2JfyEaK+5TZlY417d0b4bAioJ4gqsmS9mvxykXg5Lpge
mfb374GbAXO7GUNsp35GDzVAQbXrjN4+7kThrTmY7gW+cKmzHzf+bt/jzuIa6wC08PvvT2cKQ9UN
I3NqAit7oszRaA2YqlpsyzL2R+QH5iRAp0OUegnRrnbUeCLonDd3cOzOdLtU7Smd643WECRF1pk8
kxQu1x9BOwbUF7DatEfDjHpLsMhaZVBe5IHtBVORlvwhWXnoLm+/JqpkZAdg9Ct8OacazkeRdAJS
O7+ZN4hZ05CFGJiThsUxMCG6TpGDt2lvoo4cIF/uLBCry13uHg4f53kuGgNnIzTaVPvuh+ElLQ9L
iNF1GnJkZBW0SFpbNzwZpIV3mEGAZZlflKSxdmgmnVT6lVHe8HSF/eDPCYuQbQ9wbPwVkLHwUfbP
6lDGmZbeVKPvnPrvMTnCyeCnig9ILLMwjntscw3mQ+Ozz+hScYZgnEoxcyKOXn+Ttrl07aMqAOav
fUXK614jtjtRFM5qAi1pSLqqL++jaI2wccHcuE6YwY76gMg6gXTb1LBZZ3FSD5UsNYOqv1HKTKgX
9GG2eXCGlOUB0WWNqFuR28VQ1IAvFvQpxGP36zc1tiGpaIyarQfNO+4+4ppgXv3CUIZFeQb/WZSU
rsW1O3mbdffyvmcBr6Rz+ME4/b5nsUBUOSyMCo3pQ9B+oiPGiY+zS5B8bLW8A6ICDoNJbwMOGf5X
5naUfZCxSICa80zozNAXYVH0AN6BxWAhs3V5ND1HAuPzOdDofSIdr7fWXaKJgObI1Q2qCcWq0yev
T55Kda11m+7M4nf2r0CnL+WsatGzBwJi7czJx/KlCMU0yVeguH8x0x/G4uAQdax6rCJiGpnFmAvp
qU8+FK+KVWUlyF/lf4J5GNFYAmJaqqDuQM2EkRRCWvPFplwj9etmEq9dd/S+vAgaDzJmkKMoh+S5
YW9+qivXzvTmD2EMd9TGv93q0BMXMK+Nz7SgcZzt4o0i9Zrc/YSdgGf0thfYviYgJSfeqgKVi5ke
WN9Y1tZGnYi8frFQPwaphBXBUmMrsh+42hOL2VNvLrO7c5Nsjui6iGWmZ1ODaeq3TfPINCDupMqe
MKhs3f0j/JP1WH4RfJHQcd2/tfVbfmG7n4WhpQUy7iDgAjNLBkOFUB0Ssyt68BEqt1mgbUTPRwjC
vZB57WL3UfmaEXajD62HwSzuAngChKdi1NMfh6cgXvfp9EBuNmmREPMqoZnXlpyChGOhmye0yVD2
mv6PZmMNoFcwM8ORqWefluKXiJw702h30u1r+P9MI9Ddfx1dCo5A1ADv4B59Cpi6gKuv5mn9U6/g
F9y9qEvHZEl3Z13nfJlFpV0P96g6t8l1tXA6OO048ip4nGeDUHTtz41/u0xPQu67F0deHSds1Li1
r7JzeMHuNiaEYHnLJjrciSMnbr5+pDDdUmomTdbIaHNjxEf+7FPw3N9fDrHMy5SMOQDGqX9OMA6Z
l2zZvz2ZsW5VNrgJO+3/9mJUZtek2WSiXmw8NOt+EK1FpUlWkOf0Y+7YsUo8Msocjf9cv1MUSE2Z
Zzc/1lV06dBFBh+FmN21SdjRjQdq1pZeJb8QlOZzs4pqEnu8mG3xyV5x207o6+D4ZbHv4uYv/v3Z
R9TN75MzsgEvv2hT1wmc/g9j8NaXjzBcqSuc5HneJUQczpUG1C74pyC83tCKqzcMEGUfnAucO9Z8
CtUzVl4UUb3K/fYov4fPzfzAN9lKJXpc2XvXg63d6g19C8vy1fE+Bb6Q5PM7LCOW1SpV0rZTY+V7
MFJo/fE0Ukafw4gMyBG+xkMXxqnFnmJ8bagNx+2l6wHwZVZtlynMNjItedlTcmPG83KtTgB60kXf
GyBFa/BVRTJRFwTD0M5H6Tg6qhzGhhwyuCJhHoyC8ZxWn/E80kQG5xv7giSizc3LR7GzLwsiIIhU
ilaEYAFqhfPE2NALwhhOvVsef6d4lDg1jSHHLj9u7nBITfYmAhgt9aUh75O1A2kync/UkxIu6ixc
3D/3KKvsO57G+BWaY7F1iNpx8zdbNhIHLd14GGUEj0WrFU13e6GvYibmBdoILrK37OBMs1+uhRs9
t8Z7ykJolTV0pxeAj9P4+DDfwytmnX+GptTcv/wXKzNoE76XXIiUDo+pVr1ayOLaYIrTCjYNECpD
v9+yw9I8PVeghQ15vtsnblhwn9VKUXa3VrE9kQEAs/HSrSabdOOUtbiK4ENADiPb6ohEEY64t2/J
EpAoS7IX2aPR2dKwFmNwdXcZ6mJslFcGBZ/hRdv8gIYMwIF3TWXxjDIL4eIL8XBmmQ7X7bnTBQCk
XsNOH39VNgvRbal3t2a+nfxrHRayf5oqDcwrMJW+C+qJTmsPCT2bAloZxw4ZWmgFyQJ5uJ1+mVQ0
j2diQExPnKIhsr9xL9V1yPQMDvOxx9bb8Fot/J3Xmc56x8TZlO+iBh6PDnxN9owim5fibrzzpCfg
6jko7UiQ3M12YuA7VCq45oZC5TEB68tc1fqyd8XWy0WthaPvq7UPHHt05p1jJqbRcELpQL/kroEV
DosR5wJ/8TLooe1uU6fZir3nKz26PSNcJXsgzZrVKX59qbDjrNTJOjMbubuM8dynndnIczI5goS8
3ouK8bpV1ZetypFNw3JNJu59yU6BUaKZNkkSx5y9vvAq4W7Uw4jcMcAjzI+GR6dS9PDRNkYYC5y7
bBFYkiDpKh31JprHFQS9iFhjw+cv2leXJuT2kqyPC5+LAN8K720thcKBsiJhQdbfZaf7N7I9Ygww
m8Oh5Ulvu/Vzk0cp7S48xWNRY5Do8dNRs8OZF/K0d/1DA/BkpOrn5gzm68rfI62O3RCayAnB3gsm
g10ylq5oq2Ic0DSXeYpTEPiWQtbWbY/tJud8PTCqoqX/01gJzf5LZl3oatFh4mjZ5fUoiKFr6ZjS
La/HcTRiMamRWvkvTBhziwpgiTKUdN/wjQGVeO+IB8QHmqvRxqv0FGUZ7ElZ0ctkT49Gb9c33V6w
xWm/zgmX/0+E0yoX0ZQWGAXy5eF5nwYXC65L8uJYzwiJCy/D50Cd3v18SUWImoU00rNAS7o1epoO
IlONvKHbq03AaQhbZxUshivqaT3t17WAqQQWP9aqYrW13WZw01Mj/Bf1qRyr9wPANBAN8vrgK/Hz
GYzpmBfPD8KR9TTIaaoAxPh4E/n5E8z4eFkdQxLNxKV7TwiFYdWwEjLV3RaY0aEw2cyFzMoLUUIC
ARfmKTzxriwo7HeZwMJpqS0bcve7YJ4R1po/bGoG73spuku3UA2GT/Z0/8LCXcxQMlEhoL0WBapN
y4bycmb0X2FdTdtgoz2C9hmmIkez/5Dsq3CYQmA1WL4CS6uFlSsUDUnwOxSsPaFNr/XqOnGF1MnV
DEttCwX1N2MzCZqmH9I47EoHOObaiORNKXHOl1DjJLIrZnbyENcj2ZRrV479L5ABwwD/xiTHWHXL
NAyuVbykwzLBpYNwJqylH9aL9S87g3+CnXVn3iHLAJnsBSM9C9GFtb2pRBIgmpRmvy7y0GLwfNnE
XSgCIatAFYdDiiV/De19RQ9XbZQv8/KfB5eU81YE4gYgtbn91xocP8UxN75orXZ21eLZTD47LOdO
Y31+nkgQ7thyZelsSU+pLZLu/Vf8wLWlhpUHcsQt6W8J9KFkyIFK6IM48Ls7eQIHCqn7KV8Jspnj
afIuDa5wE8jDdUF+47uMdabyrb1zOS+uBXKKX8ry98Dgec0zGtR5+6f63aGDbSNwC0S4l7vby8px
WS3+zLzRhG8903h9ze7ixTrTp5onCDJ66P5o+y6V2UlB4DlXUUY/xqSt7UVg/x6AzVnE6p+cjjFA
IH0+Xfg9w0NV0a62LMUQnuBKh1OJwtNxBIAQPtjGvq2hjh41l+aGd4heR60UI3sk+pDUAbxmhfdS
W8sAOHB/3WZmxg0cJKHCETJlYDUXuFk6+WScFELpMVjWHbTCuPAt9lSpGKTD0EEPE0pnwzHSVpUw
hMDKLwSuF3/js/Dzhr00vg3y33M7OHHfsivJHvCPmSVfNaqGLpS+YMYZUa4BGMq6B1Of2CXieyAK
K6tQHSggaoVLSQEct6jFvb1rJa3Rb8kNem0Y1anf9BtxeDd8xPQy6Gs52Kx6z/8lkTkiWSs7cVW6
nmmoqAzip93jY8YdCQoxMjOOkp0G41VRBeS8DzL5tH0K22fPz2Inixs5tizGGK0YSPeTP3bqqNpr
SMBumEZkjOhbb9tFJY6uF2sTS3GCmQcJDfwhmWg9djS4yqPIX26AEbbe627mZ9MUs0X4bLKvA/RA
so+wp5VDgbcrm9/NU2U/B7hPEpupNY8kzjhe290D2axnlzyGqY0+gQxLay4FjS/4DiLDSgQCHIlk
O6jhWEV3GYQNu3v4tviIST8TONH50r4TpPs1c8Cy5eKNbNgPKTLvwnu8n2GLzVnfYRXb8Mj+3Bi0
s+L/5VgKQg6F/Hh20fQg+kzffnhZbJjEJQI0xgckQd1rNgD9pN1SO69HPzbekYRiPnxK5pWpL80J
pcz5ofOK6uUXirP2q2rolU6hI/DQx9oGM8QqFP0NqHTWmV+NxdtyG+6cYK4Qri7g3r+rLU8ZdCgR
fxN1SSY6PWipZybMTBRh8B1DDUok9hYnSJmp8kVsVZCU4j9TVsffLQJxr9VYGrCp+fK5CytrrHnN
AFAZSMw2PiarzQDd1qI8oZ2/CpqKBQRYPLSrF30uQ9ySlMhKFaMYml6uKPMk3ZXjMYSj2YtweVOs
Yz+gKFmBo/N2CwtAnpcYVJG5LIfKq0jVS1/03sv/oYjeS1pPfjNYNL8dpulRrTR/yHFEd7Npafox
0gzW+5KCBFuw1Glwac9v2WlcFG/TEcwSmyLf+/73zdt7nUltbMLwkZyVMpSZ3JfUJI2rSUD0AqCI
+RntcSNM2VdYPdo915VLj5/O6WDSnxQrN7B9XxhxUuxPqUK0u/mWtfmU6bjY2bhf4ZcEgugqkEM2
Xnp9U48uhUeXH1mFYtBwJ8O7+OjatpQ4lDTvC/bBvVWVKWvcpdtlb1H5N4MLfdbk4xn8KV2/WQdI
c1obfF9TxjL/SmIS5u+X8ShbBL2HIgQ993mW9IpvS/v97UGrHpMJ4fUQBySA86IzJhqPUrpRMyRh
T6MSj88rV6CIw8sacNT5FP7bbuKM+i00IvcYNmyZg4E8hDp5wArfjMpvQfVE58EvuIL+Q8zn0THp
06WVUkt+y7f5lhj8BB6xE7QZhRd8hy50HXeqxv4mQ4wKr2X4UvEmq0UWhOo6YIqReGn6w7c1TmpG
vdQqXHPUomQUnOOfR8DaAOe1BdW5+pMeehDRlQ1xxL8FuzNyUEFUx7nB/cM99thLh4MjZ+zCARfE
zHs5Kk5QxiBImnZPzGTIfvHW7yfp7TrmsIDD6MBm59ZhoI4OHvHQzQqXgcsw5kfNvLTCQ5IMzDxw
byOng30QvWD5E0/olqVa3LyxCxyNg7lOTWBMGrSDHNAKlwu/W9/mvX63klNktxwq4Zsi8+6Z88MN
nqZprtIWM1PC6psY1q8oVEV7CrF6+G8Z+rI4TJY880M0/N72rIAGgn0v2T2Dtp6DwPxky+pqtrDM
vuOHeYzmh7JqQy1aUbmkBLrVZixLvqD2LFf83xvtsyXn4Eren+GoTDxtOOyc6ZNfk9kE9kll0Ob4
rJ0O1BdIAYhj64W7ohTLPWgo5KV4ihNry8yZFukSjEsuT2mRnLPUOyOktOfzugQX5jLsVphIjNDr
6FKcuXTsXBWtlPeognvHx1vzQnZ3j7JtT9WVxjWXtbCpLEtXLH2jSvinR9h8OWjaXMuM1D5NDtPD
e09CIyQtHAYEUgdC7YZBdXuM3HEVH0njKCTp0Z1vMzS6Q5OHJlF7CKXro35xtMNvJxRKSCOdHR0p
QHUXiZHsa/TKG+LhRChIUXdjIjGyDoLh5EED3RK5L3DwRcAHVn8i2IDSRxoMoEBFxJMCZz+1DjI3
RPpFk5V6u0po0H2Pv9aEbyJSXIOuWfmhhzgI1dkoIbHdnq0lr/fooQ1Qxz4Zg0hCnhWgTctm+5s/
5Ga/cAqNmu+3duki9buMCgmxJDAR5JMOu7AO2RJyyTkFlw3yyzYx8BBmuX9ETsD7hrT9QNxyQ2co
q5bSd7YkhSebQd2GJ0YxgJ0oPp+KIcbnLoltOghEemhcGAud1OPOhs6HO8bKFxap3ZKGTmdA3eo1
1PXKhVeeVuBR+KPPIthRIeQtKfXGfcAr5MW+MAxIc1Aviq5dl+AvNkaXgD2c8fXWiqF47k7/TZMJ
dJPE6ik4GMuBTxClRUSTqP1cUF/cGiQFszkXdecpIZAgMMDdPcG/qx1bGmSnW2nfIIP93wLiRlkV
HLYLe0HQcpfjbacETSy9VBq+plHKqACymsOGbcQa+ldiXeyNEBD/2sYTnKVS/XoQclEwC5YaXMXw
FzfhZemPxGlZCWp/Ov2N+ekpGgv0lzFdKoZKXQQFyLRRimdoQaUqqwNUwRDoYDn6OnRJ0kzU8PXR
GSwbArTwV5WLAFHwlZ7/3x5GgH0IhNN+LKdNxSvpXmfnEWSCHz3XsywPsNxIdGLybI+UWuxKjaCj
RNoLaWMxDhLhqpnQFxQD1j63VJjfX3Ifb0LOudjzbLvLtUrDoa/yvc5Z4UWwXcnpc5k3ueNIw2nz
W6b3l3xkdO5rH7Jq7z4Q31yyqeavbp1/6A1lxyVT3Z19eZ3H8MhwasU6yUOPpPjuwXYL9nFZn1ep
KaBxtVi+iNOOLKgruOFg54APBwVKm7AGAOMPnMyv5fAwBdKG5U3IWRd2FqRTh5ZJ4iRfRXAHsPiQ
3w/O3ARIHB4zcpb1BAxcBuEVbWL3wLdJIouMBnWJqcruBquubM819ADx60GW75W6dD20C8lrJsQS
WZ8Y4scz+OI07oSMOGxG/ZdXnNwkRAAG331S9J2hj4ZY2z8f2BHlDjeejn6mFkTCRul+aUNIkdSj
+dmQ0lspIjZEI2sCXKo9/B74b/j6SQO3MWpw0FYlNT5ki7zgYvVF9rQSdbQdCJdv0+0rutxYwdSK
qa++4+3Qq+WOvONnntiltDq+SGrfM48FZkyJDviobrZNiWhgd3TO84ogony6EEdRyM0mYhcro+RR
qSdeFv4VqhCVp3Dt1lWiQqzBV4cv/QCHsKMtVf9pmnOmxxM5JfUpBxTuG7vGsIO6j07P0Oe5qmx1
1p5yTHKsNXN2e7ZRDXCWW4QcllELZwjjzaOsGv5uqnPzFWHR1rB2vvhOSs/+e2SQUWQ9nfgB6CrB
wk3lNcmyDv6mHgmHL2RwJ6usP3iwhjdjXkTf5cV/EeijpLnPZVhPFTHOkVTKmkNxpwU9/x29MAY0
VRcLvoqnuFdcPehLp8ujxc9fjfpa+jreD46SRfAdrD7m+oYhzrM11ey3StpIRoVz5ZMRIGhUlSfJ
dFSMPyf1QbEq7s7rRGgrW8jUaSI0JN6XpMFB9NU+GPVBXX6Uj2kScmgPYiOTr1iTTBgJ+MNZ7t0+
A2td2oKdQYWSVWHJPhbqLYACmE7AOZWE6p+u11VtukX9zSKS124BkFihA/GImknBDn3zG0Zve/KB
UeEAi6oUjmZkEk1TxjKbqXG99bME56a3YJYj5qsE8JwlgzWnCPHT5AfWh5R3/yX84fkIaOdRwxFw
O5uOUM2brhyaGmOMuEkaA3TkNlVETZmIENwr+Vdz3EMTLECwsBgnlo46S6WlaptvmHUfqnIlANHq
eC4qjxy/yr4YY43kAWp9teHbCoCg2lezDtsxa9wHEPYkvJmyAuoHOC7OpX+V6AgAXK+sjrlSWukx
fc1JlvDFAqenpOxDiBtv04torDriQwXZQ0e3b1srBpXSL64Z6nk5wh3lndug9WKqtM4xexI0EmO5
4wxIu9KY/d842EoQSBdL2IMWxJYPg0Bu6y9eMCor8aBinZzWits61Kk5vOOAGbClQ8jovL7eDEsR
BIZn88SsAV45AMIrSnDLzJTn4bwzd5YHINZAgfyVtzjkeoc+3nBAotF6CzWKH4dT6JLqVkumie0D
668t+zEMQ7xic/Hq7qDfGPHq/0RRC6J32y+nwYD9bRw6HoM1YtaXR9q4vfOXvKis5d1SILaARn7l
YQyozVgsvmgpMcrAoZGwdjxypv5QIZuqFZfy87G4wdwoDmYK9TaVKH5D2BQyICZjAOtTdRHtKuhe
lR6vOB7Lj75jUPXNcZxibgVgsP4uv+VZArJpgG7EBK611saVcLdc6/mbE+7nc8QYYUFWRWh/R44A
6C+18S/vApRcmVPn5oCvvxjb/mbss/5A0L3d3U2DBDp6jIEY8oMevc8IKZXsi29oCgiI5Y+kAPP6
gJcaJ3hWjGDd93At+q36IIyN0ewD438OascfQI8Wq4KupXrj0UpBuwH3HzONf2CIBJlpIcQF/oEX
VWwCQyaLKVjltYMl5r0nMsdka2yDMq/Vha5rRTJeMevmZiOC2TPIscP7+Q4RG60uaHJhmxSGp917
Q9J0o1sxElt9kjgjMUeE0HWwzhOQF5tztRrbI7rhSrnUXeA/fGceO6i4B5KfZcxdC9fAKeisnGDb
NRJWHHQjPqgqldJCp3tvJz0duQu2+zC5Wqh90XxgMlniu8CgWmBOTW5iS1rxihTVQsBYlbFlCgyC
844HZBCLLwXXZf16nQACEZZxvA3rbOpWUNM7AjREO6ObqnVrjM7HaOA1zF5so0GUs+1RIo2EtvCb
rmPxsAyu0VTx/b75qSgtBs50tW2FK4pReGU/LbknQzuLOO8yLhiV9KDnaDmAFkUg8NaKgixTeSLJ
vqAYNKjltVUoRvuPmoMcCcjm0skpivCmR5234PQunS0KjlUWSUtw3GIh7CUZS6GdJ0scyg/DCjWn
0S4UGiOw+eQJ/ma4EFMgDH9Edjmuw+bvvw6DILcO8ibiRxVeIral7iRPic8Eink3xcY+o+fO0xPD
AUNCIjv1lTU+SS2YzXfgRklWCjRXX59swfoP+T9H04VHqFvbbKKj6c4MT1aHy3AnJl305GTzorTx
TXvL1d4D18UIkvf2NZHfpy3sdgpD2iDWRu/VTgbzebZdnZbVCPveOnAf64ARdy7v4NpidybSJR0v
3REyXkf718uJU0Rbxhr/EuhhYZD9qjx3Wr2aYd6Ht0jjSbR4vBDlx5qdgq5Zl2EkO8iJyiMcteuf
tV2aLvMdaQR7IPwiguadbdqF4uaay6vTeKTMem/Igs3U5QjAbNUuQY5rnoxJzsANNYf8Dc5yDcdu
2T6RbGQVldEaWNPd3Z2AgI3P4eZK9zrO423BwFDbJWwKfJrrmwirJYvEElWpQAqpPGC3dL2YDsas
eqOlrptKvD80mlaVReEetnEE4BLFCNBz9PSJU7cWzCHvcbM0RgCDMy2zP+v75Y//JZQwRR1IxvWw
cCf58dPObiqCFZusmixsLfy9YZIj3iMF2jx80YuicD8g+Hv9seSqveevW39GeVpVQ21ycSBY+4AP
XQgyExlDE18FzP3tdCQGY4mZXyUXlhQNAFxT36WAjzUhrLHhhezuBsIjEM1+D5MUqI9fDMhmAw9M
VtlEeYBmi/6HQ/7rMmdAJ2IoTiHXqWYXgAPBsscgT1XorzVBRgmtEzY+ZEIcd1UU5x24Q+A8lwmD
/RG+mq4FNutlIiYJJhvTxQp29Kcbvtuu2Hh2xzclxnJbQUIU+R1Tmi8t0TJ2dA/MOW6qiaecgwI3
QVvG+C12rD8HqqTbjYxWFa/Wyw5Yf6VUl4YXsiivi76eLe/tUjKjqIUc4hzjOgFAIPN/PLcHb5hD
8EU/sVvlCc9DH8Cq/xuBPGEuCa5GvSPLfloDLPjzu/HUGbFtIsL0StXdZhPpvCWCz5j/XNtRZoP9
Bdj782lBLi6cuBvrDw4GMVz1oboLrIaJYWMdJsrS2I5/yPL1VrmBELkBX4OYUGR/+NsGLdjpHeAg
XeY22BMF/dLo7PXG7pCCgTEI1orQAvINCn7+AlSIb7b9ozrxvUAl/Ds12DWV4igMWm5pvY3B7pd4
Yi8Lr3yOmQSeWjOfpEiNy2cICIT7xw/jPX80vM0SwJ5SXt/SqcYiVA1dB9PK0lKCDgogarXNRwhw
XKt5Zj/+9DIV83n6bq4qXGZsM9y+MSTITQahYwoj1FIwdq2vXkkLhiI/Y79JCBLNn/hi7FJwgWez
49hmLp5lEp3NV+o8zvJOIy2Ww/1mzppdW0C6r604/DuTYtTMUj8z9gyyIM5QXWDSbWvkQx7Ypk6m
b+0gVy2vb+dZKyhnes8MVdM/AUaKgnDX1TXltA44Y7z8x0jyvX/yMBZvmUOX5LmvqG8iJrDutWrw
M48UuVDeT2vVo10FHAnxUFXDj2yflb0tLHHcatB5/Uf6uQbaGIUsFl9wuwBjfpqIAmH/kT08K0RT
7TAoDwG4GquVPDGeETS/AUHcJjRU0w0XKC9Th0Ql/Nj80vkOcjngPe74z64yGw23fPviPIcCwm3l
CZ/D0ahO5g4yGsM6xwm3eyKSYkuUZ1uhRPtfgH308D7GaaY8CPswrbJu0eAeK3GS9di1mmYdizcN
l3F1BoSPnmIh0GOwRonaBi12tSqttNEJpTxXWvhyUDqE/3QpJTJq1mcpjKqfpRWLYcwAqbqp73H2
K1B34AjvBNB9BSoKKSTLexySMDK8U8CbegtUmPzS5f/GuYzia/zyqh/6v6kkWB38wtDcEn1/ms8v
HzynlwbtbuOVnlAmdBHXEDpzcEgiwKJDwT/oMmXw50sci1q6xqHMRloqsrxLK/yfSKaaHF/ryQgz
Pd2vI6QfUJQQz7yRJ1Avo6rrbjfrsnuHJPuF98EIIgMedXdK2qGRuYZ0MqL0icqONAACKD2YV1+H
29cRKGXfIZUz5B9fzTJiDEJ9LN/vcFMoIU9kYuGJV5qL0uzUrh1JJ9GU9zDWhixOZJD+45zMNX/F
56zsIrWzYFxWbNiapVLPtRk3yoM2Rk1dxhPKe9FdGAhHhde1IFedp256pSam4LRqDsKNmvOfsE2O
CmAeYqz2mLMuug4V1UkMuNENvMn0vdW8mnbYHxyukNdSsCzP3wlgumIv3IIPcd4nXLVqsmU6h+Xt
L6J9oCIUTEjwHsNGcmhzh/3wWN3hKM5mIEMMkTKyUBA2L5EqVSjTsjxRrADhR0LmjZl6Qsrnm8MU
bYxgMmUOzqN9uVAqPaS2nEN+SLxfEzN0sXsgLd0eE6AkcWeXkarEzxayb+7q4Nvypq+XqQ7t6kLK
HnZsobANLVDIn3RziuxTBVAyU/PGWAh2IMKTuQ8pTibhN5hj0QdE7exj41M6IoQ35421LD/aXLt8
WCUYJZ0RGkEIkqcZb1yjdCbGJxSfGapRuuy4V+a/XKqqppJV/iua57IsxVgHPhLxlZsNv7GR9ymk
+q3BTspHuIoyetDEiv72Xne6AmNbkYSinrYNENSRRsfvrQxGAATHluQzfANI5JfaMRKFallQXAfv
gVicFnQJeeqImGuVgSbE7QIuTpRyIg/Ly88Sv6+jOCFf6EFcxkhbeWUuAOk5DYiKfC8LEH7ydH0b
uk4FdoanfwGHsyP3ZlpjedUVplcslTHDwUjpFdFVcDPv2SaKqPPZqRk62xPBaVy3dKwzyEYNjrgd
zPCpbVz0ObE45/Hzfk9pfA734vlyO8oHLy83kHChKQyTxZY6j5Y67lkS1OUg8IlAPjSgSYfeDG0M
pVNyZEnbZfMgbxA78OJ9huu5j0Hy9X5YuxAC2BfGmncTjxOnpq/lFiLrm5OgKU7G4FvfQfTbfcif
b+M8NkrdCEsvwOWCE8XkAPT/RX9X11q8AUZTmSuQmke/4bD/KewXaj/iiJuWmjzUfVy++zPpEozD
B9VOfjEC+deRBUx2In+BdvQsQYmWSVQM66bV6DOolCuYPscbX8PD341irqP8NI+8GOyX4HZl1F2R
PoNsKxpodRFc20Cq9svvTDmhBKdpyV/4qWTEDJ6kBdFtlPRYWSufjH4JRAZFilKHds+4HEqXtBYN
YiYUVI0hF5n7eY3nRXAh7M1dtWJ+/EwcVgtLfdMnYUO6FkjuM5shFdJ+OOCfQDqPRMbaQrKZULra
mqq+AUWG8hM9HZLFwI7bpstP03lFEwYO102vc6/WTFEPNEQ65bAOAiuHXTCJ/+17Uz4KEdjlxGHs
HJAM/rb3XfLqmHxurI3Z/CrVsb0mFGhRhbtAztKOaxfw5A+YcxmqdbzMrCPL5CtRtCKdHqYQmdFb
FCUk5iytTpVdov1Rzm6jj2OFZ0KoUP9wQwWl2c2s0mO/Xe+aOHDWjqMPtxzuyzTsVdIowJ0G3SX/
Jx9Jw4PEuLgyjWdkIXqyAMO5G/ZG0dFBOrJquIrqAbfq+Tgl7KC6AmXHffruaNocPfwuS0yDmR47
xFutIkdKx44OK19oGW25Y3qLPBlbHYQwFhEstt6c1zDG6yboBFV/Qvb9AyezhVRLB9jAEwSG4T2D
qMljwpwo8nFlDAOvktpsfb7LmauGaU9mQQ0em50CLGDe4uUcjfT8tH3yf7CT7h7LdGH/5pFVyDiI
n5mDBDJDOg+SToWkksSteqYAu1OCSZN4DDgHAU1F3LvuXlb6sIg5rKAe/VgE2UdC+ZwqzVKAXOkc
zzUQSoS68mhSC/lxh+aHKJCV6S1nvDJn9OlcYQjf8Vg6Lxt4NcgGhvCiF9s0L2blYLdPEvcHtGVe
mcy18XmSYXsRgZID4WdtAyoHmQVY46yT/IbsE2l90KiaIlHAEp9sUZfeOEVw4k7mDXRKElflDHhr
4MwCvCRUbkTgYrFQXQqexjsSfYzVk/1VWijbR6C3I7Ya6q283fJGIFSkTM2nzXvgkjzHb7VUZqyd
bNf4SHO0xYJldV+aziTcUr3ycDLTVBbRddbFHMF55fHgVnmAwBEQ1YAkLSieVecXxyG6nKWcvPH6
NxiyEOqGkR0V8/veGsuRRPLCvHeR8k1CzL5DCqklj6maFp3TgpNBinVayZ1VRqhcQCE5CqzJoDQv
wrJX63Chdmvs03bI/tMwsp3sfylzVRAd8Dz5EsdN9x9uyyecBxMV2QFN94Q4nCfSStl+npw0h9pa
ZH9BWfUe65sa35oPmvoBEEvRY4jiDke/ECdQO9EpbU9SKGMiSHogFUsSyllsDHv5xkpw1pBkX40t
h6wNMvJvQKIBhYEQvSieLAwlvxVCJRbM9vHiZnwDG5LNLlZsC0EP74c7/l+rA1hzHKEU8J5XwzxS
5mFAnWIPHQydjExzkS88XM1ZL1ike5TrwHqvWjKIz3orvx/LvEZmcRbZkZrInO3/ralXTqZDkv53
TiWOY/nbR4U+uUPqI6JUveyn/EtOrVRUzd3PsVvhL9J/AE7tvMWZyGz28dEAYuq5NgePM/oapa6C
Swjss6LchE8puVtgNemQiUudiq9I7XtqtHk0RoVFzXTOUE03Qc1kKc/AsvKMWLNSBaAsL4BuCufW
bEXaatdGa6Kv9+P06c/35de1tlZ7t1CJpKCITIIHQH2z0FSlttPlLVdl0WHzsH499RXhzb/Kysef
VLP+V2I3WT8SXxVbrP+Lw028CHkw9yds1llTuOEXjfeMr1tB4qJ+2BNIJbhKOn/ZPmiU9HN2Pz+c
lOdvXMN/wV7MHUWnknxoQUb8bYsFSfFPd6qVJPFR+MhKEnYyy697v/RPrOPM/ngWvH5YOMV56dmc
vxFtA0Yr8TTR35BeZMiLLk6zdn8SAx8Vk0SvaxgW3cQOc7G4MhzbvgZ9R9hNiBWuvJtWIv+VTXwc
+GO9Kj3zcUf1fZZg6c1/3b13y2ifUlfd8r/IgjSWx4af5M8TQRud6eeWcOgJPPzEo+FXWxqdG+Vl
7Vtr1ngHx2Yco68lCTk7302UqOvRxybi6b2MHdDU9YIh86cHv0IKc1Wc7EqiEF0M9V6LPmwcv/rf
zbOoobcH1YWeccw7TGCGyGNgvtKp+yAQvzpLsShWroGOKX7yvJC7z9qME9/CJdvxLxAW324qfTpM
JuIexblCmWqyk4vfXZPRxRVv4fRWKMkCE1jmYm/bMMYQp9Ggj4NYc4qWtuTnPij2KK/1eHSbch25
1AlEdlWgSIJgw4hdlLkfRBKjWZL/+ytYhwVwsot0wLMRx8TaWGB6GEBM3LODdgnnpzfZGN5C2ajC
IVEsM+tzkG+ji29vdy1ik3sbpMx6Dbs73urTjNGNDpPVKAIQrytA2Zpc1wuU0TUA5hf5vg4tRf5a
1AENK+OZpJJypast4s/sUMDF6+VjNxXYcFsrdsP0Fqm4CW/caJriOXY9Y23Jo88htEH+2ROcXmCx
FXmAmgt7PLQEGXpvRGbSEvyoSFnlykvUXSJbhm/5zSqOv0dJ8BRXkjZew7RQVZoU1MXhgoMLVTZW
QF38gQ+/n3iItdTpW7a0RhXANeUiE9k/aBDNRlmQ3KF6zOQbgWjkQjFVUDWXsEqHcSrZHjByLjNp
miE5Cupy7p1tUtZmo1tYmYbfWTf/0KygCWS6bjQnPsK9YBaQps+b0YxJWoUSqKbQ8yWC9TNTmqFh
fI8rSESk66dKtvHtLPlq/sBJl0idE7+6iVFHsd9MaIDshzMNbSGP9YRMOwC3Bu5hELvuGY3W5rcY
ADfEvv792W0hatMY6OWlvsmH3nNW57yDyMdP60GYeOfU3IGM6Z3nuxc47DVoRJ4yrgKnDFKDXAvq
cTDSY2ZDtfAqocMmwNQiKCBaNKAXh4yUh6OSU5tJCXEB2mM5MuwZu9KZCPvZ5ezmbbTqtg0igrwa
CVg3F8DATI3bcKyXFHh6kMUWtb9oWzWbxjKbpN9KXXYqg1yTcfX9Cynt06Rac5UwCTXF5jAovEPr
PWvezPmk6vF0bv7EmF1O9rZfcAjngHskYC5S/L8NMqYQ0/CrDdRlXJ6x/x/Cgc/WMHrINKSLRcxn
DqfS07Q3EBww66OAWuPlgHYbK5hjRyG6A0J7brf7z/nAUpUYe5v5Ddz0nklLZVF+fqMvzM4u7Ntv
wnkXvNguCPz+V0wdmIuNPpNS90zYEkNOj/MdYYrCx2snqC3QHYj4ml0xBOOZfVXpB5mmxTJfbuKO
Nqfisusi/80kBlgOOcD65ucRW7wwVYYtksRAMGjV6uNv8gPETeqv5R7/O3f0vacCk8bodkk2mMSd
TSze5X/b0ivulUDpqczAJbXwj6YuYqnF/TW3sZPei+bv1kh3FkQS1EMTYzIRO6lhnvzj/Jtmq0uc
GbODBcUmfnGWdX97JhKqMirFufRVtIqRC9YSo9aeDgvuF2MK9qhCY7mEQ8biDD7VDdNOeZrm+qTL
75QMNOSpUq2HfxRPDhZdtHx8Q7pz0WCrHX5ldzK0YZB1cIM/mvrWZ+fd/rKlFTgDNxKQgM+UUbgq
opxJbmnO0c2B9MHgPtCcQ6UiHs326iVP1kUynT+8CLyVoYGkJt3GLIdTtbnGNLSR1++CFq4qpgvH
80XYfgP+PdOOV4e2+UxyMpa1XHl8Pas/C0DkAzqyA7WAxiVYzIFAOrJldbZh0/nm89HXMhhir8Qo
EdMSBor6eFKZEqVGRcB/OoEB88qOnljFF2Nl42Fy2mJIea80iuF23q6xsYeIm4eDXldHETF5QPML
VIFsdoKeDVYb9y23KxAcH52KceusETmDJBnhuVg+kuXZJimSprjPrEakwF6dt2fPeMX2o0k7zVtg
nqUiXxTIbiipw+jhSlsb/1Z0zSOJWGJrTv6yGGOO6ogAm8ofBkMPjD4K93CvaL5R4iBtiXxmwccM
omAgg96YVC+chB0Z6FZo552c7ckS8BiB5edwBrKft+Fz88xOMqWRxXpt15NXfTD9Evr6216KvH+x
Dg+S+qhv+w+NW6ZaVNvaH+AEdNdcqAUMNBr07YlrpZ6iAOkm+26D7g0pSkUt9Ef5M9N1LjYHax6/
FjqN8frYGSjTKpd2aJHsw/1kCWmaWr8GUsIUmOGF9kMjA2XhkSM6gG214vcFEm5Z3UA9+NoSXpB9
7WCmH1hUmrPgB0ZF5biVQ0FfW3keqni8avAFKDpQEsW06a2z3DpgYmuXR3/NNMIgl55kBFB6lM35
yAoryB9ZMXyWGuaELE/SLUkrMNZXozP78muzWlXtxyrGNP1ew9g5rf0nKMbVrXBpASb3511PdECr
u7qqbSvkERmABTtI8nqj5wDj7ia3zpfvV5XYrGD2FQZbqHhznzPjuX98FsoJTcPDZwYnE1ZzmB6Y
ydYMnjlijWq723N/ER+k8eJp+K2Pgd8b7R2A3ImVMX8z/AFO49OxBXFsScCFK+2ga6HOV7ypBxm5
hQu+h4yQCWdwnKnPFbLIN0TS9lvCiDI/YOAw1JJE+V6DKSgy0WNW0aD/JA+MUiOpttRlxRERwgTz
dMr0FIm1bFRrS7PG+uuyG+oCfkmLxXc8JJ6wtpmxHfMP273lsn8Yg5G0zmcEUFczKnt82mF7keWO
g/RoIUPLVc8gwAuCBLRQOjnHY2t7kklum2PyNgnpdX6Vn9QGUCk72X9+4r/URnfhSqqlAPWO0iPN
21iy80dCkadzS69M51N1xTqT+J9CqxyxvKxBix9RUi9wFvE3WsNWw04+x4ideh9P2DZms9J2v1Pf
PS3Espfs83k5tjYXu+3MWSMkDpyHRAPMFbiJ7z35213Db1eQWNPeYw0fnsCOcnGRaZpHXIVm8RJM
h3vfKYJEDy8AZsRVcxGXSshN9iBZqNfnPc4WCztNlLNtvaHj/dg1CMecxH3+7dVW8SqNWB8SnSFC
3qtp78WyhrPSrGIKh6d6Uwv2cIFNJ3cQ/lqtCLYSolY8YHOIllM7auvGpkVrkl5Tn3MkhiZjjyNE
rm731AU0CnDQooYot0yVeD1oUBSJSCLSK5dXYiG6pilFCA3mfR7Q9GFVgcpBVqdZBr8Iu+fh6AXT
6S/ufcqoYmnII5kni7/Y/pJkplBqJQhXCmIDQHDQPVH+7n4vAbA7+X4J8zUtwBfKNGFKzHEHCfZn
s9nRBHZF0f7sUBXmrtUFQ58krzDLyjdk5wzfltl4RTs786IWRvHdPJb6Z0p5vRYgI7IqsPce0oBW
wS5vgbIX0C8YMZIDjrHXWVr+b2R3uWyY0NvXbgrPt2BF+RBbs+DPLrs90NjKFaWf3P+SZOBfjQJH
6vFt3D6/Kv1xINGK8yq0ADGriCxnjiIkPGcAf9BW7JX6seIeROCuG2Gfdkq7BQVZDbJSkHJZCA2f
fg4WT9KsCGb8vj9Gxa/tK5cwYTvXOYkfa/SmP4wVXtr4QorA0fOmPDxumwqe8xyuT9EGbMCK9V5K
Juo1gXqDyNuOBN6/sc+IavH/OE1oaREEDNPH7XP/axnAY6czm2b/z0tqSWt2Io7sNVpEroxDPwC2
15S5zpiGNvV6ADc/jyB7LOJH/LBnctXcXE5XG9wCz5GT9+bAtHbTt9ccbtSE+a0AC/MHlrX4G/xR
C2t9/xbKJoMnojphFE29RZVnTvKQvDiVRBqP7LeN/9QdfscLC0V5oYRdlNhau9ssofL1BNPuaheG
otr+UG+Spgzn96mempXEJn3/5FYnjVu2Qk79CGyDnmlflEIrzeHGQQbjM9erlk6o1Y0M9ZRgdxoM
BCU1/fd5LHvU501v4UKv8yui13oGG23FeWQQ5C4Gfzq9/T2/XeanQtZfDh08d4Py1GzXD7TTIR6p
fIbdty1esobET2oc0TP45F8E4lvEv7OhEJGD6xRMOPF6LqvmqrXMAqNmo5IXjO+ZnkH6fT3spNVC
8EKHMSCZo69oFBTiE2rvnCovIcDWSjz+xzSbA1/+WrWVqQU0QwITDK8xAw6yHKCHrhG2977MT73d
c2F7ZQkPrxta3UzT5C/N4SXoViGklgyFEkCoqe00IYiZTVqS6jE9ubMO7LSD4974QRW4m++DxSYt
/HaivNvp98b3n8M+1ArrZTdhRcgsHQzTMO4r+UaeJgSekufPFMKEEV4g9LEc/P8XGHF3JgCs2cCW
S0ddFRBQ7iHAF2RBtK1tSPeYVIXzPbZw0qLLzVp4iiZMJ6JPfNxAPoimyWSzaXNapurn6mIMM+sV
6p0UdjMChjfQuI+k2L2AjVv/dorhnoF+UdQwnN1HxnUKb2YcvuzffS5gcKftuNdM9sJCsVHPq41G
UBcyPv/WgQ9O53gD1UQn7LU6i7yrvXxwXKc2lqqan4XgwpWZs8F/bX78Lpv0aZAPS/egRQHSnSJ5
gY7VxBIZsXmvWLh2CHTZ4tSMbi/tiabXIybFxohAyzbyVWD3SfuikZcbTKD5JClM79LPzJkTojh+
JQwcO90fWASEvRz4D0pTzThm2V+imMDvV2CFD4V9Q3aByhmI3DGOA+x1N8V95JzECEVJs05xVKGJ
1l8dSYT5j308Cl5qg98byEjP8PRq/oz3cJDtzSeG5KFlhw4pmQwKdg++06IQ+oK9FBP6cYkvtNsm
JW5wOb9Bx1vPJz05CdSM0z2zNFPXEg73G8tAsGiuQT9fNekAfm9dxt3vhRoBzHC8a0RtToBF+67q
Yv9Y3dWMNXWvE19AIneW/7BNAQNQ8mFL0Y2SGsnU8XVOHfiA0OV+KWXvucQ25noHG2AAkcGb5kv+
dFy9SBDFJQ9A7eJGkDkIoXSMwXe1KFtx2KsLw0O7fZ2gygtMWs6PMLrDDw8RA992fmzwNbPwBJIx
KF8FZLi1b1PBtBswikdteOC5JRTk7qoyl44xFNxnFLJolaEqBhdM3uwqrk2iJgXZe3MC0HScE8Dq
o+8BrB/kRRDsFe51xwT1Ue8MpWh1rOkPQnGOsdJVCQtdSP+4adBQJGubrk8jNnu0GPUmPv6gPHn7
/cEZ62yL/IqwQrABG+zTDg0vuip886Td8k3XnPgryuqxF2RbiAUMXogTiHBx8eVQQ+PfngCWeE6C
sx2UKox9CU+rqh6M2LHR2GejqFWbBHpMsfd6iyR8prazJHos+wz5GooTryxxfWV99IM4EPU+9RYS
jhqRQUiOSmoBL7jLSEJlXWMjdYTmNZeC+jni3NCgvrlg2tPKaGfhZMZGbraLwvM9QiAuhVIw71N0
MO4fVxzeKwXv2HuEtiACSjgVaj+q4qSMjgq5np03gY6DGMI0gNAtBEUrS91fqyKl5Cb+KORDi5vW
uvNYZjJfU8tUBiWHHte0wS3bJGw/CJnVT+J2VxPSf95HMFBS3iljifM079264VuXivgdVSWHaOXm
nLqI0W3MCTP2BQdvNJFifeoiSlJSV8Idi2G/aKdV6Dpu0cThqe6FGtPCLcgmdHu5sw1GDdVEswoU
vn5zpaefQAr0XYH2eJ18mJkZgpqktFTjRMZtNpLTYiAOj/dn53vIZ7NKe9dzK+iIQ42HGXaNbvHA
+xvav50swM3e23UDV0yx0NOjiDu9Inc27NUABoB6TjXPF5B8P0kwWZbl/I5/Tt/wMpV588ni/ZUq
m5eTYzWQhoFbxG1OUiZLTBMj3y2Vrqv1XBpfpCsXDdPjCDpzDx+SPEUWZXnvCBZLI2NOIHN61Szi
533I01ei6llsZnZk2ZroIKd7pW6kC5F6Yv+LUdvLg47avjdVAyjeamMaNYoOJcK8wNz8uaIa9aQT
f/bDDV7rJteudN/dQqygoHzvOaLDHdDyBKRhSe5oCz1i6IqhVDELqZ+cB0r3DjLGhm7HbBus+Vk7
iGTS1JxLqBYfrMSpgZMJe1U84iRDByJCi9xAtyvE7rDrDW2358tmb6FqqJ5n9hfteHK9yIz1xv2C
Sxm6ClM3ZY2pIfUok1hyLlF68Ejpi2tv1sFMYdxCKBj7RbL7ibevUofFIi6IniiS6X5Gj8L+fUh1
+vfvkf46rTE66ElHwanl8viIn7VPZ0ZTWCy9dYrN14RQBMgwPKvg4osUr+ESm3WEWUF5ZR0Mp9CZ
Qmv9w0OeKXt8AuaRDYEXzqh76DnOayfmkchjSLOUGUV5gy0n80TREztvHJNw1Sn3zwu2X0ufpI+g
0SWpOTfVX99k936tKOgNMKd1UFTCTESo23qgK0UB1ynAKQboO4BhrpmSNTu5xpMYVkFwhWSczsTu
a7bpjwisPNlR6s/AyJe0kKkl7fV92njTQQeEAlbrr58ld0tLCS6/Ob0ly+Mo9CDOBP8NyGucC+np
w6KsWI7+KsH6iB0We5+/N3ZorBOmm2rB5qX2rpJ13umqmU29TSLkM9sPhY1YQeMBLmo1YfIJXFZJ
zdsn9iRLCpav/3nTyBtLFPYvpQWl91Y/sm7Xy2IkX6A5BMwwbzeJJxPt4PXTkstizvJ+OVNy5BJR
CNG1RtT+1vMx4PcQlCefm5Si0p4Hplst7srop0FqmGArwa3RfPGmQepW3vXmv0qDemNvqoYUNf7K
ifFe9Yvk2JOPMLuwX6H7z47pnwDP5/tVB3y+PjaqviCbqJwhgJGlBxtx/3zc0Z+0z7B1SrvqeB6V
B0Ut3wON/XR21GStYiTnhmZVJ9CvJcHW670wDNGosMayuSqQJzsW0KBOAmHp1DrM+hh0gU0CXLSe
38VkRHkeiEDhvCpBcsqnkC/FgqBkASFpfwgxYGJ79nduWpdp7pWzzs/lgMBDNEzN+hqzPKgctytl
DWLB874SGRTtHA88roGBxTfFD++K6IwYDUkvM4Z440maUG/wtfk2BRHC8qRWzpa+YuLoeSSHahdt
25eYEZ8M6/mdTxY/6RQQcbN1t6tIvZ6H+KR7N7mtiwg2hn2sVEBQjZzSWpA8vadaFBBwzVPdffM7
bMQkZFw5XZo118p+rnXjWIwOc0CM4fc3Joj0A8PYRRK1NXKJSP9sW5H3CYu5+KPuD0bkVRuepoLZ
U34Xsm/BcRwZCBKTmSPwaEgoVkYiXDar7ezTA9iY2vLzL+C4965g9LixQvuOS5BdMTJY5pO2Oc6o
De8wyaBu7A5uaR/qZAD7kYqLQhlprf05sLJh3pwwnzdvn2LP2OYL0ojmnq9NesCigTdadbGKc0jc
D/SNGGAOipCwMOZAkEKLQPuutLmWmGIhKOl4FXBlBWb/oPFOLaZdiRkL9tpkYfwqnamZbfED53Av
ygCYyYRLs19EG+P0CVdrReElQVo55fBzhgerfFRmejEEb9A78KNNB8m0CKmCwH7fM9JmvDLPd6NE
5T81MiqwJC0BHW9l0rh6tIJoSsqNP5orzsr/X37A16S+1HlG3ChSJNkY/N2wGe7gKcb9n5MkqTjv
ArGVtIbOnXtFvOaogWkPQRIc3hHY3lGM/fqfWv8jT38SZMbMzjX17rot4XtHgtCQCjPgiwtRIprX
IKA7cKFSCtx15+zyf3IqQ2N4vHnzfVdYrcbpNup+R7VeACaUv8HLXIbaHAyxYwGEGrNixoHrP6d1
6KX590s7CwHNA/JCMauY0YuJ1D7WjlRCffd+LQnFknz/s5pUx9GB4JIzrE1qr7v3JAci5Tfslcuh
QWadyWf6c2eO/Bjq5CUd4Dz2K39KZjUkCpwYgRMS3vwJ8t7Jt00YLlRxcd3dNg5VTI5k2KwjntRb
lt65Wmt13V/+uGW9VW9yK7DlwLmnTfc1jKFJ5wOzC5kd4mFSlFsB8ewm/FO8kRy7sgM/qNmKE7cX
mKDIzsZGyEZYl25LW+4JytlCrh/a3VO9j/1xy0m+IcYZW8/AB+87/494GMYGtmL20P/T61XfSsp3
CFv75tSmjPvAptt+AZhX6l7aAIPiVym/Ijo1FdAeTRohbTD7xHTJxTiOFS2OCanoscm3l6wjtW/a
za10VLvNZJbejOqgu/hU7fGfxBLdtvDnweiriqNKFTKRMAX9v73dI9GCfphgU/PLxQvNx4REA8p0
F2u+vTJCjg+yNodvW+/rtBhcVEGOQDhz95QH3VBDVF0UCHTuuizrCdp4shyHed3ufFKvMjrIe66H
CMMEGltsNTTIXN57sg4yTZ1BJUJ/eRhZwI+q1dozINQDlszPwVxD08fMGYZ3Rd03Wy3rCnUujRW3
N+QT+5M0YIDfiAeUUqIP0IEvPEk2NJSfYRX/OBOUaAjliIMwjBFgUGplx5tffz4WIJu/yq+JaoKA
uUMK7bE9gW2i2JZs91G2azkvVDJ9BNN5C6pYjOxlOJuhVmSObZ3ghLXPS0Oe6f0DwddT/zWxVN8H
Iez+DlHoP0NuvN6VgBoNd9OgWQiB1sQCmKHLPT5vo/0AGAc52TV62pPlzHecP3pC3ejnFp+CIJYg
G0djdN6O5HFprG70vAC2Lwiuh2ZAcI0XN8YK0W947d6ARuu+iHLzIYdB4+wAN9qdzMbV/PXOwkZC
7PhLHONkvtg65VHU00apMMg6YZUTjm7MFLkLHaemXcKJP2GRsLMjom8mIWjfrXlW0qqQfSt21kDW
KRbTpyjv+e9n49k8yb9cA8yehG9pG4euLB03xuKqnnDoYGMm2UhJPFjigok2y66edAfnR+fISWtE
FIQVp+oAbIaEkSTVpsQqBnRHznxdkY0/CMprnPSDaQM20Hbf4GQHxlxOfKfmBiZDmmJkIkSFcj2e
MqRgtegLB+4dTaNHfOBQoAPDkYQjbrkORgHM/kg690r49KGrd3DtA1re4D0Xeq9fsR8609McRrZ4
uJMF1qKFveT2iASek3AkFBU/b2McUnIpz101qUmbPjIL13AoV93DOylYR+oT3W2KdRG5gU1yHDtl
UMCQEGtN4fw+47yWojTVm5KO69yI/dvA9f47WKtO4IGf1GR+Z820G7YMjuJkLzVqkwKUcrka3/Cz
dvcCoARa0cn05GGmBUVk/iWSX53sQMLj6dANI2Jg8CMrBjPWLIdlb417G50syI7Y0FRKjijBbE1b
tD9Di4MUOAllv7voe6GcYs5ADxdAhqj4QdxQS022BuRkzp9aCQ+8A8Vuzwj34ndakweV6WKDtcpE
CmBH6XDI7jhBx1WNCldPdJ52DCirLNXKxUAECPujrCra7+vyIpotE8NXX23Xy1G0JkYJbugfVjgy
xWSDISPKuJR4Ty7/+6tUzWfKZU4CIf8NdFpM91W+/kABHYSYfTmaRJS7fIHQPmi6OO8H75/KJclZ
mBCRYb1pOVTB0k07R/WnH2vY71ufCP1kV7Oq2VqzBVfNDYW2T4qlh1qQqvpmupD1+VhZrpT7tyws
sqv13UVFs+wwTs5BPhtFI+0KFYoKTDg/hNjCZwpZaENzcYBa9rSYNuF/+4jjI3aRp/7VMrfjQB6w
Zzs1LAQ9l0ety3LsWP448+aihXC+DT97W0c3a/VUHjrLILuDX2xHL8O495ueTYZ6UcTq1A9p2+Fq
hWGJYDWd0iwxUXe8OOuRFrnDWtsUpm9D1hrhtPWchnQdEN92EuGoOiMqkFQsMlRCUTJygag3kn2V
SDQcbq0SulfpotuA/z36agSlx+uvl8zo+omlw5xlqtmdDWkjwEGeKtvZ3DMCtkRnWwip1Ohm0ArL
8ONONbKgif0kjVqH2bvvl8/gPyrg0A97A6SMHVgjN5/sHkY137er7rgkkBb0H0yc+YLJUqM6pmPk
1gYYolbWPv5TXtZyER4CprU2ywEfapBuGCUZamNS4yDpVXh7HfT/GtGf/tBQmQlRPnJA2GOBOCNX
NNmqnywcTLn3JRp2GmbX1dFYkGZ1SuTIc7x0een6Yt/1keoa8/opVC8+kRQiirKl8wQkHV0LZU2h
7Pjpk4h9F7g4SV4dbrR4ovfRib252BbHN4G4hEe5momFWSsyOkPBlyCsOlZfS41W8MsBUd64y7Bo
YPQ5l1gy8EJgHWAFUBj20MgqyLlahfIRLznjseCzOAbQtYUTj0FdBPV9inIM2Q0O22fXWcjH0h2d
qyj9H9KlPEw/9yI6Xh5/UQaz6vVvg7wTq2BCrMTrFGk+A0EFBKmSsbAJ+eByYyhDgcRK6sDzXZsQ
aW2tG8Zo+yq1nql+HSpZk1cVQ+IO5jTfaiGxkXU1ifSoZ57+Ov70i+pVDRjJEMuFCdSp6cfI3co/
qSma8YmqIBANWYni/CDyP13c1HPmCTSgv8dR9PbanrQadmOe45S6UeGzT/dmOTj6gAhEncdaM7/T
GzoXQRja0fDKnToa+Kt+UrBZNKCn4BZHDKuWDWqnrDOLC1AU3hcreEeHmy50PXkEFvsyRVA2JPKz
8P6jZmNhlydrtyk1vl1t6Gtmcf0VZaoP5bd2QOwWNp4LMfGXj94V4XlEo7/9h0vH51jf933F9ExC
aVPglE2MNaihDJK6HImMyKtUI0se8Hx0Pf7DO5b5FQG+qARHX/vWdv2aZeMZ/TYEHnvoSWRAlmhd
T4Mf9BCh1xZhI+ixVLKZRxAiD+mFLtGaQzgC1XjowVSv2mrJ8SPM+yhE7rTFpFZVUvxFNskj/ch6
VhH5Yh8LMWGP6BPxM+rEwNQsPF2HfGqCFZQCS8iqWkbIYFv56GJF6jUrSFvCRcbxfWJzU6s4EGEO
EPdkyygGFU27rCAkGpJ/hGSHI8rF6EMNNnbKj3YwDEYaY9uHiIJed7SXvj0MfrpqjULSxRQ6G+tA
srIcWmpwpV8+mFlaQS7NbUcodL8PHGZLgeFlOxCT/WUk8vYFcqs5sUtp7CGjjxZdfcLoW+NCsNGb
DK9s6EfJ/3lLtt0jD2yto003EJSEYYFA1Yl94+rbHned7sD/TczZyfxxV9CMPE8+bPSUbtfKZQ7t
SilVQBNQBOKCgOEwQl1zYz/mSZeF+VIThsCW5obicQg/Qsi1XoIqMwLq4lWP2OBQpr3a6IQ+kmgi
i4200LzG6XDGwfhOK+0MG3Vv63SOFp+JyhT/OwDXg81cJe9s+MIGezTshddoMdyQ/MXoaUYyJv6q
Cn53t//bkkrtOpfbuHQEIHPakHdFRaCS9UhJn+kJknqs3QO5+e/dK5hK7h6biu1lffqLRg4OLMiT
vmLpJI4T3bQo8lHvZLETtWGBW4Lij9k2I6qRa6X6cmemEe2gx44AaXG3zC7H9pNvxlPNNR5NZ8fY
wtSlRZmhaddD8gGIkEib4OJUHseyh7WA3o+x4rTrASucapKmkWw6I+GK/wJpem+OYaxoaGoiU1UX
0Ophy68DHTs27mfF/iqhuGJtZiqvJh5zfvIdb9odHeDfZI8S6sIUkOV/ul7oVLydfOJQdtvnpnvc
+j9iOsS0aejEEpl/NjLJqzCenlYNYFW7f3+/kCUIaoxhXX+8OID09+bdLjY3Qi9BA5xKlZ7ejY7j
hC30HSQisHTih0gUpbm9JOuH3LFFGRM+ijFbgiBycHHZyUxHz6SXz9a4TyeAxhSNcKkDEzXonahB
dIhdBKavSrvOHriXFiIG2RgcW9tCPmweZ5kSnyYzO8U4tEREUILtknJ0/rvfmMGLBnTBuBtmeoIq
9LN6dFn9UQ599jj+GI6LBHHUt7Ja81b/gz2Mq1reImXIpivYPpRrauyXPs1U3AcZAtrpo5Y+Humr
ipi0zxl3ozgcfQ+6skalqSPPz3QKEj+2I3uLplCO7kN4MMXBb1fWkll/UrQCjY96rZOWlr1mlUcS
pf8HtmX3k6qw42IjV2uvyLmks2zydV5VjMqK4TdtTRTpQVlwdZGNEhg2KqW3zUH47/3dCWlCPZin
tq0C0hLiz/9JsbiCu+VerqOJ/n53q6fAGdXd05xFurpfz9Hna62641QsjCYJLS+Hw1UjKzshoNwY
KJdF+BORcO0O6L5aWi3f7N+y9f4I03eVoXGrW2a8KWvIfBLAT3paW71GdZWLSmQPRm5F3GVxEmot
6WDy/yJRrOARYjk181q9t/JvM5jtAyLjie99qcV9xMtNqHOmEeThTz0hloTYTikjxSd7Ql8lRzPN
jqsPeqzsll3HkiecXYBw9PWYpOvvQB470FjM+ausdBYPTkrZi881WItygv0WgPYhRv24s1DfTesM
kGY3KEFkX6KUdvEajOXAktdZVrXy+iOqnDhTYZmbuwcx/md1I+zymyb8gli6InWcoCKUURdfV1p+
OmBCDjUkzq0vvy01DjDwvq26dV2CMrCLayBDl3cTd1eW9ENlk2J4FiyI99peTEYAGlMRbzMdS8Di
InZGQw9WRL6oGpYXrVAyh3eBlYeAJwuUTaG84IobcCxWuaI/Dtz81zTlKgtEJtDB1B71Nc7hqeeh
6s+pn5tbTuTcBR3pZE2khkRTBx4K8/41OSuh/5UeeN9RoyRKxSJD+8SNSti+87xZrHdkLR0YBrDR
oOwWRrab1AJ3NDWhk9J2RHzloUUGqWjbBvuY6TJcXJlKtS95fYatGWhz92lrSGETaczo0QrBbJb1
taKB4jcXQDqnqNmVS3cnTITve8/W0Fp67owefwdyXBHPqv0qnlM9ZFJNkXKXx51Nqu2lL78hfKFt
G7KAiYtXk3JNOrLp+C+qa14+vMUZfVcDHf6XV2YEf9KRfUWUUEghE43QI2UpgPx2Eo5Swp9/yzdv
Mv91PtWitKktX1QI2p5FJgOE7u/usv6InEejLMQvO8SKCIxAXGUcMjmvRrqwfhQxDU0i6W4ZZGhk
WK3rUww6gG/w/BAWZUMGuUyFxxZWw8AsqlTyJPfwvzl9vevyXOd73Q6jptqRhftFj96lVO2sYWTi
mzyuWRKaAxggnwr93VgdTGKi6PVE6F4zz+M56uWeXzNK+wk9I7+zpFqFHOsBeQ7kkcdeNUs1fzIr
pn+3lpFXK++E/FIAyMZ/OjllTURF5zmH+4Zc1kJJWVgAxfvbK1R5/sjuLP6Nmde7xdk+qE+Goofx
JWfMzoZe9cD0Jg5tBLP88t4oFZVsIrujlO8IPm7T2qtDkafMxQOcnb0p/5SW+GfN8SAUlsOMwDSJ
Jd6xELKahRaQWdbISpbbOymbyzhlnKtzkV5JsjzI2Z7GYxJertGaTAMmRWIa4rk3WSwJal7GNrL9
CeDLhg/zTV0g5gH4YsDzJG1RwHWSkJwRRzEdgaPaJyYRXlv+g+rey9rqMA7zKqJ2o5eM0zwPqYds
rtiq7usx0kiWCtBrT0IGnQGQTs4POaVkEFJeXevvXD0XMPIKVFFaLerAP+XYHBwwrxXuvh8AM8xg
K9sozoOkSYsFhHMNsohh9Cv0nkIXmHANLI41fmWKxToX2y3DqDq8K5jiB1fbBx5W7K/vM2bHo+Ms
3aM4ME4QRvI2jaxPKx6/bN/zFZeewUXfKDp5j+ELRxkMQT290jWPHB/WPz192w9qFXlXubkghblA
QXXrKrRHoseHmNnVQ5FWtNGePdm8hvijF/5+Xcqv52eUekfxykFZIx7m6ddCc1Cb5otXKrCK9z6D
+5DM3L6Fvl1wWtC8eFdcC+nWFwp4/NwxSuv1ky4iMY88uQHIKwX9dH/f+qNoOCZj/z2MQvPMuPw4
ZbBmRFfjk21bcqvDItkpKe1FpmsDuWi7kp4dC6JQnjnSaVuzRcOvlPG1f0cPv1OGYw2FjPoBc03f
DT1OxPxtBjW6rHNZOd9Kyd68kdQ3vFNAO3lx+eH7W5BACv02Z54FtxS1Sedf6OMs9xy24NFdEhBK
hATNO8KbZNpuJ/UCWUHMiH0zbkVWZ66i/RGi8i4wnIBw/jcP86lAy5f47rA4Hip/v8yOA7BXfO0U
IFzQ6CaGyiPkwQAIjJpA70aRdGq+aeFgZh3la7UvOM2XHmRztgzqG7diDdD+4MIBm/sQ8iYw5299
EIIMuuogjp2XIUiRZFIEGltKX7+kBNqPAkzVBWgfyK4n7nMwuZHKQkplSjG87mcVjtR0sJgLy8Zl
PcK67T5zEKUJTKpj7kYCtnenah6D7IElUUdoR6gdoTSQLyP7I6meZA4mYHk89EBBki6I12c9vG5d
3dIXXQCawl8pRYw29UBMlA5+Mh6YftQ05/UxCiDf4WyLBnOuTPApLB1VWSblx2tOjsON8iW4H50M
GlvQWPB071/PTbUbgM7SMliPDjWp4C42vb3SOf1VC0B92kvg82s1lUE3rvByim17T9EzSEKztQSk
60nPJJfGy4K63V+Y1JXvRm77XuKS90i2BP+P+EGhWHPYIVjUCqKUmXhFUyJ19d6FJ9nZnMqjav5M
OqBeMmO8GEC2FjPaozBoWwjIj2AsrrfXiwFYGWJiX3iduRT62Wt5TJzayL7f0KGeGH1loraCx3Rw
jpgUKoC0qRjWMegzBFOXvktGNPBDpfZF/dqbSC/pDbgqJCmS39RbdenRbOXY7N05Ydwk7Jj+px4d
VGBscNKZmUeddb/ORCp+WgAQDAkbZaKavnL5ASBFpPzubT5HGnsdOigomHTKzdfGrMcs5UFyHeYr
bBvS7odXG9EYRlXyU71cifLy5dyu1bivOoQIJXQpguo6S7LlCzWGegCdVJbe24p2ySVJdRnuzAxK
z9ko5fh+peZs+lowNR8AscGhDh3K/8SN283KEYipyu0GafdgPy5Jldvo08J6vaOYcJAlf4R5aUWY
Ad9MH+Kc/q4ikS+ts+G22N3IvQ6CUu/mNlTn0m9gxE/jkqmLg81GONgagaTrUp7Nra30s/a0o6dl
IxO0JBOThy5QfAzI+M13bxfQAkgsLgckehxmX6pzdtLrAd/1cM8n4Ctggoi8OwCUuRTuH8/lJ+4J
tMzOeEHkR0SB1daHcC+UeaWuNAc521jcsEej3TbO5J/fzuNO9bBgNL31tON2miP4sYD11lq+5bX9
UkuoXvBPWVB35gvLAlf4+NlmIEKNb2ctunKDjrlGFZn2xttS+gvI2Vy+6LzONT67qJbrusECFK1J
7hwVJ4H/rwV1b7/RrSVnW/2Do6+W1GqeDBJ+1okJguFD3udjIYtCAEx1igCvjSnVSS7cAADW8uOG
rWBsWwxOnmUipWeRgivoLZx2xXn4wwPdud/rUrR0c6tZb0wveE3TLOpDO5vaDbcKNba3f+VXs698
ebt2si5MFL72P0pqxD0Jg9bNejvPeadNrEPMGSlzFZha45ZAMP4ee19xKUO0bv4kMPaUqEf9schH
as1VbfctA0Y1JlJ/TA/cGKMZURAcafjJq87e2tgODYmDD/5zj97Wk/Cv0VNNbnsaNUXf1i2ayqHD
TxkDO5OrSmUyDu6j4gu43/0HUramw8DLSXmXTxlZgRYY8qIbF3LWdjQpBXVgx8PpkY2qVYu9gm04
yyFt/Tf+1JdjXvXbUDGVYrBZJIfvIL0sHfaxSgGyNlvTA4yZONV/hy4zf6Yc43HZNYA4Sjz5draZ
hkQG/Szhx/ZUpTLmIHEt0Ee9WxygkuYXdfhzJUXpYI25wUobodyfgu3idClRBCKoU99y8GS9YiXA
pCFxvBeUIjbzWR7fUxYweWP6x+B1IPeX3m0x2xKy4J4EwRqCNaFBh0WG2LRTd9Sq7XyzUlHTH40w
o+y0XFH3lPRrxnc60ccD6u2V2Pw9bIuiQYUmWkV1iNzo12uBEr9rWSGZmmkuZ/o1L5mcgUWxUfRf
ZUFdGPMIoVznmTNm55wTlxNKe+nzfThuspQpQeiGDhijZAZ6QXTYnbgBufLV4R9DOnnEmRZ2AHLV
Y4Wyxh+iYTGMuvTKyHzvnRNG0t5idFii2K6gGbgLdG6Mt1tak/vG+h0VbsubOd4Cmie4DrtfrNDY
dX/7R+AI4e6u0P/3P8CPZZvAHgn7QgJD4NDQiUv1aEvJSgt59IKnl+684wuX6P0nOXrVKG90rItW
9gomZwkFxispM7gJcwd2zYNhXxTwf9aHvErFePNHsc3BZiWzjF7nw9Y0C/L1GiFyN4TgLs4CCF+a
TeYp+nd31FIHfHM8ADsnFz0LI/50izsWRQVbdOEz3oRuTGwRbl3EKx2EXKYM4/ZZewWTfpCWNVBf
uLspEfMYdkW7gYIDQtAXAGrR5dS9Q46iu9eEBmmN7LDhhlsAO1I0QD7S6+zUohboVMOe2ENBFlow
6YNm/JfEJbR+wesL/RgkI85LRh41drgHfYTKFR+2COuLAgIs619fZYU3akR9MPUrT0VIBJlFPrFN
onnNpqz4EdzfAxr+Tt/5DN0s7opMkT9hGL/hIiv4JdD1I9P0FUq4ckS905gFHk7T8q6SDzqVKhVn
/Wat/DNlhHeEmFreCr/bw3gceV0RAeS3lR37DBRYVKD1EFMwmXNOnZx9aKpokS1u8XC67LMXQxMz
N6nprJO0khhCGDIveKjb6xzHVK1tR5HBwjXxgg3PDstLyZlGmKS0wzsON5o10VO4IJrlPL8HbhsS
j/cv9NE/91ZdvbzVYchSV7TzD0yJQ6OOMvp4USjkbVXMGRRjvFqsYjTDGKcDP3KFKIGdGTMEeAdq
c6IgDncODk1BRfprf7yvAWeuECbL5J05tNsaQZyi2KaxiAJpsnXxx0GoSIWsohvbqwwZR6pZ2Eoq
a8N3ZgSdFXNtfPco/3QwWC4YR9RsNJHoOfNjYGDxNT/nsAwm2fiupIdOQKLPtqHjQvXY3mvNnuVR
x6UNjpzWpawTeDBvQDV/JzXmq5GBmQz3MBfV7po7l4UWbQZtSDyp/u/4eyNWmFRjyt/DmiO/Q0dX
YKf9TOG0z5g7EQy6hKnM9X91NUN/0+Ad8U4oHIPVIL7i7w2POYel2TnAjrBgU+mka2UrAQtgWpnJ
7ULIXJ6lB6zrjyCb62okJOK3n/64rnEvRICVulbs752CsI6c9qAVNHJsQRcWRMyzWTGC48CxR7/6
F+TXV3WA9LS3IP9aZJOsMsBJ+ZSACEIFInC1p3rV1bzqDoDCXjPL8MFF45dwrZ+cnMKkm/tSAQfq
rYOiq9XQ8TAt0nF1fcoR457SKWYQwHiqR7UFdAOikcsw+UhYaYExmJlji+g/bO09nzEg5k1Pmdex
Pr+TEnB/7Et64mggZYyjbH7jjuH3GKslTmDQRrv7IOICw/GTjzdBY9yzghs8ZAgiJt3vvUSyJa1F
swot3rvlKRgKdWA2xB9esh3H/cSsVWOnzm9FVyZ50ZH5pE/8cRq+rTe0NFdUNl8Gyh5ZBHBNXzDg
GXwgP1lVA7uFOaGnf6NeV404gNkbullCaHLGzMb/I1IBXGEVMsLUBEpYpp+/BVyO+i7PWk1XkQfj
vYxMYUETa2x/GMbNhNfua6CauMnmP1puCXKMoc/6onznsEH9E3tGYtmSROLg7FllaTY45AaAlDub
qdC5xNKycPwYdYI+dLDHk+BlHz1SQFHHVVzdoMzOnE1qn+Kh196k0iaheZYuqDIdDCPjNopDZntz
i1Y7NijKBdh5Ojut1M0gRx/2KKLilNMgTKKVRqKkT03TLtEvLkZzqZ56P0EbBF2fkD2BzgpMjXiZ
5RViEn/KG6Ih16Y4TxkyxQ6Dckf/oooRV5esvMIN8//bXq8MwiLJZBsNR80rn3rkadoFW+RzQRqp
YBjKEDHE8V2Q/RYRx6Z3SAX7uP3wTP3NF1UB/vJ3RvyPq5RFsgpOTrldR59GBxgTFDKwCtvBVec+
0ujVNbfsiQhTY1EGmpYv6GgaJJ96PcBNYKjy9dbsaCwrQJPmQLo9PbsG0NRjwz1SKVDWBuLXKePR
DD79KX63ALsgOTzgPzTLp/x8xt0JMy29VMFsbQKj9jmQ1EERAyYVqMB8fdFKaezmCTpifqGMOrY+
AqIi0Sj2ItFrMT1tEqhyYe6vPW5sLHQsJHEeUAnBb/m40Y4Qr4oCXu3j58H/xbfwHIlwyJEeegal
lWZUtOBD82fYXGtKyX2+EbgAb9AsQLvcr921zIzcdQoRHD84pNLJqfdJaa6bLEIzJAC5tyI30EkW
sdo7U+m8WfsMhSWB67aT002yYFtlpbPzRoK/2vJdXjIOzzwSE53gH/ITy2FKCu3JzrLTni755/k/
7MB1oGWNI9OKQzEPITRtf/Cl325FMA5XmEj1w+9kO1mdiDztu/xmRnhJmclRdIgM+8MMDMmvMoIW
82kd90MnyqUDeO4Jztuvpq+/qfxGvc0e5eO1KcYayMEKeFxvuPAK2hIlsZL6JJkYdzWZrZg2kgfi
35VV4iQQLvq3J7GI4NJlkwD6t1Pn75XoKBvC62O9CGSelD8OysKvX5gQzQXG1BD02vRo3/lqk/nn
MDTOmrWhC7bks5aeDyw4fDsJvlxBAjt+Dq+V8T7jt75IiBZnHAq5YpdTnACjrnWl53ieo6hbqaxx
DRUgjABMQX643wH2PM2vo/FmJsG71fl7KcPojsWxSZU1rZ2HgI8hBhDyeHJlJzJrZzPejOJ4xO3j
CMMb9RZAxMTFMWMGuOO2MOs4HCAIgLvJj8e4oJqNCeIABQk8XHrGjvJukcjfPbDsprAEzm2WSWM1
bvlx9sr3CzbDfFYDUP8C8E/IPs2V+t7ZCqqI6z5x/tkMlGZE5VI00Fv3vUWHmDjLnscMooH+QwJ4
DvRqc/vtpKLtSfoYolxsx9Ar8gEtutWCiFV5dUfbtfyfgSmtBp6awlw96tiZF9cVKUcQ3Ti+1A84
Kfcf818PSoUbkgjbTfjMH9BfLTc3LGYWOI4ef1vmU0Q1IHpC6oxKitDmV68SXVmWnERK61sgTRbg
syuwtwq0xWKnzXOOyoW4JYAXDIpaS6mwIXRB2IZOeT+jjoRPcCPdE9sQmegGxDOh91UxXS/ANk0S
za9iNhngeZF8+sYSsRarjf1JVofCayb9L+Ypw94w6dtojlcPKAh+YBjNYJounHM10zY8uavM9OO6
Ikf092jlx6MZOHagnlMWVaXLaWFAUk9kvN9ORAhGDf4DmYfCFt6ZWlbvHdo+xsyCpANOlmlodSa+
svt/r1C2ODJdD/m6pJgT9Ggk0zCwuynI4iQAlvfRBLVVdncprPuKh3Qt+PX56yjlJBrNzA9eVYyT
9s66QTtT8CJRgG6qhx47Or3kvKqZ0WU0PMivofxpUJCLSCq0ZP3hVWLnPnNv0WKs5AgGoI9zQPqf
vCRmvJnfD9KJ5r+tr65K2USXq6yWgZJWM/UWUugWuXFASsfY9gTIOlwmhFUMh1tmdBPMNywxS36y
Faoaq2N3XRuVs2uIvXK93GlYl8qG3fEv9oGbXwn7BX24XLJIIHxwMkLutQSAKgX0oQN3nSQCJdxB
5VE+tGE267cqaN+4mwHO/7Eun7e52WGpbSCDly3JHtWBWgI6TN68IVL4nffULgTP8DxLpF5XCk5b
G73EUPSHsyIKxBWTYWvyNHuQ4rtMuUsmL7ffH1ZlmWlaNuFsnRvgsxYNP2A2e1IZ34DZXuxucZjT
hmrWGcgDPpoq0CuhdXkwr5iq3YukPz9rnxd/QOTsU7c1SwVrQdOGHXBooKf0kVH2QF2mZaEDXbUT
umO1ZOasj4fxiR0Sm9MrFqbX4MoPSvRcVFCgvcHcS4nvvW0kN0cx6buifi0tcVg8777C1htrzmbG
ho1HKXa+wsNOgqnz4gqrFwGKA0tSeE229MsME18kMJO2yHM7vMlCwsRXJLvhOF/bU7q4HMuPieYa
hSJpZ5cKYVdxZmIwh3mF6uDs18uiwJGAobTjy+XAuepyZa3Nfn6WC7zqnj4gecD/Um/TOI2ve2v4
oo3NpH9H109ZLVNtkVRnoj+mTrhWehE1oRkuGkwvNrtrBFwM4f7vSDE3Un67iuaGxE7yi9z+DSaB
fXFBJUm7wK/CF5D+CU2GVTUfgs+Q/LXNr3DmhlRd8ud21EPuTwcri55Y4gE+aC5lWte94pvun2Bs
l843bD8mZHTPKF72KkOke7cwSwas2m6AGQxU3hwm6X3eXwxIUKAfAcufvcyexCelZ8lAZZf4ktRj
TUs1ebpgFLn5APQl6KDvxJ9V8DZf5xAjj1GjovwfxpafSdIWkniWDYKQ5kOA9w8Ig3IhRTxmKIbr
z0BKSBVTPmePLAWkJW0u7qRTfYFoRtVlP2kqiuIjr29G7SJkboK5OPCI9zssfl+k5pP+U3gQte+9
d6cBAGRFqPPG+koKJREoQMxJn7LbGulTwxejl5ZN2aEtVHrSZ0hLSbNkYcpYcC30REfyuulRfLr+
8ABznFH4QdnoFOPmlSL1fIBH+cEVj6QjtVPXieVPGI8GY+hJvCeiAiUO25iGEC+uEdjldW/qr8jA
0Mm2G5xcg8hpQsvn/VcmTxv0yQPnMZfP9XGpmB3f9gb+H2bjJz6RofMZSTMTQ3WIlcQHbwqybV5J
ETI8ZKBL8r5Kr8vHrcW7qBxMvSFJy97jlwAE0R312YDy3V2jYbqpXKtIUUUpXgIqCX6daPRfhVO6
vFdp6yrkj7UI/pNQL5h4SzTSMU9TGnuGRojMZKma1/LBDyJtXCRUph0TyQbq0hP9SL/2uirOerXo
BfXiwO5hel+w8b3xK4PPGu0IQs1PB+IobpJESUyO9N1RWlrc/KEajFoOpYGpjJPYwAm3EixdSRsm
WTxMY3qlb5m6Uint37I3RTKitS76Dk0wQNqiNJofnaefKcg7PNOcdBrfHpgVRHemUuAmtDnKlrZg
Bx4adK87Oei5YkYPsJB7Ad2LmzfHAZUT5+M6sjMANOYsezMx3RDj8DJCkaKXfa5ekjwxd0kn9f0Y
3tB5EfzlS0kL4Y5jnzTW9+m+pUQvNCz/S9fMfLK94b4tEGuAV454kFs+4G18wrDLFIsI19bVlaL9
vY6srdcFg8ExdWIAGC+MUzvGok8MP6mAYq8bPBGEePzrvgakrALanMHx+pIqvRHptm5ifl5KOjeN
CfzJ45ZZ8xzuKMNJKdZ8opGaOuOwwZ6ymPjfSDNIKU7ID2o7YmYW6JT47rnliVeH3nL2Pzs7dunI
igzVPTT1D4msZF/ceiudkOu3g71TN510l22Zn4Eo21+DS9h9ZP/qEmKXhnILMzcWEaKVLc3nrNd6
C+glZqA3/EJJXtLI5QIkZp96TTZqSGXSNGquEXYl5BYuzqn7G/ssPZuQBUbHsqyG4a9Vy5ccNl7/
CTQU31/1stSyR6lN9FXT2xyjVj5SMjQAuL0dOAeSm/JcCdAK9sg9+yeOAIXTBRMY6XVXpC1UY1qZ
F+lvZ02EvchomSpybGZXzLhCVDU7pIIi24ISick52gUFmlwQ6YH3b4kFVS5XMU2KOeigh2ebb1pM
k00FSTNUhljwx3KvawnohCy/wYRi+Oauy77gJSM4qRP3lmdlHWylGGQ738qwnX22xX/cVgcBeCso
uXzG15EG6TJPxlugaK4PO24KQpyW7OySsT7cs3LTP23NWZeaORkgtT4o2kDC9nXEfHF/55+wBH6e
JvxfBiJm9xB/+fRsACUPccAXmqr6xzc7FuS/pnLNw4YWB7aFDKoz4Lh1YEbtO53VN4Mwc8Rd/2Ms
iTY1bIvj6dMnwRYdP4V2iwSHdEnkJ+5wA0e58XUiuzpd8ZDhDfyDYpOrt7DGoxbQVHKrxoc0nTvU
ifGcrOJbgXUeKjPhkdKLGd37nFCdDdheSyIrmrSx6TDhBQ1oYdo4XGbL+XMbwaeGjHL3gFeqYioY
ZxVsaoiGiKdMjrOShxoo7EfAgTAD+cZOCDllgOQK14BgqbX5b2TRDPuZpS5umJjQ5/850G4GoY3Z
JQ4hgdnEW64yv9L+JYpujg5AviqaCF+uVO1Fr/1yQu1ARb7MbWHTBKHYwJoNR7/+c+0V3cFcV7nw
eO9syYFCJfrEl+6s/UibpSc/Z7MZKz0O4cTq9GxU3IsTFMLp5nAF0930Rh8E0gCv66aaJDK+hNEL
mCZw+zAPeyISZvV24ZyZ06AeGEZx+Ki1dkX7xCcboxLeAF/zb/7TS/nA8l88mgTxC3sSt17OqtQn
EFNT/vHYQeQFQxFanRQlTwQObQXLgKYrKH3BI14iUihJNfunxWael9pqEGqSE2oWtTUWfpcmZNxy
TtWAw+IRnUh+LJKSoBfjMD5VwMUkwI80ibYkCkp8rOaZJPDOpDMaBavSTA5Z06HyCDRFFmDZwbYj
nP1CKymPn/+by/uYpYIyx79XYNSDRP0bu+QouPWxnPoXxdn6Rwq1DkXdUfD2MwgUYVLAFSTkou4Y
cVCHX/SGyhgst9PkxxFTd9unJHh5GD0HLKTEOM2gL6j6KURDZLWubanOibBqPQisesqtPbIekz/5
BNmat1Q6BJgA1HmWQ6Qshw3zMRFUCDikSmGlnOA8QIWgOfoLGYh9kHRsszCYOiiyedP4tlW0XI/2
Raks7H+gmIG3F0qLA0BEcWx0OS/goP+LkuRDj6w5PP7tAWZ/fub52VYcxcUm9VYSae0Wb/y1UMQL
Ezun7nH4X+r3v4YeYMSmphvCyr8gIRH/ISTreqqRZxFSusnfiQAppkqfujKSHnHj8ar5bLCheSKT
RHMn6rsFaYal3YuluUeGxYCZu4wsYFjxgl0Ki4+6d5IjV22lcyKTBTlb0PBS8Nd3ciALvy0JDqCn
UBXJpzizxrt4TFOf4cUGESGpdGxPSUvKhArWQk7IBSUG8+9qAWmSUlXeZv4qo1+67N3FGnkzXuLg
TVATmYSvhuSdqU6uV7MmTQKebQ3c2ghSy8IV7eTW603RzSDWzhDNkOHvQMs8g81VaRvopeY5prKp
v4uGc0TqSif5M64JmIMihs8aL7tKr0bxzYHQVEIvD6Rc0hSgh6VhUebrEsuItERyXyzZRIJYy9pn
+V9bEaIe2IDxIZwSuAmBFuCWfRzhfrNd6iTVEJwlccHQ9xfzjTwV+zkLf8j33IaSP+yM7lcBszcV
vyF+51Z8T/YsvGSeQRbgylgeAazOZbT5UbIWaTU+l+O9f2JLkZbeoOGQs5qGxdY8+azN7cftCPvk
WjnN7+ylxh25Nbs/upvv8Yat3yh/8/jfWaNLFpLBkVCr5RkdFf5BEH5zeY57IDFbSZSR0Inhqtk/
WBf3P6FUqzXDPPPuFhbUhGzRT5OMtl1hh8tyDVoXMi6bbF/OtLhKxmEXk9U8pkWGIZjeBiaVkINj
0yJUy4udnYoaXC8U1dZGF5NDxEcowqkblwB89nwvdw03OVOABbzzdkQojN64Wrt6VCsbnxGfuLRr
3wMxRGB75tOJ3c6+4Lr8bDpTrHFhPvFVha9zHvPIJ3c7z9QVx2DrZh+C0w3yBQUHS4CMdJPWnlld
IN2onUYGRvChtnJ45jlxI0gOgZnHKRRXJPe9fZSDbmqd2gl8RrTb9QqIB1ZoJ3ewihes9qLANvFV
P9H3FCMKkfWltekFTe1OHDuMDykTXRNR8O7SHm6jxcKiicWMakChyM/LlMK9wFjtxPiNs9rdSjGV
EKodrgZdiaMgV0OFttRaXqAA/oW+NRtFyT8CxoYQf36engt6ysJ19dZSvjQzm3dgMbHwo6MDTkIU
+x2qXpqbrCCaJ1sylD4M6cMZInk5IeExLI299IMCKkw1l0eCKpJ25wMU5H4gaB83q3BqQ/iSZ/l7
oVwe1s+3fpBtNTX1m+QvhaN+1qukKlA7MUH7KHIbj9ZJTLWSmF9RXfCT/7qx2UEXRlZ+PboGm/AH
SWmHIGLub1SxTay/WXQMc2NWZyX5zyLgwvQgH2X2akJkuek4gNnt03vau0FGbDSdZJZM3ICBkDk2
lR93P/R/ZOK8xsD9mXi2o7xrZiVtIKRiC9+mJSQblZSgetiQMV7411XG9WbEjsjt3T07Oj1wjMgB
vYUuJcrigNL359K566hCT9r9cJj8TsZz8Sy3RePIqmwORYbBmriCsDdHxi3nVpXIuA5cdFR4RYjP
tqBgBYDC/RFl/6BhbpiADlqcUsjsHT5W6jfKojxvfDcSoeAL3+YZ8KLYeUpe0KOkfZD28hIx1Hh7
9vyR5AIG12Vqm360O/6tyFEkH0l4UxcMLVPqIsjNg91u69dzDTn20epftTJIEDDprOKs3DKnvab3
teU7Uz/4c+XTFacFQJU4/o1WjCHxiOaA279Tjiu3WScXWari3OXNIILT5UYJ9kTRCeAJHQIw8qd+
CcSbr1/90PF30jk1fB2B57fuNnaTrdnCtvTlH/KQvlJEgJ9JyzcQCof4F8siMRpikbGzwpfDlIXY
vNmrQY6gbkIJ0/jfoclsTgt/IV4anpJK9YDiTBkEmGRQRctai+XXiZCtHY0xhThq/49IId58Wd7A
+nRzOgiVMLmloGrs71q/aTh+qfunVpLSBGKAK7n67sxNjTcUjJ8IEMnftchnpsJ7a4Zx75fLHdts
ojrjjS2JVwBql8+dQil0jnkXHzeLPWc1nB4qSku2wLV/N+jZsZR/ZtWRAe1YQ+UAdOvYqZdiJTtt
LezFkBiAReZjas6aNL9raaOcRrG6lFyXp08LTraSdSbvoUYTBc3ZoZwF8rxxQYZZjU5qleN/l2uO
A8LZ5d+9UtnGEAiKeUZwESAs8As6cYSxE2SgSJBAf9Qs6W9cgp3q59f/WFGbHnpaKHJQIj9yPxot
XMXSZpwYAAIiHvSs9Q39qUerQ9pOe9F87zAXnEkpk4J39Zy2q3MqlBFLH8niZZ+swuHC/Y5Q20mO
ppDUAyc6fs8pS8ExDrqAAYb+teBVzfXEzRPzQuEo7P8Y7700OYXI/bJATq7ilarxBmJQ1GqPrMwa
1YvS0mq7oMxNzJY982n6eSzEkXYIOC80/axcYgXFiV5TtxocKNiHli7E18FCK3hnbkkda/qRZ0hx
/FCeMLQjpgPCFeKlcSIHRBgcxZ0eOoJccj3D+bpaNBW6bm11BUc7RG/6zalActIUX5Vw6RBrH2sW
HPYT5TWjHknrwdlJ3YX8bqqJo2mp0OtRbmvFE+JSbT1Vet8C9cEcKZysw8GakokXXQf6p1lzHv6g
qlz3Of/9gLLpo/Pp/S5hNKwzCSj4tFfbvhXlQeBnHrpJmHAuS1+5VIe22EmgX4ABhcrY0xAmshAA
s8Yn6BXETFNOSGzVHczBL0H/BrJQDPUapDeT5WFsBedNQXA+z8xG3bzYXLcjBnx0DUxL536KXZ9e
AJve5Y/qKCqUTVCW9rtRo+SE3rWFRPKacnNzr7AzsnTaBHVJXdfcP4gd+0I9Nl6JkjxPvNOH22Bf
YKGR0TqyV8sdtxhMFES+pxlTQE7it/a8ZzP/IJixGl9+3HpNGDhKjnTA1abRasDXqnmK8y0vvuMQ
kRGhuaHT9w1f0PRysFgOYcjjODCXPw7YafhRnLZU6PJVayMASEGDlwAsCtQ9oRYqIemzw/KBbtDI
LpZLZLkuDluGoA54vy+2jBtCi8uYOWJQs3akujzDXuPkkhgyDSp74R0D/EdC0ivWnCpBX1zFAhPf
Em9PDV2mjL7Pw6hXA5tDqlPFa6HeM5CO28KnHeKrWCkKtQyTjAoSF0YqHGcY1OfvFCILmN0eQtS+
cgo68wJCUkARqcagBf7P4oMR2LHQqqvOaCpSW8nr2Rp6xsMEVtYAqaQbw9lB/S29h1jU8gcy2vjE
lmUdqWc9mIygCOKOQV6RTi0NogCwCKLxKAVF07kiGbo4lA8I8zj9VvDiOf/xaBB4WuCIOakHANB2
gPnbj0P2IoPY5XS6HIDuSdi0cuORXoScTfqA9M02v7h7bHNpLZVEkfaxCjJy0pM/mT99uiAYZODU
5slT+uRjZpD7OAEmaDlsBAoUsoWqwahMZrcr6wjoUZ5OyF1a0wqqPZPlcs8Fk9AUs9ECpv4HS1s2
rIkvTNf8KAqhSr1fxKgTrLG+pnPJIa60q+y4geTZ7ydJYLSlNfRPiHOoVDma9x/ZStqHoNqVj4uO
JKCtKul6Ob+ii0AbaL34/KZERxCG/cXUg0P2iRqpYnoBHcV5n9XuMGn4fjdcLXNHoDXGYvmGudXw
dk6++DnXNi2z8cz45RK5lD/yDaSXpJTEWeJ5YpF26/S4bPUKF3LLt7AdOhW5cUlb+ZQi2p3cQnsE
Ri2XveXl0fFn/2JSX+FGxEE8ujzRojZWkEENRLlrKUylJnhHKwQhM48amMYQXhfiV/13g9o6ZAj5
95EHevJSSURR+y6RICImJbSfuSW4EdqMSm7Y67Bj9uyUdlurRmNU3drLJQFkW3UTMMcqwTjZ183F
NMVvhXQVA0tsCSUoRrJqU203th32rwQct0miXeNf/aR8ZpDUPJ/RQvSS4vOXjKEhw8dyhmK2MLBX
60bwZZi8zBUU74lDJylsicIWGok8Qt67oEDJ2UVPN8yqHVV3yi8o8iiNFaVEpjVY79FRk6RgK+21
Og1Wv3YtxGhrO1twvUhTioU9g+SDDP/Q1gdut1cWmN6SV7VhTZ5iid2Bq8VzVR6Gpq7tCeJ9cn0b
STkotk1z8zNZI8cmyyPtnA0dl/jvB61WUOWNZ2l8P7Ljls5w0hyPXqzxFOGWStL05N+vOgL1Nwic
t0dYlw00opoQ41/bQn1B1DF5TQV9PcGv2c61XQ+RLIvOZNY8n/OV5oEOpnUxbSBTCkOmiaL2g8B0
Di0GxRcg3c64Qhy09O2Y0FN7FItzjRa84YNjkjbGm9kdqYbmuJXhOtLpu9zLTpLRvjVhf1Q0sqQ2
PDr4pKKLaUXPKCotM4ewHwivpKCS6rjmhmbXmoaTH8/PhjcA/UpI28EipocgFHCJ8lkOXgoar+/A
aGxAdveElLDs7Bv3SNVpsf8XvHDl7IBmNs0TeVvLzUrR13Mp3kasz1P9sMT1c6lY+hGhlfxJzjAX
iLPJIyeBLEKihi20V5aphp1IrtT6HCT5cG7s8eQRDG0Vjo5ElY5gKGt2fmqLx9zQuSxY9T7mtkAi
5pYP7uCCW8SsuInXBGldZelAFLwYmJjEnx5ZO6OAH/snEdxa3sHGULjU74xRGODLNwnPvU7BHyZT
zQTBsrHys4/K8AQOYMXi6Vhdm49ZmvN3zF2LeLCGqkH6lZHQmuLESL4U+n7PbF1YOqHgs6nZgh/F
NLlpwitghG8LZjWmc/hhV+bT3f3DxJ6vZnGqLSMxX4ga2om67xroka6K9z9aK9vYcKuv1vTVvlr5
8gY7pXOlcql2dd4L/0Z28swj0sMfNV7wZtrl5TsQcayhMl3rq9bhEnQARXlQQCqoHceEKXPoU61C
X/FolARVdaPYJce3d8ohuraw0D0ZurQONs/05nOSg37P29ZTcFoL3XQe7a2L33GQlfI+FM7cEogF
IRw7xXvnr/XeZZwFb4C6N6t1AJIiSYzaTYry77rTClGt8OMjb951XNTEav22CrTwzdO7DqoQp997
n0y6P1bGN9FxQgY2Ub74GMK6yX0UQa+QBAtqMgla1ovs+kaxedl7rKxy3eFufwUKEx/famJqOfne
7C6nlfrYA8/8MxW26DE7fqZEgbKORRAfgTRqNkjpf9gYXgvAYP7dDAO2ZQfH51esXrqz++DgmAEQ
e+qDNo+xW6qcwsms7arwZH4Jcf7Bp9/AkZEXMoobtc0hWDCXiI1P+g0TQZjvltdwruzjMp1W2CDj
k4yTJPl65e5cLNVNTSkLkTQ8hEXhfOmKHxoU82K9z1yfNyfCgLI/ARMYLC85FXE96l5NoPpoPUAX
B9n12+Q/wTupt9tnwjqRl4MEHNEv6imgZyWn/gipWDkWH1crdU5klNYThiCaaXL+MfFDjBdAGUlF
OcyTAQLlW5N0p56myKyK51lU0jFIFBmm1ErrlvRY3g4ekmKzihicMBEdo0Tx+o3uNjD9kNGYq0oo
3ztKU5RKIIlAPTbnD/Co5vPTx7nyt7Oq52tIV80ntmY8N9l3O9226o277wbrwy9DPaii68bAgU53
5N/JRWreFV+rmL+raB1Z8OHXdJ4FnkpGAGOtDMnO6OA9KIAVCL9ElGr5WO/JzmOEk+gxlPjw9n4y
hO4Wydy8M2jcP+VIMMoaKDoUTE0EKmX3+kr+BSGj7YqzSyK7V0K5rSWwVAu9BuRB3azv1wyOK7zd
25S//PqlxgeAAHU8F+7fhZWvwxlx5RJh4qGy8OTEv/i4SWKaFEVk+xJc6CI0n3KzD2gmVVaocOXT
rMdgwW6g+sFW4B6kR2wehh/klimCpRaPKBxi1vhdMH5azH9AkTQLNeC1hRVc93M8x5yW0cfa5ilp
worjwQ9z+QxOiI1vSfzi9l/7enbjaVyIWXrE7lO2TG016fv3qAXrOdRJfJRdewcrrXNUWL572a3b
4V+AMVPieLissJUUp30na/tffWdtXlCWfNs05EMdz78lp8HjQEb5nei8QowP9XsgM1F7fNnJCGNr
Cni5LwH1QCIIKhTvOBXfwzRMclcevSXNOYjFvLHoiFVv2s+b4vfjpny1+Brabsnk5yE0F3SDhhQg
ZbN+B749wwTw8O6QlxN4xI2pbfEBf6Bu3ONOa8sLU2P+DK8giCDZzXZacnHRmtQ54dY6WqCea2lA
hkQF9W81aCxcflBVckfjZmxURmX/4DPixZAOca3A9nQ9A4X9pBIXKdKQbniT8htZEB1sKmLZAh7j
hoPe+UV1wcQRVaZzF/junDjLI/tpnq+FUohuNco5nIurbYHr+ER5v5AlSmqKlAxQc8hGd43n0Fxc
GVnXr4E7YufCHUSLjhXlonxfJXMoG8WgdkkqDvGhAsJkPHEDrrlrgtmm8Ly4bFedwoA/D3L9GYQx
mVvXc5IUpkDrapnhtNHVyiBQl9EOUG99vKqBxotd2Ak2G3Xwvflg0saM9w4dM0s4IJAgsUqUwbZB
8LA/NWu7WEjdf8BjMzUcth2OY4NFHdr4LK7kRgp6CWfVlhCs9DVKRuggIDDW+UpKOfc84kj4Zd4l
XUVNnXMudhXY1PvTMkWK6LiS6J5RynuN2G4HRDr/X2t4o2GVQm9KZBqrfr5xoy2hATZraJ1Ev1AN
bOUsBx7aikdcbkIpFyUaqrSvd8en2/RZoGwr733r2oQPLKwrrsa2v1iA6eQlIuISFvnpaaWI/X8e
RCXPgdQJo9ZzqF2AAovCLSHHWCZV3G4pS38NaD9aFzFxilIW5LoKFyhq8dD/ul6W5mRfyFwkBHt8
rfv19G/Jits3dHrdRvtaXMFmxZ1R2WJf+2l910Q4V9Bh92XUIAmCMZwEg+/ICFQsXAIQfJTkve1Q
hrrFhqL3DoDmOY9JaeR00a5x7eTJtFltCFsJkNw2iflIqLhl3dQDz/H2zecGlSLpM5boaaFvRoFa
KP8v13gqLpDclXrCopJ+7pL019B4bAczItxm+ixu/ljQyQpTY5IYle8C+bEOevyMzkS7Ui5duTNX
Z1H2xQhHtaekYJVCM5wvvJYdYpBUmH38vIs2Frl4wxqUTy0lOKGB/anPZ9ThexqxjO6INUpEhq/k
gDTp9L/5tvUhjciEDjFbsrtQ2WlOpJKvJVXwDXJ0Y64mVJG6R1Za8C1j2q3N/I4ZXF/lm3hEeOlF
pI5RJwbHUUjB4FvKJx5g3Opb5iFsrVPc20vHILgIZ+zvpBhcwm7tcNHgEl5sH26PX056oGeYeJxO
DLjMr6KjAZd1kxhRdx7gGZ7jmevoAxEWyxj3IozUBtoAKWQU2Ceqo8l0/U9UQX5Zp7Ni1/t7ZROr
jTh+o4KX+WvkjZs9P5zws/eV8npCK/2whPURW3PJX1DRlZxhqW6kIU22GU5u8u+jlUVYzxHBn4kc
oE+pJ6PgHkHB72HlFElztjPODS7XYeB3GiHdsVG1r7kpvcG/D4AG6hPA4I1MkkyxZK9kmaGbANVo
23IFDIMuDJqbQlEhCz0r7ZngL8v6DkM/q4WUI6ACQEOwD44wfhFs+Qa58XR45ZHGUn432OxJmxho
bXP33NydHw24EA/dkQReFoa/6OtwtNtv7ok3tdKYMerTfrh5wkBl1YDx5juULCbcDd3jcRXXVszL
ph3DcBJqZoOanvgfqVdA3tqWxfO1kkfyr/po0WcDdyZCda5Ur3j7l1a1ZUJtoVVNHsRFFsCuPeyK
A6JGgpKZmWKPy4PIo5oUe3939TCCMaFSQZCIBlx/VVdoKTs9peFTtUHi2hEGHGyzi4NfolHTOiz/
Fw4CaW/ICONOjvDEF1THdKQ9FyMBgEgw8XEPXxvI+jZooU/SRgf1PIxGJN96iCXQ8AwIsPs6C9Q7
NnE/jhTDQFjRB8Dulm4pB53V/yREv3/gEXsap36P7dP/gTGTwE8Y41pBVOYgPu12QFY2tSity0Ed
BnGm+o9GXEMK3B+lI+w9yChNzFTowXZnodydBkRZZMzRzo04rl1VAj72G0eOhTD3lFbIwV2pF2pW
h7TqZa0ESSCpVh1Qv9oqIEC5GSCPX34Klda1sHm/xGCU+OWvuE4NJPvNnq/6ZVsVgO2YpwM/YfV/
x7u5efJsrPWSMVVNdgMBCwq/Ekpn93gR+mPBQwZyA4fVGuD/oUn/dBLevWiIgFeNqz0Wtm6F9gQb
jRXobq8tZQPIXUqB53aqtZUE7q7QXN2qUZsmPqOJRYMxkiVthQb+MoogP3/6q8KopLtwPzo8F/IF
2tkUb4w7nC1YNIvpG2tIVHHjdE/Dsb+cd0YrCSVq5LyqU3PHksTQYcBuvDC4oeDrXwV4kB8P1uHk
9Ggg/x4hrdQzY+v8KuMGPIIXtlSaO6sPd21h7REPQVVx7e7o7JwKBc7VV8cppNvKVH0lYDVdR8bh
Rf4Mc86FCFjOy0ahs1bqQByE6r8E6FgAL3+TyHWw0bimSiI494A3ZquZyR0Pg17EnIBsZvavWxG/
ozC85qH4GbxCotMPKYSplP/Zd2mZO8ovcRe32wTBdguXHh6orip4AuYFkqYR2u1lNTgpaVEU0VVd
58jXIxmWpl8RXKbuahV5SDKTgfaRT4YaoB/B8BYKpTwxCurZTI/VHNEr1+fQAqNBaXyKXPtQQDlQ
EAgBVrdsoFOk/UiYBBnVQ5MY9/ZBMqMkkBiF9cNnmTaJxnzuvQBvdlOKH+1wnsSQ5xoU5xXP9Sp6
3UNDCVGQBJFHWKQjTsKVi1pAub9fYgeE+QIRuMHI36c2SZCXZDdojPcVG3nSantPxfeIqxtUuQVS
B9ze5+p0FYf7khcsvWHiF04ZvrIbywcaRiHwZLVW++jsrJnnaFSe1emuHIhVCT6zVPcB9x0yZHSu
bSQu76jB22PzlSNppQpvrTauHSCRkcKxuXZYmykM3Ffqx5d/IEUraBkdOJz8x1NBqllJq2jbVxWb
h4jtwUPpR02QdI+tE1qL7VBXFLdohLU/8Wzo1vgis86qhIT6GtDcplFpi/oTNjocCZdb+y45sGo9
cDgZM36EOucKJLTzkja5lpNxH8hZz7Txxr3pNUWIV2x9jUtdaMiWfuryieI7JjG5hGMAb7q+6TiA
pjSnvmGhlwtvA8UMh+u7wVRtgwfWTSWdUKZ3gkLDB/P1OTMOL5a6HXKMDTHXM+8Nad2S9oGouXxk
p7ETUMqptEg/rlKCxqW7orhr8T52t6CTs8i83AmcOpov2Le865qE/fZCB873V0OLq5yFvcpJiZht
XmkLniIWqf0x5rScudAAW/3N46tDf7VsKrinUovEjL/hbEW8dBEe02zM88Lo4vLz4aahRsfVOmJT
t5otl0Lh2T8O5RbAuYUfAjfgzxeNfwuWozUGuoMgfcvGqE/fqqjCz8ZpbhLhind8qDHy6Htk8GwB
6SyWPbP86jxxLiIjobFAwP6d5+pjxOa0N6CkbYAbB1VkTAQ3k6TJ8PY6r76oJirHoedu6MKa/iSv
xRF4OOq8VsgfgIm5MHG9P9cb9wMtHa9NebSB6G/f2+y0DL75B3pA030zLQ8cyJEMQIus2j+Zdtv9
4pagOxkgCWOM2GMcWrxhd9zYw2CsU9kYo0Ed+iIvGEPxMYFdUOBXSKQR+9zHKjJLkGpEH5hRgMv/
VXtVfzks3Cgc2dcwQ8G2EyYBaG6E7EqqcF5Vn9A9FyIr9B6eGnzvGdq/iktyow/785BysgK8WAG6
6NyHZXghFTPyErEJ4rMaP8wsfis/Jq1aXDdJ1HaJokv2SllZ6G6gCSTkQhTbfVvTtWJ50IfLU4hp
Dg+NaZxuKe5zVgC3Mkv/We8SRbBNRny8xC55QipNd+ln1LOiD11JQrGpxOA2qQJTCTgLAeLRX/Mk
7+FQCtZSdQbtO/JTnphHbd5oacVsU3bb1Mcom8OhCm2WGaI6diJnf6T13cAJDjEgCbxwDynkLsl6
bxCrCDzYSnZ3A05Jw8QijvCLYPM/rTA8b7dvBzD/XmnCML8vmq99v1nx1KV0VCP8qtJFnxf9Fc+C
W11OoMdudHF6jXJY7VQBw+lPMBcAvy4moPNSDjt5yT9XEXu4DWW/argo/tZ9J7ZetacnZh3lizGA
n5HQfSAufmDDaCCMOw4X4Jt5wEBakFDdwX86znSCVfrNYEEruUXz76GdkoyEik3K9RBzB1zVVZDZ
WzpgAuAvwwxhHXTd9Yu8A2e5YBSGSl2LJCiU8nlvntaR7xJngAF2orSsdp4pkm5VDN5cKLgiGaMk
NaY/HGzBcKKS8UQKx9IRkT1+NJH0EXtHdYCcr1DW1AOpHPaOxqDmS5Qal/YUJ3bpMGUZ/h7pZyRb
qNoEK8jSiAp0RujHe20w32DUgEz0xAUmzr2xf0U/w1iP9imSJSzJ8QBL6OfXbkQIk4bRBsj9801q
lsv2TSFDalAaZ5OzuEpwYL7Nxiti3lsAbPu+54LKrLDFY8ZShATa3XkxluxGEav/B7b6KbagSo4m
kuOp1BsRLKBquvNq/rCJuJw/7LFbJjENyhcDGg/3A42YaG4X1wm3Rahs8tK7f5YdLEqQ47FdP6kS
udX6atvHfGif5i+JP2iy4tNR1yX+YX4MeWfYSWAr20igkqcEaepv6WAd+Q5XmdhphoKtSURMqeAx
P9w20cxjlMxQjZMsHoWDN0MkiFRKqPTCDP4voTNPfk/OL9b5uD07LccZPb6s33zxljjYErhzTq7I
QF01DQnMkeFj1xNXBk/2OxraMou3FTqhXBhwrl5b0RVy2H5+LUpg20F79nRhB9H3ra7uFvJoLrA/
2O0pcx11n6lX/OOyIDm3UAa0zIu/B9199LrUGHXgyCgjJny9OR905aMRAYd+7Sp89pKH6ni0s+5V
tD938jZ0lRfA8P4bF7HXm0YvwlJGaykQudKDLmVY4M/NJY8Acjph0fYvC4Y1b3fOwWpE+R1tA9gz
r3tyCOukvb4d1SUaLWcZ7bYvVxbvQg4MgEYGF0+9JQOmIfW0cgers6XXqiTWnCG+uL/jdah7duAb
rUTEUkYs0xd1JQJ2uiXMoJIMqvW8eX/WL+sHNHdf73YztDr3cBfHcgE0I+lqhG6+AjTB/3xYz6Y9
KNUt1JhGuMF5T3mlNDhUPRNezeAZ1U4ATACifrRaV0li7jVWMFiFm4gapIYaUfocLPyXxDSZd5qa
zHSHd+GUpjhdnQgSHahqXwQTmHlxLmMFytugBcZ4nFONoxCcWw0hii7hbQQwWoD/lqb9dyAgvjGj
ygIWLI48KM0hkoa39VsvevRutaoVs+p8S9Wr8Ar2bmVFKtGP61Ck9qkw8nEX3CH8CP3BuM2xvt/3
bYfTpRDXFKBuvd+5Kwm3efqY/bzYXrNshDSdJtJu1w3Nuor7APPLpeGB7rZYYJcsmDnfB/V/38zl
+kB+QuZot1LkraK0UnjZf8vYJqXCb9hWoRBPSFVoMPXTn/9ayp/+WPaJ09BdN8pbTQdqtTv1fxzK
itW6p1P5fSkZ8r7C50kJJHLyKlrL82Q1digKzpMxnR1BmXbGbu0e5pxgW6rDIkd5huKFQuEJCCqp
3MdkU2zf2GmqgT+Z53UYxB+xU0UB7aRLMsVHV+Uvrg8CkBhtaNUnnBuyGtn2OsliDvt3J4Iqlewz
Bn2POzTeBZjqCd0v/flLJU9RqyUgHc2XG7ENDOxG41Ee50TeyCY//srZxqUVZ8ywThzO+WAF1nx3
WPuHfdlik9eJd5VqxbQM5Gu6WUe2VAI8mo147hejei/o3c13m9qWCNa7lBEoIYlKpEqrMByUpdZQ
bKXrnmsFRuoXrAx2k+jqxxaOX/ekoFUZ3U+dPGdx48QOfxrNjO+A5Vn/xFvlTtcL7gAmF727g0t4
Zfyf6ozILKHzgrQc37XzVbIwV3RvCMSazPK2QcpKCbunAL3nb5bdmGuGrnDPkcqaPPfqKDHezOnP
GE3uGBDQQK7dZBtos04mN+nOEzEnocJ0/xX8YYlipXQ6Gzuhi3aPYwRgopPZjEmW2NXd7zhbjfo2
o2SDHiji1N9APEZDpnh51dmdCaY/gfRec5AK8oFRk0BL98+2MKztWVA4AKLRyujspl1iJnEP6GQb
fSggCG0RkTGc7NASFg7i1MGenDLQnI3zCo8nIg75ilGE1UAqsc9JxPvj2ni7w2Phtxko+/tb8QK8
1D3RPggdDaeiWOum1hw46z+bG019vo9uA/Cv3hheGYSmUzLAjxfILt8+WFTo6yOswdQPCBRFTRe4
6UqpvvzP+jNJO0NoOQO11ekquxlCP2uBs0QiNZbXPZG4vONKl7jdWK1PLbwAbyJCBZq6HAlwxDTL
nBibe7140h5hiZyBTZXaeZdsd+2uuab6Bge4dUscpao8iJ5+Wg57ihvkqTEYwHHyEqyyesFM0FsX
MGF9tX3EvUn5LaTB1B/ppEjn8yalUtZZrMbmXrKJGyj8fj0N5dYJSsx6rkq8oFPoJCc6Nqqk4HL+
2+iKA702amZJ5sPRgLFGcc+lhMDdF6qCLTk78daTtFFwxZTFBdsPl0Pnhy1IvhtZ5Tc/zTmZiUJI
1lgxxT6ZOYhiFNW9/TzQZXAszEmq0BNq9qWoCBuYawjwhJqP0nWX6r1PGeaqfGeo3+TaxCULYDW+
2dK/lmC5OT3dOV/L7b4t954vPLyX83icE4aR6Qj5JDuCsc2AYz2F0JE6LtUM4eHCYTPreTsErmWb
lkTd7EaJn4gqneJGO9hbeZOZ7BW/5EYxlWuqeZSMtRf5KwxajfmE6KcPcj4rldz0E4gy5BXHC8kV
iMtMcUCcnsiFLQWIA4xKRDyMfizv/bh7YreEjC1layPbmyA1amfvPdN4+tJJRj5N1/5+2LDdHSNV
nzEGRAm/g06QVja3lnthG+7OuqTV/XhxNdMOMIs4Kt/RBvA+P3k0KanS1Upb4NUvjQwXdR/DSodm
fSdyWsE6sNcZuadEplArQEap9I0w8Z5jHobl2+ujDuFeOUWFSiuzUgDxQ8k7RgVjW8KABjen108F
Gj+FcL8GJO81gw+q1blOp5vGgjRVJ8oF8XM1jZ9kEjr4FTZc066R1Tqp153IXbX5q5/rjwNY8x1N
ENeV8BqizMHCJKSjDzHss91iD7GMTbgJnWQlSzIz7kLDFuPBVOuS/EM6McLIKgbg1zN6Uzd3E6QM
5pfwwSwD4z0oF/1Yycckex0ljBkkw/AtZcif0IpuUunh/wzhUBO6axrfYNX2SJiqf1aA3aWYSh0k
Yvo7dEJiAGutzjtSEfzqDoCn38G+WWhFtD4vJB7L1CG4QD7o4fSRJPrysWJzTYmMMLIckINPiZME
7qnr1QGZMzovZDEe2l7QdSwBA8E9zaJJp85xs4dTIHNwEeqAN/yOs4JB9x2evYkCe874iwxX8sJZ
DUAfwPBd1wPi1+BZkHDo3x4ZZ8JXVSE/srEf482vWPerABbHz7ByLcmElLNUmgrC3bWI7obvxkHm
VntebtKbtP34N4wYySROfMS9T4yUmK767UUPuJQb6CNkQDSgBSveUP3+hg9/UdH0PolyKvZ4jCym
GpuLvLMerpq+sfvKkyakooTAS179SvY/lkeYANmV7SeKVL7DqUWNZXr6QBqN7xGART8BvHwD/9YK
hDdxS/rVCSZdXSoP5uKalUH3TrfJyXS40tI0pSTrByqVukN3IMID5+xm+U9x9q0NFv5QjKuouZvl
CaGvlNs7mDqx6U0J9lAxPpRAfiI0dmFqtPjAGRH4vhP/LmRXruk0vS9d5EpjMg4fVa5Dq7o7hlvQ
TcGfYO6YWbG5wKcGXUe0IiE82YT/BFAwYSBtOFrlxsEaTgYMt+QydpvlZwZPWsSBPHcrB95pG6IY
wbYgF3bgZghyzM0zAbz91XjxYVC7cPck/y7al7PiqlLzXEBHdQ5qCoLPIzH73vrBj8RwEO232z6J
I8QbzDVqZlIk17x+Q2IEgf8pRVpMCw9EaWt0/wJVEm62HmH2x8xEMzJF7n0Qm6ZNuMg2Nh7jt/pb
ee5hGrl+n3vdkvQ25I2wG1BBj3sZFmKjg8vlB+Y2gB5nU/uZnjC+PB3FmFgaQUwysfTCHBcxhL1u
Qf0KJzolCEp3ABbgt2pVPHSjqhp/JmB5Kf0iIxqm8ByVqYFUMSCYP3icFIzsH6PEA6eq28cv1h2M
xN/ERyf1bLlEzkCvKTLJSHq1iA2X9QwB6taFyxIp1fZk8MXz2aiFxZOtkRGtn1HkO3cRv53rXKXH
cMqwtYFXziPF7gYWubr0DzPjO6HkhLCrNQd+bULdLJViRy2OD5FZwoeWFUdX/A/nxB1R857EomJ/
pmlQhugHHEN8hMUvmJ2rrQopDR6XN5Nmrv+lEu5qK5P80erpm5IwoEo0gwluARemO5ofu+npY+xy
51CMCium2UyJR3B6erwWJ9pBJOFjDYNfugHmXETFpev4P0Ed8j8B+DB9IVTUUfcGtKuWl3/1Kft4
8nTJSDlZ7+EbX5PzTYTLu0CUE6t5ofn2U9jjMBnSY6JFebua02gu0RHHdX+k1hublGEFj0IePgVn
6cD0TQinKS1rM076gu9NK+9ZquWqQnecPRkq/AzDaL+IikvI46Xi8xcYLTTd/EqdIUaX1RLoYS+c
RyrWviFY6ZRuYkCrVlbThbfL7+dwcnhSz0NtyQ5t2FXwunTXrXPonRHgXm39UFVn/8LRDiT6Vkqn
9WZb68eM/1MYzRrOK2CnNsuVlmdWiFmk7cV++p3KuMRKqIgnZW2q3Lmc+7J9ayoOgpcX3EVfT/7B
bynjdCCf4FimmELBJAs0l0UmJhNomJbZMA9H6sx9RSTwBogyyczyI3giZ+1EwXTAzw4ntMNH83BN
SN1l82R6IYUIhAdwPkhwAxwZYjrwptBodpnBvdEiy9BkPuEpk7xhFlDcjAP86DMLhx5iznHBYCcd
NbTTbqmZLyGNfMkqL8H7G/miJqJfPBCGvzH0Oz6frSIMDrAGLbUENn8JVDo9wQ3sw7Sc/+7YkmQp
z/i4OFrKyMbpmobmQQHpFVcD4O6Gy7jTPujsh/oVTf3LZPHa+R33W+7CtUnHxa7lvPZ7xMt6ILFp
QyfBBHVDVsnu2BMArobTzPKA/TaTtHI6S/hHOvN28fVnrMLya0UoOPQictkewyCK4fcisJpzoU3k
b02PNJLlIvMqoJbPAZALxHtWPF0bSE7HK1BkPtw389Ll5AUdTEmE3deCm3uq+srn4vK9HeOKjH1a
VtiiNgoNwonj42EEVpxBEKjymZSI75w7FL0aThv52+59Et6MQyO26qvsNtZg+P0B/oA7iaHQFXvJ
IHqozTc2xGPd3DxbW1sQhIqAa0LMZJPIiczahK/TLkIqjvSHA2aXytbp/6gGJRW8iHd4+psrvpQq
jhhca8oCNm/MKtxohoXaqwscMlbCAaDtEsOmxLOoT5XTAdki/DZ6IKx0dsZn436eljplwUg6U30g
PjG+dSP1dzSxOKWav5Q4NMvdQcB2TAY6Oz8QEBuz++mgJZqlhqq7B63TrrM88iqo6aA0hniFcRrT
/hT/k4Vs++7fBm2gA1jQ5e6oeKK6xDxyCVUV+BblL2kiZjoNidalP+JKignI7hlU5Q9cBJv+NkMq
fx0N82yXTiEaZ5nnYeuPcMVPCHAMdSJIdj4C59xBqXiY1Cvp7flIAMlDP5MV2tfsDkDnGrIYX5Dy
MEr9O5AkZAeiYWnW38dEczWn4L46DZgZ/7C4aTUHY1AC8luKt4xiRL3Vtm9y33ZMqanBFwt0VkDb
lh8Tw4AYDsZZDw/yoTX/agvIyXM1sE0xrVJkUJWGy4h5qL6mzkyu7XHk3feu153I7gfbc2UpgvjX
WKDY6zQV59iU9w118fYTOxsfIKrGJJMO3DXGxbxqinI/ZclGbZ7WbQKRMDcQMLvPdPRurTLpyOqd
QVTViJ4VRT+ETdv2CYvhaWO/hpFKw7cTPnqLhHHDRj2bV6F7+dTNv8w6YBrzhhWVRFIJD3h/iAyR
ewH69Fp3pNtMWcF7j/qg9vR1Ya4rWX1ctB9BeKHkKSXSg3fowcOGdNmi+ZfgehSp+B1kVMtW1uNr
ogZbaYz87SArOvq4xaQX0gIaB89wmAjw/im5gtBFpR+Sn6EM6GS4lmJzVw0e6i2cnxW7sHwJHKG5
M9sQoeVB2qvWN+9uNFDNr+4pHmFCb4/4OUr8kStUDIihhhdIDlenDQalsH6hTLLCVi9TP4qWSLPb
Y4uu2MsOU9nhqxzvgQcIV8bVT1ic+6aP7Cq89cTJeGaGSrzJM6bQoUBwWsPqbXVxVHfC/RTWbB3/
5bv/DVa2h9RarwowCL/+tGzm8BT9fYEtX6WSNpX/zlOmpTNZVtk/znPeUmJxg5UeQXebIKt0l8kR
yTes1w4VnArtAj3hwoTj99uKuH0v12ORUdh86+/u8e0HNVokALHEbSXa5qw56m3tKnbGVaKxzjSz
pLXPaHpYbbBRfCY9IccqvqTuPDTw2hPyyhxfAWaxcTWxqLdl/CtoHi5UEWtBH7/JdiWs+u5+5iWL
oEdCue1DfhvuX/4surelr0+EIxjYrpv6GG0w9ymy6Rm7CNnrNgWKL3L6sYqH/RDXGNBeVQCD3e4v
PiLUblu2bMuQlCISvINvaj/+PObPnnRu5DQXeM4JePA+6FLNXV/mWDj2B3Thxrk3AJvynbXaeJBD
GCWv+H9WZnelUWEWS8la38DNgT5KRhBv45s3dwP0XkofegAOfm4E/gDxWWL/NSDyl0Y+UySvkH/E
IsWTas2+D5M1RAMWm/YXnm7cqDoW2E18a1MO9oZ+ze9WtiARZfqLD+3wKOFdX6bMtlKjrw2P3zln
Ktvb345CKmEKE1Oc9isNJ2z7Wk2luETF2T3pfP4W/YwRXOw+7VyxFoIt5DWjrhy3caI3xHWQAGCt
khxwF8iTNjCX+ACAI+xW4dro8VY/hu7J4fJcgTth6I0ZXqduMedxIHr8ZuErOwbENCcF5I4URNXh
rMkwMqye+COTC4bCJ6PLLCCiOo69QV0IgKf0JAiEShcp2PsEli/nWv6lxRIGsLYMolGayuBfuU5V
INNTneyXbBdqUNoAkJkSYYoTrlRS9PcuLCR92WSCq6jeSfrKvhYoSd+xCGXQr8komf4k0MchRBhv
CJEDXXlkgWjE4xJW/utJHbgNK4qhSiddue3z/fkWJqlhkuxPAnLVRMajQjifL/lUb9x5qENjLunr
UCMdinyDLNkK9j/jg+hqNTWo3vJs4hPnv3YEbxoIthgg37G/XgAgY8LAIZuXXIDg/3KZNkg84vbJ
FvrZtqnYZYRChxFVR6pVQuGCBK0kcGcPYrcuuqadCO5NP1H5qD40LNh0H0c82tOg+4I/eHZNppOx
OeDIB3qTF9kkCO4NFGMLswU4/Mr8NyYbdCedueMoqTeZolSMM2anlvfWxsfY7eJM+0leZXY7+UAM
pFvwLnGP32f6XM1zK4HuwkySZMDUMZVR7gZu0irYrTg4jFmacWV6dF1uc43IzhmvS85Pie7tDyRj
6xkoo4tZ4i2Cs4Ec3n55EwSTyBHeRs9p3cJxUEF+nqHWBtky22mMfY/qGn7CrRMnyOrsJsqFTciw
DDo3ntaXoh08z/wXvTF6A+u4MXSEbFKybO3kSXZ1FUhz1rPBGnLMHvaYPtVzfOH7DuThfQv99wMT
jci0S1MKT74Q7bw28Hx8Kn2sbIVn5KEb1oSZaaZWfPQmbhpJgLyfwfg0V+iJtXXsj+yjkLRLbkJm
AWeKOmmwLecLy6PbfrkL1fZf5ZQRCrheUGjy0Yr+OXzxr51LDPa7CatVJm8P9L1fXznYkLfCU5yn
CdCkU7Rixl+mgO5nF4hWeI/8/d93R5UCDLIKCcQoCzIrLDrg7MDAyRvpzX6BvpMKXG7oUA1tzfKN
tCqEKdphAe5QrxYCyFTox6HKWea6Af1dFS/ZSTBC3d7+3Gpw8Wr+7DIgnl8qSmtxtWmszBE9lxw3
G3xbVMn5KMQXwKKCQMKpv9QG+U1J9DKGJSkc+gieJVy7JahMhrvnLcvVEgExg6SXEbZifJnIe3SV
k89Zux1sAOBbGDfjU2pQzOYcWi15MadjlLFkupza+HY2xJmYgI4f8aUhTl9MkIy1Z30bVQg0XhAU
ptMpVW7QXLQCEIBEC0AnyykCwC1QHw6WM0010Q/aXpMSf2vRT7g0xiwHYqndtVL5ErNckJqU0jZW
GiBsrJ0d9XW5VK8jNSav2J1daDehvgdXH94u/caElf+PA9rXRGlm2wQB3wrNn7Pv7k5UdswikpVb
zLPA/Tpn7cvEfLvlsSyLUH+To51URzkDrlb1nDCbQ9/J55CKqERUeCRGqn9y4od6bHq6h8YPYKgf
EzA0u3+SwNlH1COEmQPZBFGL7dT4Ehwrms3RVvgHfWTyx0Twd4QhMdZO5cymy07nY0Ncg1nziQHS
mVt3o6R18aW5DmQ/1hBZWiVDqFuPs/FrHim+TI23awzV992lKqDA8EcFkVX8SXPgOM54u2XwHwIa
Pp/qGF0oWUnacVCPFf9BweXbWfeYjNBp5JPZnXI16WinSUWgA+mNQsr3spSiaDhRKBfKYiCb5oHC
vD7CC4sSHMdEQxkgEtqICgbNkyGc9Vu8Dza6ZtQs7w/Wgb+LHvOjoOpco2xmEYAZD2bBrxU1Gmvk
Lo26OZPkYxLDNAEAXPm/7+LvwrOerfXr7eSxRBAEf9rQp1Uk6i8w0WnhZIQYsgP28TgM5EJdLD55
xgwTWigC3+4a2j8dTjD8Wd7vFscq3c4X3/O4zQCT2hvnD1Z0GI8ZHBfAGriOuTBQpevZw+/7CuCS
aCY8T1+qPVtRhHz7/HPHxIHzub46Tm9bMzUVGj8C2k5LdMqrUVrKizScfMB5KLePPHoxz0r4iu0F
g8T3rmYcBd8yLTxnwRX6Of9EPktkGCorRykhmoS3V2zjtX6bwTtEfk9qRE0SPslNzEUjvepiZH4i
7jEcKSS4zCQFFY1xDO5/lmHbXF5rQrtE4CBtJ2EU82TnYUWRrYm1Fyo1Ht/1nyLIsvWYpnQg5WZi
G1T883tU45LvO7yUNEOX5b+s38trID9kgDgHq8gP27wTXC+7Igy3KVZxiDT/2m28+gLQRIXw6Q+X
rzJptaW6JwTBvI+t6GlAOGJfwGk4/Hpj7ycwE4B3OB9KL/y6EYT29noVK7jT6NdcMMUBClrhiWuU
9grIpre60hYS5B1AZZ/snBPMRqKxdqS2FmmGil02v82zyH4Ha2zuoGGPaIIkISJ+HOquOvdXklbm
b/SS1yznR/ImbZx9b+kpruvB8k6q6sZ2bZELvQ2bOosmcaxDdTZyb50IcfURz3v7ZyIQOU0IfniC
UXd9Abw5gDqHe1rD7n8/iLt32g2sV42n187Im/4OakgEMVNSNCnQnUkNwqsCiohDw+qSa4YbwTFP
ZKJla/ncHM55vheHQsVhG1Ll6AEqPZKq2bU8BQiJHAcwMoHLDs5qKcdcFl1H/plmoO4c1JmE+l2d
DWDGIGHosZ2t/4/+yUIpZZm8fHqfmdpNr1HJVooCbahczUtZgng62JTLQBCqZOKF/Z5H+aQpF/Z7
Li2fLYg8849v00tQxduhMxsfLOXMtnFlaVpyfAU2cg/gRyM9yfgk3PbP/CUK8xQgqVSWrn1NLf6m
yBW64A8OpKZOb5FoNhy/SBi7k41Uj/Mld5PT+xlBxBlL9eWm7YG0ek9xDYnXjQBmFj/dEPzOf+7K
kEPIxxbzbAG0qWeIkAQi1HftR1NNxspve/UEO2lXXZlTzlPgfwnnUocoHgIfINU/4NPnDSXB3KRO
5uxbpi83z4kjhcPyLYlf2jG1MuNYNmnolKaaxS7kBho7rO7TfEM840gyeFzvC6LW9Lpy4fXOjfaQ
LsulW5x3y1zNumtLyRIwsJqUPp/jSPmRa2jqVQTaVz1tvdjGVfN75MkRCvR6gaFcYKqFIiqVXXEe
sCkkHvAz1RHTss7uz+4fVzt662PtY9cdCOXhMDxXUFKRKSFc9IH93off8B/FFvQ3c/5EAVxvFHYJ
6TN7KipSqaJtz+nqH6L33Unx3v+UvKr0z58z8jbPbOlQt3Xxzby55Q6so89hXmCkHeRBRdaNIi/t
AULW4FcXVm8IBOR1SpRLjjCvHBRfp6DbxJO912kiqiaFXbV+r4i579xP3RgC0iBoFclC0xpNpb4Y
8aRhQlLgl1oXD2QBb5gE/svKn/lqqNUPr3v9oLwLL9Dew3x1ZxnYQag5pURWVwGOmOdPVU6QW3Bz
YtE+xin19aKqVBGc1j1rwgVJ9z3Dcu2prUkIsB3tGg0KFmTb0NtnBfnlF3vyUDYq8lIju/8MuYko
3JYaEcWXLungyoL3QjKVm4S4FE7KlSyrrnLxCFUVhWt5Ya3KYv+o4jqqtpyUwaPd6vejvY7/T5Zu
9/ziasukFRiMDSN7hDVQuyWbHU468i8yrEBogqXjFGbWFlLcUSpJELtjXMxDvKdvQ4fHj+W+KMwt
YAX8NTQQfOa76uE6u/WnUq9vWDFXmkzkeAkDZfxHYxT4esn6IgHkGE+oCBNleya4rrchSjl2MVEp
AOV4QD1R2G/sHZNS0DtuIhDz0QU2/SPX2fY99hUPPUOzVZ/ZQvzJ4tjjo/5rQUTVeJR011CA8Qow
UH+L5g8FovPMKaBx1sNwI6EMwfIATAQydejLicxZpsXrmXRH+lDYozzKRDXebKbNKXB5HJ9z33le
kz32DTB8N5G/BB0TAQ0/1M5ZYY16uM9p0XVfuXfyW/X4MzxJMhvJG7n0+I0J94Kxdg4jsqrnFZqw
5JAHGoQb6KEYl3e34yFevCX6KIzQqc31sboxsqxHQawQd2lTuxlAtY+MfpiY4dVd21uG2u+OM2yb
KKfZVQz5vffmoDf08C3CZdCCcXJUxDMVu3sLblBr1DNvqC6qAe2ksuv3MUnF9jmiRxRnl3V0t+o6
rXCejDW/M1+34+oTnsAneE1w+47umfgkqBh7zKR4j+9BAuV2yBt5EUCBNQjLyymlsbmLecLged/H
xrb6lJJGdW3mWHQZuv5/OHRW9O7Nm7/Dc9weT7I1y01LBNIrYKElSRQVhtpvBC9TB6VyPbH2Ekdr
h1Rb+dBOxNwtCS9D1dbqxzjb4LnOCXpv3AXO+o5QqhJSDdD6X40h6k46tykkdpgU+qw1IyN2OKsY
3AuWNRtJmbZfYkNHjulyTOw9ImBbqhtYPVyif+ws2MmEOFVJn4D7NudAoA7u+zagR8b81sDbp+iL
MBJ6DktBbnYSeNYrVPTj8jrGTzNh+NeUc7ViDukxVekmlBynMQV3tfoSDR7ffM5oDtgnLZj/kpLs
ArXZIpA5O6oQ0bTdCPfc8DzqbysbaTh0IYBFXuqoS9wcnL3VKBwT/qIuEn2AKas0MlJNHYjcSYT3
sRA5PxLq+/ABUJEY7uzHoX1euLrS8h6xlD5aHRVf5OZjCCZpDLS1tWkms8S7tRg9rZ4vQeo/UF1R
Uyvq42scuassu6ibj8bpm6S4mrbNg0mEDagmTlCxwKfFaYSgGeZA7OepmGvKGyEHkp71GqksCFhV
ofHIMMrUzI0g/H+5b/z40Avt8XXZmDM/MNfJBL+u5BtR8WEDQlx5g/EjLEIRQOIHmpXl+9JHsiMj
0HwUFAQ14mFDmic8fBkJHlv9GW3Q99LK8I478ot5diVdg6Ce1VkWklsRhTc1Hg5wEDI4urhtdy3r
ESBXaeYn9DrInMur9uvXBpam9JoYpA/EXdCe0xo5tX1tj49UW/oYJmmIq2j9szDhxGGtIVPIRo/f
bDLg5SDq5L7iAPATMHGa3/OlvDhzmRzu+JePVS4HrjuTY11q2HiALrJDISs5mBB/owItg/SKh9Un
u4BeWicoVhBQ7+pfKZdhjyEdFeQ5XFVewNPcK89RNOnRUwyKixC5Inw4lod7hSAOyOEOq0Pp03vW
VPuk6HLt1bbB75aNvOJogysjDWI5DgWVBP5w4wqdXduxZ2Z3e6X4TyplUan7Ya/lJu/x18E3ZwJS
VyRr3bvEvJn4sMKHqvVMYrvTskQVLxh7Xe2hxOdQq2WwzY9Xi8+LVXMQuvwxrMe+LdbDMu/8BB9Z
giL1PyMJpAcyuyNqA7BaWxAzX9J+x6L2jIbcIkcG9/HdvbGdBVTPba5vAOD6wJw21nxANM6ekpHy
/2Kf3eZRBoGdW10RWlaBehTTr1CV8sikch2u8EhU1yjZAC26wDZ3AamkhBx/HVmxkC5St9WD2VKF
QcwyfR1581LnkTxaXvhZ3fYd3f7jNWywCo9NLy/r2NZxdo/HPd9RJytAQpH38Eo8MUmbthTcGWRS
ncatuSQGVvkngqOJ3TU5uoWRT8/gI6muaYaNtsuk17tmev2LV15kAz0E3/2+GaskrVyj/TsW++P9
LxCyt3Ou60XCHmaG9YoIYb3hGLXXJlo9rGYKbjMzukg60bLb08e9Rv8Xaw/MfGEqNp+IbHqnMIJi
B7u0Gx9gb2Ns+pqwqs11O0JTzw7wHZbhxlUSmsTwmQelOFCQ3ygpbpPHsaymbcDvcsmpd/6wlJV/
8npiz0hyfoKjAdGre6bXgHwqz4FVcsUKnTVIYNcMQuCAyZlrANdyAZPOLHJnYIWg2J1li4x2pLy0
4RoP7/hcFSjqw6UptINQXbD2rCWjniScSFQUGyxZfidRTvIzB2lO/VZTECrO/3YBa5uRsgrzNNTz
9BkKyYpB4D/V3qOIM10+rM+0fQDyYNp1EWLnejSZAYrvT68UPGFGYo/kFZzZ5wNbFNU9V6OvyWJZ
DXObr2GBcysmlH3/VJKdh2zoxWKf/GjZE+xKO9Hbf/8rBtBhd2wpBYZnvYzJaTP/kF8VYnRcub/M
fNKeGv5j3SRaPritypAwePiT35JWQG5Oy7tRg/oos4/Tk++fBzHKfWorfzd9ZSmbupz+tCB9YxE4
8k7FuXp26n+qFUxL2zS+8embe/kix5k16kYD5r6km9Ah7pSLKO43U2Ph0CVMZ4nYdkwRq/n9jO9z
/YkEeXIu6owC40nNYOYbySs7LlbyLFlKenb8xUimuPTCKI9VsJ9e8TUnZicV4vjbi/+fqwiNMl9J
Bv7fYWBRSquE+WaaTHzi3ipngy7OqKqpKgjZS+b7BpxwWVgJqXKZGEFgVrPvqwGSkAvYbgd/S2BP
z4SxQfGlJ2kByalaoiW8wjccvNM17hITWjt9KLW9rbfmBr38to4p+xKlM4M/x573YO0l5xF/tYk9
NS0MDEouhtiP/7yNWdHxUJR8Kl0hK0/UwNPSe1bC+Zy3HEajd6QHNgCPmei5OcgiazGJMpQ58WH+
ltpAeVY0/uNoz7mCWY4abTVerZ8z0KmSMI4WHjv05FN/24JkiYnxsr+HYeft0OWAApxEu12TnF7e
5Kl4iXLoetmAeSbbfBpsuMHdMxEr9Q562E4I1rhVsMG+U6HJbNFbGKfChH254vlYiUjAxtT4JnfS
zIEBJMuqIK3F9CNMx8QnpUk7WQZFIod+qDOoeK2t14c0pBDs++Z4cv0QAWLUByLdlskYPmkWusue
4x0dZaIupJBTJM9S2RndpsBlKniidWN6N6LNChH0z1OVTkE/AH9dsiiITc6Ou1QlvecSlU7EvNtK
wCjg6OqfUxCjRB2XINoCzM00ZYPMiL1bq6lTb5CxBQCxAqHS7nIU/E1+vZiBEaKocm7Xes1DGTOx
UxZ8nVmuvvjZOboXrSQFRhFXHH4eVctRP3aEI5QOGXGwjqSy6I70CPu6oIFZbB93B1QxxqVHr/fZ
dek4YNGyBTXc/Vp/XOs1r3RHoBDhsp5SJP8y7Yp0ebToZaun+/bBNVapK1Bq5XiiDlO7VNLD1MO5
fBbgEcAvWMEELM4LoQGL3DKmixLJnW421dz4ZZ0n9Z4Dzlwp6oWVXb+Qgzm8C5cey39ivkYpboUZ
JovD6KTqGb9XM9hN/t7cq5DFE5sQD1h30tDGxa8ekxqvngLt6p9VzgU1vA9SBc09HrAaFRPYRTbE
zSNRuaMVUcVAAMa0actgzsB0hheCWMH4G2RDFmc+4DSe/QM/+ey2UBSjFMybVr6t/telYcEIB3mO
0LlFqDGfPgidcxROgccb8hPrIA7THQwFsBSg82/FoGvV7kuSi0crwi96BoRodq1FTeH7sFN0FGs9
D76+O+3+SkiWXgL6JUBpWTrFPoxlP1EBD0bnFs/h9WIZ/bbIBwn/U5ryYnYUeC16+jtK/NZ/N7q4
XET3pU8q2M4gYz6aiXYJJOPF5sc9Rq5RiMPtNqYQZJfkTDqCc1WCD2paBJXy6B/z66Ptlikki/m1
YGg+pYj/eBR1OKjSYzG0aHb9y0Wf++SC/rPJ0zhpCo0tsImonqW/3xffliUVxxBiRInfWheezC5j
dn4e8HUsaWETzhi1eyoPiTid/NAFGHFupCmyGnK/84gWLbD0EK3R/PxNNsmxNIBxY1dP4k3FoXR1
EaGtubJKvGBsrrZrEAnJCVGbH3JwQFBqgBHzFFbPE0HpI4OF+LzVVqZh2OK6h/VkCQeIt6UKmSqE
6fmNMd3lTyXUyacYIGyrmYkDUY/o2uv7P8KgPMeNzy1MDEfmmJmX3lbWr/g9mBopH2bdF9TYL19R
t8OgclIZaqVHV4yDhCfnwvmkrcgSRuwbTb57CDABiK+sRni21AAc/tJj+lMVLRJ6x5i85NUv4qp4
Q+MpWJPNCXxEjzyD1MlmOUzYrHmkbSb3QbI2mixlsJP+PWR9ijgs8KLlrSVDTfciYLDy2KqP9wXb
xfPu2bZhHBw0hQP0fci6ide8jhP9fHhZ1pyWmatjwTgd1/vNcCAKWY3Jdp31q/kWpXzrT/24mxqZ
opxjkipjesoAo8zvP08jAgkAeimbk6rv/6bpCMslyauC/LQqqsb1YmNOqrmqRoeZTzs6Pm+VUrHm
j3wUBxTYksfWXF9/7Dq9+5Wm5W9DWpF02DE2iJ6J6S+M8xfF8Lk7zPdu2Gp8Jt7/CIhRpDlchf+a
yp+UqRfg7eAZmxRCpbA/0Tfu5aX+TM21Sq/rqNFV4JZT4ziNajchC1fvAidMYFCcrolEN9t7sx3l
V8P1njFn0wVqEOvEv6PtLGFRwmPvz2agVfDBiuVMG6TBVcwRs9G1NZB39Nl0rMs/f3UNpyFGv0ll
sPWTTQMdNG1/nQ1efmxcmvD3R9zqpo8As3O7FaDZGG4/1WBmr+wTZgCrZoUxzR3vYRjU2FJBGNP5
n269ABarOq6nJ/4dVyKiCcTSfzPB5nOAxJBiXjw5MW0poajP+vC5fgLZnZtsI/IpFcGiGw0+oURK
R5mE3L+u2HQ1aPc42GhN6PYRgEY1N/Nz0KlshDNxhmsv+tRJ0aeXCLiwR+RkGH4fC0RD37zkem/s
e/y1WLs3zfWfLCt+FplwjZOeqnqcQXO7RNErnyMG/vBHtPQkCTuc5uWfRxH5phLwyHv5Svx54feV
LdzkImJyumtDVgcAmWYJ616eUsWZtsHASr/62caXXw1C+pmOPJnfLr5zq/aHcmtSjDj92ZjPxsG2
ZGaNGJotW433fQ596Vus+iY/UMdf2IDGBwFtGust5KDfepzkEVzt+m88NE3nfN9CH5bO4KxFFaHh
tuM/dVhZoHgQBz9Iuik1/Zn0zZIP4uV05WsqnMlq6IOAg49RK8RdGeNep56UrkbSjjzk13EJC00P
FisW6kynX2eBhi46b51qEwM2PdhAn3OGKYlaRg4NC+sorwZdlHwrsUlHvWfnrG7UOqxtvctmK6rW
/DWg4rtUgJHWadwrtGWygW5w0+wPvjjsBkjWB7DNay65Yrx1xm9yE/3A176CWBmAtdtLEMuFGlRe
6tDV4cUfOkCc4xGk1v8GQPJNPixvz37NvzN0WRNRTL/xEORmTXZWv4GDyxO7RVX9WRq3j3hkkphx
cM478eMPsKmJOs/FIE1qCYwJ11ssk8+V1LqiqVPyQQOEpQjpUwHIZBWypd0UlwXROvegG3eMZMvg
t2rvJvcEdkS5SPusbDYElOGRQ9DODzYunL1k3iBL8az5Zsz8X3xT+GOVJZM2hmQP7mHuXgRn2TGV
/fjlUO0PuOPPJy5oyEZwgrN3xHAGYRAP9Ec9KerQM1nHbDv96ZMyJE2Jjkj5RSSkVQxrG29Lopya
SC9tSXO9zfCu0Kp8s2VvFAusta4AooIbiDjl9b0nCgyJdq9eKcIBnkn3kiYU2lUlaf5VZDegNlSL
/Yu3F6YS4RAvef5cfeTTksw14FyJ2/zIICfEbFVMv1iEpBJ+sJEIKR0nnGIw1YBra7jQVewFKaMk
ZHMDZ0x49FynncBBwjYdqdRZGZZWBhMJBHprZeFZIlaUdhTl8cZToXN8voSFb9O3SHMBcEppHlzM
O75i1yAhxSbsukroJREhaRfUeLG1EbCNg2Mp+EFpWSD1XD7HmMuFEhvpxP+YIrGBWWlHO6871St8
eMrYFivh9oEu5flr3rBayJ6t+fXxOlVwHJsrxHj119Yll5KqeokV2pu1pcC6BeuZCSv/Xx0eEMRX
qdcgv9d+nVcNGd+IQAI2mS+Utz7bIP2xZEjauPUavGTlMNf5+GODT/SlG/ONYcklpBAWS0RkVCUE
ZuxgQXu9VE3Z/kl+1Q9NB0XsOcajJiq3dgOTOO7G+e1KF2gcWrBQchSsxanB1eLCbnjB77Td8nV3
jogm46JC11iC04SCWvdsQMGO4HspWuRMd4nIREbE/8v6nukG47y2m4LSy6L0GlQk0rHHK37djA9J
+Q8/VO4yzjPLKQVtKmrLwwZF+Y3JxhBzb1g2zvUca+o6dH1kofF4wDtY7QqhUcLG5RU9ZZOyVlYG
+9CvYSOD9gFKOX83655i15/TkxqCQjbQRdKiKTN7u+dBXjKVdSGY7xVQ3aFJIOM3wj6wY6OSiGLH
gpLzL9hMLpGq3de2N0IJSefH8dvEmYcwcdkKhN4UScaPnKpqbSI2fc76E3LfLw4E7rbICrX0EN4R
aLBsEI1oldK+M80YXOWkeauhTlvlCtkXxmIMHsJzMwk0a8SOJEp5+CM7+n2MS/ZJRntdLV1e4OQ3
0N0p+HBv1DJyC4pZYDuBrg+jtYTzxb7TChhbNRfrIgV3ePRxLS2s5Aqf+di/6fxzeC6jVNpYrSP/
62nVtE26YwW4SE+sIRsowQDBaIP0bSG2pvKKLU7KYT03QyNCLqL5UWw0eWHZJ1iQoQjd6sjvi224
GI8MVwgJnU92IMNs2R5UAhW0CpB+QJ5vK5yCbtuvzbxy8sf82iWMbCvtTiGsO3JV5GYzOnGW0XyF
hI3Np51aA2B+OvvUtLOW5ShwcMLx9LwHd/SBd9Kt2MWsL7Vxa7T+pgQxfV2ZXbpnVel2hde7eims
369pWLrS49gIVbUcLpV0XwiSe6REAZTncExFxT3QnljPywuM8XbQyUSvI0zj/OIifPqg3Dssdxmy
NkTRV/CIDOzRHReEQPL2Dm0UZeQRum3BVF1cEjx+Bqpk0vgEbnRzJdq66pR7IXHBx36931AbI0Eh
7owF5LhDl39xbyUylx+yXzTk/kOpDXEPjb5OtAQIhQoNwaU7B+ynXfw+cQ/l1TDDR/h2vz2lN3ZW
pbZcyFKTuULS6ZjUTz4nEDy4Q4UZ4qXQrP2t0nIjW8VXX1zwUzkPeX+ffNzK1aBeWpDgD36Ypk8p
qDnvLxEE5KRMfjku6hm1JPt5M53ARp7Aut/38+lrQ1fOteA4jsuyYnfLDF5CuRvVhUyt9ghuwR/l
uUl9596h9UEfIk8XrXkyahHvzXinxI+U4o/yisIklEDy+Fmz1znAN9lnn+nCVWIvleTdvL6Qpylr
s77z0LAsifiML88aPiVdBvytteT/+X0zL6zBws2fpQnkA3vCahVZ0CUk3tz6xS2ko/7jP9i7MDxQ
6s23LXaqoYupu4/pVjVR/jv2L6LS2csWDu0TZZvUJom7q4ZooOUBVoPB7kJCqDgP8YCveRfU1NOR
vzB3iNzKXCQtQKkrMixJH/z7Lq9dLCQJKpDBnv6JEtWAixPK6Fxzmmt7tr+Jsx2UFiX7oEoskzcu
wPROdFQERcbMXv4ZoY3Ge9MZJVuziOGFfQfeCKEyjA/8B0OhDpYfaqAwImet56mYdEVu6V+FgRcT
66aWf2jf39vY7Tz+Xdt5hzEq5BDvYAWLxjXgNMHC/7bebk4vCbnMciSPm/ormhplOUoFLo2ib4JM
Lzzw9C/3+wql1DMU9aNVjer4Wx7xB3XeAUcgLUAqu6Thb1gdSMLb5deIN6dIbV0xD554hu1jW4d/
0GH71nVVao+IRWr7O/cg/QJFrFHgFFXhIPsi9t5v3xfMfZ+BQSVJeE+obwI1hFSuycyQZk4JmOSJ
stp5zk5qhL2fbwJDxa+ByqSlPcmzI/RiLf3UjDw/ng8GTlYaAtxzyyzHo7Z5rBbhyg14xg7K+ud7
ippBLRMANo800CPs9RaLnICS2Am7AE6Y2nQzAX3nA7OBS4/mi/WUffYzqDXsnqIhMlZ+WQQQUYA3
vFJsOvbAaPtrSHbwsE8rpT844FALgMw13/ZrDWfJgRlEeglFYHZA0QdN44sQaooZeN5FyVmcB1Kp
FHBMwDtNMr/AxSztsgJHni3/zl0aMXCyEHzaN1QGiNZ4oNPvq9jwInzH4BE57Sw4fj2BCdc0RUJk
FAl2Mx/2ZeFTT+E6GOBq4f+EiQHYbFIR072kC9Xfv/T2onm86ARbEuREgWr+XBZj5EryLbbQJMPS
LoQg+rRObfakM4W7uaXJY6G/o/9O+1aEASdCqS070qe0oOS45WtNPShgCmRhPZ9cYIw6XdMoythD
Dugr7mlpLLWy1x4n3tKLpg2c3UENw+iecwyIJv5uO56YFdiw7VVTNRQLHTPFf7VEsFzbcVWAX92h
Oxy2fYmfVGQaEfnqgmB56AQcoQsBG5lI2N56oMAmt3W5j0suL7ursnSKhlqhX65tNAoQ5++LRhNY
PFJaFws0jGLjBItPvcd5Icqy460Zc7GLVJhyeR17HKjYRRGzA5hJoyZ4D48YA+5Sp5cFmZYTjYSP
6HmlvR/4mrO3KaK/Cz99KQpS4DvtSaT1NyItygP8FFRkD7wiZcTGVRft9vRxk1AX6QRxIfF2MdND
pK1qeKxryStY1+363hfEB+aXKUP2X3347qeZSVEsDgaLYqciEk+7GOaXJ3XjxY0XabywkSrYdmPH
/Meh/VYia+B1E6Cg+znS5iOmp5K6UKPNDJCDca6MngE4Flgv3vOZZ1Bug64YLQkNazzOQd8ubbS+
CluIKyr25vacad2W3tW829GP8Fy8SuQ5wqYs65PI8JtimJROSoxO/lE0RQm7UdBLMSVzbo0i4w1m
4HG2ustNumSfE0WGHDJ/sM7mpiAQZOQjIiBpLNXaVDvMoGj9q+QFIAzBq4zN7SmefO8dn5KA7Ql2
fi4gR5leYNQcv/DF96YV6rvn/Zz4PN/Av3Ol8v9AHWWFH7fwZVdY8h1I2fbcfvoEjLiV9kGqO+/H
Z/FPh80gO0zbN+EOlDjWL1If/SJWcKcYUIT/5IPbCUiDVFmRWTY158kHwJLK4pDsNdxA5/JavbNX
zJf1VIbA1oo+qfdg4K3bs5pDASqp+GCO1r3ZFNdio1Lk9Ze3pIKJPyi+l7yup8ZESdXoVwBIexVt
0a3UykeDKHewaGBecWgafIqFr/sTPwYOGGFNuVpEuBDDf2qw1PcoSrWp42ZklN0Q31QY+LEKIgds
rt8ogOJbmTyHhGtbrtfPF7I+L/hUM1adluJOckul2Lcbi8UJ5s9mzY+7Z6Gjmfnvm2H7ThDpLHvZ
7V4xkqsU6+Dxeh1BzoM0c+xvmdHJui/ioXapw0De0wYh+GBQtHThrvlG51tj77jfeZi4TYxDqbst
aRHcOOna3hBR5+bl2rrgLb7vfH6A3EmGr1EpRuOyE/W1JHv7dglLurpz9TwJi9k+iqg9EKiS4Vvt
kXkhNdmynBSzuWhW4gUtxHes/vEFJ9eQMGe1p7bEl5SaEEc00SiKV0sjuS+40wVVvZW39/AX10PZ
uIMbgMDVu2+xReCAJeHZNA1KSye8hTUe9BE3O+1ob4S2MYgIMULqdZZ8VJkTQ2R+54nczbWC/8LK
lBPOYEDkjtLfuDnFfl4zm9zOVXJ503jTMehq7oZ/OXsOx1ShFLhNRHnO/djuMytP5v+99LseSMOC
Qbo5/tidna21bsxmBo/cCieEY8xvZLdeXiyAnx9RT5/5sSleJ9grw8PkQem63g8uTqfn3+FLuOye
fhwr/kzTwT74XvDJap7kKJyTyaCocvBzfctq332vDToPh4RXGhB5/L6Z+LDjm2WWnq4odQwUJRHO
JkQsuF6JuMq6i255qp4F2U1ZIHhC2Vn8o4C9K8Q2awuwtL7ywdgxh89k8QihqeCP7hbfTCjvAS1S
CpXJvPwqPQW5HrGgznqBLpVvEwIeAml6ah1ZLnE9Z72vOTX14nHIcJtGbsxUdLnZMGLg238TqSdx
xFzSxHcOou4Qzv20TKeZprv+fAlQv9/2pI1XTLXsuFx88BEdw6/wF/33RmonJUB4aWxAY2SagMUW
82SwuyJuECcxnEtywkJHL1p40L5Bt5bCpFstlO2qAm4yygd0TzsN86IJtcP1SQ1BBWDjqyMBse+k
lSD6hCGBSzVWXtBXfD1aPKNCCeE/MyE4vODVsk/zx2vS0ggxP7gnixWOqmHDTYvq6fBGQIGOCmY2
XtFRbd+Y+SXWT9sWME+Z5MHiOJGGMMeN59KO9nK+Ircf6V1KT7JptTxiT54V8FkWUDMMGfWYkYIS
kvcVL0nr9A0Uc7h+P7eWSMAhjI1CNJiLUps58BkAtAYc87yx7R0nflqS0POn301KLZMlKjmsImQM
OZUrMSOQJJG+NK54A+W4r0zWdqPhHk+XdZNlyUgKmahXrbX4ERmIxwVqnI5nrv0I9/kKD7ECe/Z3
QiP+194eBQjcjjmDiz/RsuG9S8xKfYhbX/9yTW+dqub4hUgbrIKZh4QfX53nEn4MN3DhIJ/M1e5Q
UiMAIDjxw/iDRAFHtshHFGFYsSSUhu+n4em8dtCE40l/1Q3pbt+BhlgYFnyKLdTw49dYySwdo3BP
eoJsBAUgBVKEnaXzPb5ApTpRF4P/kzCVRHmyl7QENRdj8rksX4FqK4UR6/PpIp1UCQoRUi7hb3by
XcpRi8jgJSgS2XY2+q9cazBbq7uD9HHwbdbmnk+ohjva1TEpRJKSh7OyV2vxCkBl+CSGkBV1ZSlV
pSfE2b0zbtVbblm8F2QwR4SVjfT3ZWIJSOKQ5/ucVvCJKH6RIqowgeIe0vMOIv7jQVlexvpKnqwF
ShH2NTh1fj/U7vzkEIdTe9jQ/KY6+kir8p8o1Qt89NaQepm7csCBg+X3vwVxtEzd9S5zlgQ8qFzt
uZk/7a7xSWlfHVBUnlaCUI6FadYU/bnv/DhJCyPQqeh6uJ8NPkdHzS2NteQKPDXPDB5C3cVVn6ET
96+uM1BKkK44bDyxXL0vydtgZ9+OCQpkqSNC3E5/CuLEz5lQd6JAp4lxriU2oFPzw0gLoSLSAKKa
OOOH/7+aM6jiWuWfBq3JHfA4sVzqxGa/rZ0hUwnqynG9yC4bNx3Oo2h8Kh9UScRpKtKofKexonIA
ejPixZyRe/1DpcbPCtWyn6C8oeTLiNEEDS0M318BAFQx6onPlkTrHuyXoXvXDGrgUKmrzhmgHGTK
5nN2tRnLb6y469eZVY4C7BGxUompBp2lAKwgpPwOy/BFpp0NAbXBH5qPjxJ569aNbv0u7W+CpEO1
6gpCzXDD9RmdqC+05WJ/VUB2kvBmmR3aYyjVVBDkBsrk5RmLWAeSUpsyce75PWCE1Z9G6G9VTMbC
aj0gtxuexBznxM+tRXmM41wvhn5L2yz/Esy3WJ0u9MYcwW4vRBAjej7yS61rX/vVmEmiOBRLpEAV
/DVmBh4GhBqcG0arat1OQIbKUHNKNpN+1KG9Q8Jy3t9QAfT6HimuFmRA8FnCiRh7GYLQG8i4/FL8
iR2uK9VquCWXqsCLstILSLv8cQKSNxCYW7sQgAu3jq+9oOU1Trc4XXSqghHDypvmWr5QVdr4DoDT
bkXtTsXiHvoIM8Wi9ZmjBtWgZXOttutBEOFAXM0itaYllKGeIDkfuD3Nrgex5N15vTe76ZeaZD1B
+QtXVUF2Obh+01CVu50rhmuWoXUn+prFd+d+kEaqgAFKAlE8942lcjSHUjgl/sJv3TzRwc8oyX/k
+KTT2xPNzLYJQSxC5Oj7CQDdAQ+DB2IIDNJ4HY5ifAlA6G/Rgg35ilsPLRLOlu3QaBvX428UE49i
rbl3nLLxUAcTlUQMYs3/NskSp6Cx9pRBzZ5fcU1KpdmYi/QMffGgSJKUoTQUX4eS8X7VjpUcWuXd
qVhlMD/kbk1DQmm1mylEdeq3+6ClVyvtltCcXSiUubbZ7pD2ugcd2oaG+I7RsvRqA1K4KIH625uq
Ghh1UU4CJNHSEey8miDWvsEWk0cwFv4n9L9h2dMsodHIzbNPfLc8WSXFjtQfOA3awhTZWKuU9SER
U3BkdexCu+nv4QjvgEOnJKxQJ7F6jhXD9Qlu5c7GKGcs69Nkd3i1j/B37/VFL9vWYUPr8gHtdNx5
FFFk4Yg3C0BkCB6fy9zEtq45K70quAF0ZpIm2DJIgmsm0EQiZnxxPFQVGYQTIB7J/RcOXHgJCqoP
JBLUauWPC5s8tTVIgx36FGlGVqRCxXHQVzzo0ejFE+6SwtNZ4Q+34h2JcKvp+EDkoJCK7+Ui9bWe
ybHH8oEmxs/QZx+Jz9CC6qXLzEE4oeSoC02fYYUhwBTmj4qf7hjVFQAHuJGk//1qhaPRHkoHGd7L
/Nx84kLVswq7k//j5ZBDKq4UVHQmkEMHPGJbD+PrI06iXZk/0/LCc5khDNxGE2NsKUy83cFMtwKa
bC5vij7HjKMdFnD4IoV48vIG2o06Vgw1S+bU/DEdXS+zBR3U6nu3i5II19SDOwKSLu3YgHfrd9cH
0py5bcbd2mkjEliH/CQvV/RjLs6s2LaVPOCapRnCGnjQi0iA5ACe4urcGMzxM8xRK8RdAMf/OiCk
ZS4sZgdTb6EppciJGSpir2OuP7Vl0zrgV2hl/C+Ar0tbwZEA8nO+pU9Z5ezRpqZD+upqj6r+ZSkY
m0ympK4l7lEvzQrFivBsyoOmvw0el11xPciHM6YjFYKzWltYNR4c26/Owa77yrspMUjGZyx0Uss2
PsSRUtpcR0pql7bcf6SODEQ/+qVedEHS6fiYO6C8RRFa0RqahIjjBzvov6kgeFjSQElTuCXetgd+
BcM0gZbxAqvXE3Vd5dOC/X61mbnin7Lfpzo5/Nl1CdrzBoPcB3YiSYeSmmYIt4jb8k6+PqbO4BvG
9LYdRCfX/B3v5XygGzxp8bdKIntqbKNrhHPaWtJblKUC9AT1Q7elOcD5EF/NTTvgefA4DnVB2JZT
VM5IWV8SWO0WTU4PcyZc9fSf1th6WwHnUqA3UNF8/EITPOXX+rSVNoHdSEptb236gs0Bqm1gJqSL
cXBe1rpLsWEUXWnC30Ha5gSKSFhYyc08Lc4r0voOz3HQ4pPXt/hgbpo67OluXIidrbSz5shhu8hR
gmq8m1WwWmdLu/Ju25rFHYMQKMGpULqHAUo8G0TWMn9yZ7cJ1OtLR9p1EL1u5N3AF8uRWP8R5Zht
7Yw7ZYBSeZempUd8RQo02EbUgyyZwEMSM3hXr9Vtch1I/JNBvGKkMZUJt+/9mzuz4Pf4/tSHDlFx
/RHZE9ACAnqrHk53O7QVFXLHV3tN9SWiPD1L0CenHXkgDz7tugadG920VNChGpjv0fDTOQMY5nJD
UXoVos3LzyL4Jj4Fz+SRN0dbQAyXabOoJAzz5tcKSuCtmtrauLfYJ2pDm6xKCcKuH+9X4EF86RdP
OCOulrNt8iJ9Ef2nbfB/MY3dR2jRuPBdFdMG7yzSt4lfLtEYlXWSQcJ+ffubjU324/gMBMYMuFrv
xDaVHc932s+xbLX1yd7OYyFxGo7Oxx902J2EzT/rWZWcfOdmZ9xJWtLZHwkWp7q5zXqseXBNNpDD
BW392HenulillOzgr0U2VAfRePSqiqAzC8TRRZirMUCkFapxF6edv4QsXRnLTBG+LMzor/2OIBxs
+73Ghlqf8bqFBCxgAhrk10Q1JQ3i110a7jCipxNF4yANdoj0YXMnCNknkzWvyoihsV4wQoeLhQNL
Yls1uey6uGZJ2CG0EIe4MqEks/OiX2KDtDfYe9j5WVwDQ9brYuiBgQMu82dRLODNAPVoSpQsT+cD
M8GnlzDfOi2aEYkZWHfGDV7cZpYWmbWt33ow4rW0XckM7nBLwKAXAVcmtj2SpzcBLBchGYGrxzt9
BlguwUGFceimvPXF7wz0X2ySp3YBJrhfrOgRj0U1z5bGlO7WOdkY916UvSoATkTdZjR3sTMLw0y5
ffiKXAMJRLpiSC0RUJAOBsTX4l0ieUlAUW7pXcSe9jO6hixxSE4pyJ4RRSvjwePlq7cDEOCRJsZc
pP8x5rN4R1xJ8jbkoxEqTGKx3Tpb/kSLTMxC+rp1aH3P0NVTA9IUJm9wsp61vKb1GZYiOB+ezKWb
JpllrSXJpDVM14N2BpVs4mX157dB86lM3eDF6/8DES6iBq8SB6uObtZceu0WeZqeI9oIKP+McPCN
9MbX8StpUPAOo6Wzbm8gFixnWTMj08rf0kUr93FwIkRyjPc/8VgKFNX7Cc/ddQY84cY7iMr52+Hu
rN3/cg7uoINog67O0twVKSCgiQtqwYAPet5U2KPVUgJURJzb6CS8K2QJeXoBtfFxSFJ59FnynOJV
M0awLHLnL88SF8x516LaK0HE/plLUg4aU3Cf9P1EG5wm/7udSSZ2ocvr39nNmF5dIMOdmhCfmsfC
2EyI/Y3E3i/w+zYpWsSTnGTizS9zoK2u0sA1ooIVfgPEYz9TJ5sKLd47XDyekKXzOMt6tiW95IXk
qlCEjveA30AaeHijWbfYFVuV9ve64niOu/mpJotAQOipqZMWyP+hupI1PiPLii08irEsGq2q9moP
Vm4vjnMhXy0TPO4L4BmX61rWuA4wPUdIpAFfmWgzKpNPHb3w9WTmocabmTYSpfxqE7AcnOV9er1r
9E7/Ti46f/wGI2Bofcqwjc9hYChuU3JOG6eYZSkoygXE67319kitv7RPRTJieBjUN+5GaVzL4fCH
xR2MOcw5xgzBbPwPkMTIBJKAizA2pxhF8favs8kbHzRsc2BFsHuKiOXAY6NepafBqyGgwNHeDRao
/xvV5Npjf34LFz5rUMlbuF3Pe6i+9/4pltFl0ZqaAS6GhpOJyE4bdXDbq2GhE+9j1Tf9nLLO4sgn
xPsBAIN8jJZj+lXj7/sox2+132GTvNTwd0hF+KScANPIfbGykjBbHZODLcQQC5d6CooF8CeYlo6N
9QBDpoBPSC5yLj+q8qeYAWLhnQFLTJoAJIYED9siyuG8zRH/5Jb7vA7I2p+RZmCMp7HQBk8ZrJs0
DYG+afB13oKdF8gEUhVzoKWoFUfJVqSwYvQttolQxxMhjVsiwxKRpPQskslE8xoVdL+flPznf5f+
ZkcHiBVRUqJg++2Y83CLXHj1kvoWcIlZFjOIMNYwgYxxrNvnTQMt2vMmaSeS32qDONDqGeZIT2DX
ewKIMjIqjzFqxspSNKiIvbNWLkJ3A1YWOqV3qs+hpBJ2VtxrqEwfr0Gwf+IFKKYsBsiV00qGeoz/
aCRnm123X3emHRRmpJ4FWekm9sFPZ0Y3OGUHLzaTEzvjEoD68BuvctEIOaGRPegwdBCaQtarMBYu
2sYXEP9KunFDKk0Kze+Mkyr9L3ZrcdESia+kN4XS23EkLWaXKOpvsniKvaWWRgcgUIU8IT+mpsOV
t5mGtLbvTDK3z++wqeoP9VScAlYjK6/6BNYQXSoIPFxlijWOIUtkOEh0odbAducRf3pc0rjTiBle
h1DHof+AcM/sPGljRvOupIc9iwyF2L3C5E1ECI8rJG6uaa2YmkF4ICDTI/wptr94O6vCbiSznQ9d
ImxiKoD/k0JDhhlH+Pcf8mmOXRoaebsMkRfaEodeP4pljVQuQpDBFHvDVTSGLt/IR7eSMWLqnkon
5j1i04aIlIf4hXC9rjJgiGuqpe5M8vXsGrJiDuZ6BvPKDAgw84peYFwKmnUWevG8VU7GLElePsiG
oUeHpQ7p8IMLT0czGP8XfIotDctNwTUXM9B9LcNw3yfXXabeoBNC1wiAX5UUmxDJQHiVvaKGZRzP
0soZS9b7xf1h3T0Ji+y5uI4OOF0CrSE5NbIshd0Q9e1N7evU8UXCkPFJ0eFDLWviUs5mFPBIrgu7
PV5bnaSViQNdzodS63uecHd8rCjYZarPBE+z7IKa9E2F10/oe5lDihtQZ840ycixg85hKN0v05GB
Ga4wbmZwW10S3XzZJBmB8rlWQ9gtLl8XNYuOaGO4Rtho/iu9EkfYcrAMbB17ibu9gUWfeG9ZuR2V
I0b9HIYMew/D5WRiQmk7iKqYVUeO1rKXYu05fkes9d15wOwpmHBqecLd6ZH/Rh+pZZ4d16tpRcX4
+yCg5C6lytUpNg/oaBjbZZomKPkZmoh6NtVvUcuK52ttszdM17xDEfZ32X7SR8dBDOFRz+4DXzoa
FHhKWlELLMwjLlmW3cSovYlBlTOuro5tSyvjzP3SEkOQtNV6/j5UbUcn1uf2qeKQAAOgJib7L8zA
pKwzzUCRPROHyZ2kAdw2ORW37hSMXk5KFg+fgSBTGwmNrHZkHnNFsNtdHzTn4CdXaKq7ydoEl4Ii
qaPkn8g83+dJ0jYTWYhmXTZ7Y1MR3/v5D6l64wBzKdPTitR3ZsedcC4y2CLTDbL57kC9cwQgtXKo
gQrNRCt5Qlu5bjJvA39+vSrwlS6Hwhqh2ThcSvk8kAq7puufpnJ18BE8oS8ZLMcBqTpaBnc/WOEm
6hvCv2Ia0VkZ8urXMQh92esER10DtoP+AsBvH/v4YXK2/kiN6nQL/6x06tnqa4XEoS53APH+ORoG
kTQ0zu9hKanEUZQl1fr6bAy8gQKRTYIMyhh8VAx4OXiAmP/mJT+JV3iK26ySXHumqCMPBrBgb1H3
aHhHeM56A1TnfdetL9X6GP2tIF1O5XXt5Cy0niseypLf0TJLRGclpZcOqd7kNZwzTkGUlybjxHCq
3TXNtB3e8VwW12egygdjUCZ2ywcS3ryZqZFN/0SWw9UB+eGaGase8JZNXrmxOxbxFImBtUHyHU9k
Wzmr/2tQSBCxJCVJyNpaHdmPvuHkmrzD25S1NsxDFeMClQXEJX4/PQzBgHYxMSPjRi4j4k1YlgfJ
tPV/dszyPYLDNTW3UrKS/NasI7PcGBklATLJEBTzakREXKRhUum7Qv8mFV2b7mkLHEAwOwC77GyT
VIwd6kZRvXwaTUe4oyRadO+SQclO2QoZjyWRbHDEaOKYQwlvkz2A4LmetFJk5CIWiWZ3gA/Bi8Se
rOvy76s0gPrlT2A/R/EtMG8b8i7FdVi7tVrLwJHSEZvkJwJIA27ZT69l8vF6gE5AV9Brz3UEdNxb
V0HzxgFTbhWHgAp7ziEmW4zK3eOCswrRfozfnP0U3Mn4ojuanYcbTXf4I3t9164RYzOWHvNvMbc8
C+rpxaNDZO7uvve4+BYxGT0e/V0PBTLxTY04ylNS3nepqE/ORU61/m7RXpnnjKENfBmNf44bUbVG
7e+O+On5hBeNfQxwU+b2qeuEx88D5FC1iRRn8y41syajmWCMmdNcWoBueWOwvpMr6BVyvywRDDi+
XZUoPrEXjnet2D07MWcMRJv/oF3GBXXErTkehxzaTixRLHWKadjAULRhRf/p5BI3JA7F6CWlxZAv
r2SPETFu+K2+FEuYgIqkZWhZDKvBdJpbIMwynkwSV9n52LI7KRbON4StW5+gBQBrvZxlx3z416CF
F/iSn4fhS8T+sgLH9nViGlTG8Sv5oER4M66Y7cl/e+g0d8A2YDnAnQZt/QSofxmPx03DYd8Sy6J+
IHLjj+h2n8GDHQm6ZnfqZMsdTCdbheYIj6LILR4X/EaNPPODCwvLCq4ZFp77Rwu7vZHKRHQp2kGU
bIiPzL+hSaHgETl/FEjbdS0eh6+5tyS++5QYndh6KwjDbBc8jKEq5rWiuLSNYOaUCoppgSrEPuX8
7cWKBne0gjGp4Hcy/BJyo3lXQtRuQqHyV8BMrZ6caUCofpXBmcaMVBDYR7LOZ0b4fZZ6T4cWnm5z
zcf+z4TDphP+K/630OLObWhydj/L5eeBl57S03G5oAkSRbr4MraVWdeHO1cQ5IOesstWZ/aq3ts+
IGJQCHWdwNhlShPvI7XZwOxbc3aopzXpfBBxfKXyJk+FJmxMjnEZQ4N7OwsBc1qy61LfBytZtHqK
p/SM00bEyINTec985LPXDXhXmIFWc/bISfflMHcaAdZrhbRgF2LMvezDbELQgLN4Xe0OeWa/evU5
WjnZIYqcM8afhJcx3dn9H7p6O6oN+l3UagzmPXCiBixGiCkR04oh8E6Ma5giUHJDLAcgfpPGa2i1
5IdLAWBH2/2jcZxlL+fb053Eh6WymhtoWe4NRfvmCKYfqhrHjK6/KkTKSyzG26sKZ1d454e7Fhfd
SjdJ0/ST17v4DXlyT7/Pu0ZD1DWY9qE2RX2kBk5v/6k8v+oI/bgsCHNUo9i0BKjJuqx+jydRANbf
oMDRJFV5Lrni6JCp5yqodyZJQ56m6/iAAtcTDjo1pB4GcN9f60Jm150Uwpc/tEPZa6i112IC8eA7
7yGxKRCAKjWbw44WI1e17uus70SByWML650zcjqyl3NIWR8TYDSk4M2a+ij6jg1R8uUJrNPA0DjV
gXbd6umIKC1W4Au1W6eNSNtPj6WGuVDYhJGcrD5Lms+jIbpxBOWGiOHHMoUnBwLstWrJSNGxpzaq
sn/29nSYLEvc77xyfcFQTHgSjIGv3Kau3UeajmdwmMiTv8tRTBxrw/NByNeoWdCp0LF80aKcxUXS
xXUSADUnpIebSsh4KbGTZst/Zq5JaocJvUQbb+1PRfarQscCnW2ZL0sj8vMmGxDAKqNt+XTBjtEK
jggFPB6eNPElXQI6AkNhu/SrKUoBj5pLQddrWd5aDLXwfapX5Gz7sRRMSVLC5LyaOOYTbdgqEBPX
wNBKiIV8Y3WsnzBmQXoLZM4l4Ml3uZAEgnwoGR5/6c4czcXsxIqrjK7tqqvE1uai66qnbscpBFZn
6HD7TeHmyEKLUz2LTqh9TKiWO++3kwKmxrgUVLEvGg7HsmXgFUM0G3qZX+m3ri5FXFVlgPEoxss1
xgB3urNFjfnMJHQJ8Zb+lmvaPg9FSF9p/wUErBdr5/mRlhQS+QnEYKoTJ4Ps8bvEhkw7ex9GqE4H
zgFOs9ZmEI2mucqkac/0gQb434iCBi2X7pSuwqjW1RkJgoD/tGRCjp7oT7WL4FQwFzr7Ate4wZy3
JxuUNppCLJfKMKQi19tYX3DxzchsAzsFmyMWNcd8PmmnaBQxNnRvnP2LeVBGn7fvuT/BcIQ8//QI
Bed7laabNpCKzFUa0i3eU0vl/hx+WcPyyEKo8fMvXp14r+IC3RBZA8atThvjqj2GPrjQTsU+hgv5
HjWtavH4bOI1kzF2LhQYuLAeH7rszye6BYGbY+0evwcArncXGVHSWRhpAHBOlIRhy/uDb82+eBNa
fVw7/V8/dlxTGJ83B/5nIpNb+b2zktYz2scixjK3Ax+cP8WTqBj4CsCotopGbnsIVyiAxLzTBMGt
bu+fT7oJ+89YH1vkN+t4VRPr7nv3+TDUlBPZB22AD9X5bWn1vmm4eAEE98e0QE44GjuutW4rnmr+
P3Nf1GRpYpjZEWaby/h6jyCL0j0vuWJzdbCLN55s65cpPl0WevG4aEwe21BfqEYtUJNAbQ5Akcfs
+bg1hKP28FtJDm4nghiR5fqAMZ25BK+xJfZd7DQL8Ugha7C2kiejCr/ntF4p5hUSGeAGqcccv8f8
+CaDNMnZz1lLW1V4siuqre+YkiVxBJFN8vcfR/vEkERfJbakZZU3rTV+tOBKpwamu0spz+9idt8P
2f09XR5ZGHdRIPijUNbJZm3GNIQe41L2Dc+wFV7jpmltsqKxT3oNIpt/zbjg1UXyDFtaX14ArKRQ
P705WPcX1b6PurLc+7WQOAu6RZG+9R83lSr5IxzoP35lapL8+2F9DFT1nJaSgCdpvgucj/Ci4sUl
LTf4U/yn8P6qyynX4MPltLSwdo22xpWv2MpWVdpxPi5IR7B4H8GJ8JypK77Q0iT1+kn8r/X7GCIJ
TDvv7493/9LmbkqD8zbW92NtcYCHcDAS0GKdrNphX52nIKqJnBwrARspHjPMulKJwAXKdCKAjw4P
8xKICqhrQcQKK2mm/eRSYSC4cZokcVHjDWaHK1sIJjDkqq+57YeG8kAmTj+gmqerqo3HPfLcTWkg
uL8neX9n1iA3d2l3X9scVsUccTqmk0WH8Wn0RQjsx0Q17aWlMrlEp2CNnKKHZdkcS6QOfnLvK9PK
Py960O74cZ41KbBf+QjqFXHW3KYn0zq92sVHjY9JOO/JdJbyo4imvkEzlTX8u2IwZIhy57D00z/k
f8yStSFb8d3ee0NZvhl5wSIBgMPiWc9IPB53JICmVHQnRlHqyN8kym2/mdjSNxQlC4q3SL8cD1Nc
QEWKU6z2kqCWmNDxCMJbPXchhIOqNIOSnWIQ1tJUfZsNWqnOrX9iYPDrDDVXZ6vzml+z8QixLWSz
w1bLOMr01mQXiV76b9FtcD7HwzqvmiWYO8jr5IGU+AhCXSInE/NEgP17wctjMK8SThSR+z3R6TIe
LL9mHf+X/XeKpLmOo0pcLBcXmoRpawbJWYd8D+YYnGc0gAoJnyM+3cK/xFlKh9lh1azahWDc9663
YMyifVQQyvlEsmZUKojK8TSv94tt2rmt6mrfsFHyXftJAe3AFKKUZwbx5BwwHCnI780q4IMhZ3p3
4XHUvcdAaP6mUfkPgF1eGdPDsJaVsnQ0KJLhLT3YYt8hpDkuQyngEf7Gju6L+xbYev4d4lD1psSX
ZM/FcHYPMGezbjDOu8MD3MMxeIRaKzycvwzUJVskoL3HhjSbANzxKx8msjpwuPOL8CmkFIVZtkQi
6aQqqmUG1PWgzl5nvic16zdpRvbRtlnh8U07c/zUi1qVNUu+k2TlN1EIxxEOBu52u/tg42c3VVC2
l15fXIh7JhdAcFWS0vGEJNlbnq28v9aYmNl8DACfVJ7XzORZQ4/KCW2E2aaWTkwroiICIxLmhgW7
9VXbuLsrtiDrBzHpSm+ssCizfhxs1oCZ8bZtmaBRaYqFIkAevIIG04dh3EO1afc3SP3sXx17kZzo
oNsnNWoZj8Czp+9BfCDXd0vQSrn1tkHRXwtIKi2BI3u/GL0gMeLVaQ50O0+CbGUDRBCm2F7zV+aK
i+6AnblnGIHM8ueuCmVQdy9OvTzbcoF4dCBX6qWHrTH2Jv5j4wX9Pco7pAMSU+OLgMVx3SA4dg9z
+5sOzkRyNgA36vFBriCgxLM2HNhEF0fCaIlXMSgezszaj/BImgsxXnDJzmkSPD8QBk5h/x90wB8g
VHVCV2IRhwxvBiWuzwkzWwyFgdCr398AfFmlZZGdSgicGpN6Xwwz6fVfEK9479l3se0HzZsHO0MJ
aJcfoCre2ebYxuemTe3afcvrmg2J57hMjK65H0Po90Dc2LeJI1PsJ/nyi16+PM2XCsf35qi+GgyT
fn+MW+aUuEPHLdkwyYZlBOe6C9ckNAyGmwfqhcmm+KT/jROS9Xq+TB7PhKkXF66MtvY1uibv+noS
zJhKM4hWEesovdGRaWZUC7yvaJTu/UrIqIDX3ChRd4CJO1d6KgFrvqZMAABpmL3Lf2c4+9xaES48
miSvjC3B6WM2nsAOuwXT+0MzIO6yp7gDdh8VtW1MOSjz2G+gAT6yGUsHDzx7JUdC8quh7rRoOSQ0
FqJV5YInxYiDTQFa/1+gcPHcb7Kre8uoCegTFgVTCyyS/4hz7yfdRnxZJ4Om4TcB48eT9AhpKhZL
W13B3ICj9iqCZaKOh466X7BBcIP6BYdvrOO2phLwG7PeC5TRfT7CyApe4b3JZA79JI+w35u9V0k2
nTAiTXmO+7XCWS84Qt0GtuLdpZPRBfUC9hloU9/hM0pqdh5vfYIOrU7kLys9JGkBUppIxRAAlHEc
yTT9P/MnsQMG++VXbNDP+jxKj9KMFOv1Z3ACrHuyFIo+1etZbww5pYWAqy5KVC2FJwHlgpxir1SU
YRx2QdwcCfy6fz6hZoHeQeI+KgXQD98+Jx2C6YZwXk+plUUki+MA5MLkG2yXsI4XRoOIjXuoISE2
5xs9KE59euF8KZ+dEPc01xFfP0a2UEHKoJyyTOt6AFtaV6KfbfRQZz69Qx9t8e+ZF2WQ8zMnKjdm
vI38VCo/KiE7LNJS5aD8D8Cpm7oqSgjU6c3/pblEAXARRZGuQA/BnJJZcXfALJaDkcX/laA89Y53
DI4ltXmq3F+fa3US6sCJ74aElyVbhcb+6LgqdJ49DGNt3ezGckDqSomP8mcvHfjRnhhx7zXyaOYI
XRgpNYaVQNlqta/RUFBJ6WzfZKZK+TRLXHam65KDrm4vcw04jmyFb6eLrtF8cx1IYYaCKEDyqBdK
cenD4MdBBSrvX0oMz/nc3Q0125cyxPwjfE/Ey8V1FgIdwl9rLtGuyfVsUKWz4GLO0Zu+E8IETI1w
VA2JST/qtYnVh1JNv1FouN/9rfTxlH2VAEVfs1TdTqTSq+n5do5HBxD5lXsiV7wKuDOyZ3IuxMe4
TaBz+dOoqR5Jq8w3UlC/AirEMMZFdAy8oPAwP1oeevQyGGc4b+JKQ0My1fmHVSrn5BSJEEYlEdXc
NvkyhZwfQN5DM8Fg8BVg95dxbIL76UE5BSOR0ACCOTaGwIFelzviBg3rHNN/sqW9wioG5WnBLt0H
RWedF7IiRyi10JgxiqgiOOgob2r+CrZfp3hrMmynNLDAJGjG7wmVPKzUrCs1DsVXtL8ENmeZ9AUE
Ky/E6saDPCYhtz6qfSYNoq6xgUnHK/M5RIg6rIwyVYu1ooTGkqzXLSbXEBki3y+vVkd3+9VjIj4y
dXRiV5eOx5wP4JctEANnXKox2wninPDNgn73/SmoNINxD2fJg0wTJ7dvIxrHe2eZMVZyQ6dHdxxI
fx7NogPzsCOH0nwDxJwHAzVupZBrj6WfKj8zpiVBi/D5QWVGQ1BZ1gwzSnWtLIQETvwvCkikYSTS
yKLY724KCgT1PXLCoG6lV3cncvuCuWczCyUDWKzQ8vtNKjYpKqI/wxyobR+HPRLv68+YtufgITWA
v0QptAmrKo6Z6nd4hxdU2vS3asKh1a3TVQl530/v5UfZBnCgVc24Y0nNB3mzn2VmrRKjK19oVpLV
lVznIWLCWfJXVXtcXW8l83zOQw09UeKZIIB5JF65jG+5czzqDn5m7Jxc1eJQDesKWQaH/FForJNb
dcR1yZOLBA5j9ZIVHMQkQL5EHdZSHtk8jNGpQuyKQa+XDxvhP8+z0pqHY2pRvjp0lKAQ5yC5sMmu
4lqHKBPHhsKHGDjyc2gzxL1XKsQot9rx2kc4rSyzHKhr5b+pxygRtc+HMzcbZLggUfSbQNcNzDaS
Msc7t7qgZT72hRIaJBDIDg8HPda2hubbwBowzMN22c4l9QxVi5saNIBpMOqKhn6QA26kKQ9nb31/
0ospJgHL0YOlZ+S2XiWxgHnFSHL47MI5+K4qc/ZZbu0Ezv22cO4mbaj0lYZ2EaSsWkVIFLWKOg29
Z2pXiDankoawMb0Fd3O9ulc+zWvfG+8EhThwBRCJDkb/RuSiauEA3aaPOZfxypY2rUQzeRl3oYTp
D/5P8H0FtUCFANIeRZ7hk42VRoAwk5TlwlIiMjdcPRBQkj4QxWBSrCnVUErlSlWeJCYwfA8SHyKU
Pgycd9YUZXBCPmmIp7DiOkEfuPV8TIdb9k+jDiu7jbrk5rp03C/s00D2sCY4fGFfetwfLZXwYvBT
2K3MqxG67Vja62mVVogl0zUHkslS0znOGQqMHr6WDUcASQZqQR2ONrNDIAQzFKUUgvHAzyl/GOi6
MMrKSsduObOLLbXWtwgtavXMqWfSu+nOxuc1wYUeouTANuCRX00pqKSNye2dJ/ASIP1pX500Mks0
BZWmaWxm5DXgXkFLAc8gBGLqF2VHwxKdzdobHQB/MLvWJcdBt6YmyA26zayM79xOqwljYPvQ3Ujb
QiFVyfgoXE44+fS0MtRa+adr4SPGe6l8BLdhwqcxqgOQkaabFjD6QmJNgSZ4V4Cm935tCMHf6IP3
vYko5n6DX3GL0Ozwy8WletOopzPyKaGpl9RYQlzXwMX9wSjktlhvRipq9icJ9NvkI1p49FtNkb29
+KEUp6q840GQgsO+yKtRCFTz+LswxxdhLIXnN/AQ2DTYQm92SARpr18w+jJfrk9merL3zqgjk8By
P+BddWgW3/v50n+TwQY3uBbvEOUX/mn4/b3PBo9oBY82mIFp32LjliDRShrDnHANoRrE5WbQyc1S
09OZSbO1ywekcWIT/6yX11hJzhYr196pjT3sHcqhRVYhLM3fGGJ1Sm9NLNZSTmB7h4bYN1wZXnrM
/8fa7O9AIRSp3YHXU0dU3geECRDSunk2RTAzImNGw0m6tEWP++qRDKtJNhYUYXjPt+DreBaHPjQp
4BNuKOpZz2EPgL6EKt9oCp2ayH+6XxA4Bnhmpz7s9Evd1TiSoKOSo3NpWEi7XsdVQZAMfEqSabBJ
ZY+HpEjNFB0tlaVoNbICduGfgkQWRbGTdw+/X5n/76ho3zTEpNUixCbFHMHgf1sDW+udkKp1A02J
hSwjAY2c+hnWOpE2EYXjJx8uhg1P+iwADdwi4guG0XNqcizu/XaJL+T2Yf6wVCToco0geBSpUe3B
LrgOoNiTF24BAnVRVCrGlXNdmmM3MVONq+XT9UO0e167PQIE9qM4JUa/eu56QphzidMKiu1BKn1i
jdEXa8xWoB8rMW2K/Ik18m8KJXXg/iz1sQ+9NzeNL1Rdzh7uDNQ6mqGRGuzRCu1xWld5QbASlLYS
NDVNcRXt2cy8LQBKNbA0CpZGBSqI/q+++fqSFkQ9x1JbtVWiBXf4T9rRWKSlQy6FXgqcO/PXpz9+
HEG5BtSzVP9ZF/D1cwmdSc7cTsuW/pqd90d/Z8NYKblYY73fG6z4XgQ587HZxGg2yTImdKroQuZJ
8lIDt++VOQQKvClm2gne+WQEXVMAycTTX1c3d9bf1VjHav5+kZKMaytl96nk6mfVCPN+rCNCDa4U
5G1uCqvgfj+zBhWQrOBkb4u9ZW0wufCVtVdjHQn5Gri1EYjlx/l5DeyDKDVhrczlFhE7Crq4opYb
3zKZOW5xCVBasGyxPCKppldMNUaqmQmE2M/IJrRMVWWj0AkgDsSPL0DkuxnGb9S7dhrZT/FnNGB1
G+RHMHkGi7d1GhPmmrHrKeOj1Wmd2QLe6ilL+NLS2FVmhElP7PXMlhSgOa3pYiuXrsZ4VFTobPxA
NeR9WRQeI7zyRCWKx2euYljmidTMYhndciz94xAfPYnehNcGSOhNBZvASgjtQuD35IkrpfY/DLA+
ts3EDTXuAFpHeSekrqEi4A9nMfS4jeEtS8Vh1Igv0M/DFXOuFAAZ/JfinZILxpv6vuzsjk8BcdPd
rKjEXsPWqiCzGgdXhkS55+9DyT43nmuyBMgnnI16XgqpAPBYyfQLRaAbRfhwiSmvDfS/E5uVDi6o
GFhFbLRNXaevCzZOyAjrehaeLWLggtsNlNx0bZzyfJ8HwPeij+ofxTFReYxsjd4yD5ppeW/5kqnR
PHYSDPCYF1HQCccc2zNUJhH/zXrYkny8PI6ItSDV9E1zctxAu6SVMFjUo9YMn8smLS6v6y1CiI2v
fTsv0Dr4V+PlpfwYoRohQwuKAIlrIGV/h1PeR54LtokJrLBM0bxuW9Ogp+lYnzBPvS6kTTM7nzXY
NoqgYApq/CBmRLBs7KGJH9fRFk7VrY86fMW8kRiR31oSwPf5DUmGGIS1OffSUR402O6Qzg8OHfNz
vJlhxcqQiCeh/yfjvGUxXEd+OqULeeVSxAmnCdnopzgSstVEroEORcw/Ua1HOti8vGPBv/2ssNy3
OG8Hq7iEZRojIWKeLJJ5GKRIKX0aSnJwhQgc24y6bEsekuwwtB4EG5PYUBAf/PzQ6u6q6CNpZGUl
RsbFkEiKvxfoB7gnEqw4jDaQLHonwk2HOf0obvXSf+t8ZjWk7skSbVMjTRLGPbx6LbdHNWIkGgYm
zBW6yUtEulm+Maw3R5FRZXZSxsMFlYSLKMkMmMOaYVJ8OL7d3KXR/GiyPDKLNLFrEo5WGgg74iY0
vo8uyhozYYRoQ+9OAjpVHmk36MAEZlhB3haH8OtFysndyjJpb5ByUWEdsD/QfMGtPpRh/Ht1ZGbz
DY7ryO2H/CUdJSWQbIiWXkYj6IKAm6vgEu70ICV8lsgDzF0NyoUj6YTe9KF7rI7MIoYg3mSlDkKN
vrzth3dPNR2oYmoQkMdyvcjy6z44SxvjNdKBsmY5lHtKMYsGR/ThzUb1nFC3Gc7g+RiY6RHkEp/b
8Zfb7NTE9ezLyz7yo26l8HYOX1t/zQ0XtPLeKSto6dfPMY22z8Ks89rF5uQLXskSNLlwFyEAql28
hz9toLi7bvfNi17b70uhWyEUtPCFPZx8jOpo44TSZawFjjwb8uh/i+YCcj6HoVE2GvZCeOi8FFkl
/GKhyK8eMX6AP9PbxqXRqCm0GrqeHeSAZhmSjV9rAJgfKALhNsH0Z/wkspQ07l0mPu6BGUoSt23R
t3W4LbJ7hqJO70ed5axIE1r/5TCuVC6tFV9cwivCSkG9KGgATifpT3wW0d7qRIaf2XcFjlnL7hvK
5CAb9WFDXbtqvSvZ1OjdSUD2BLX41KVAwLEZFO6Qrw3lhN/z1wTShrnTSWWr5YqAsb/BhpPQikqR
CCYGgSppzav+IdNGpvqgaGgvtFc6dsr/41vXNL5uLyhvT+Sejs39dnhYl7dpYMd6t9nUgaxXLmUe
LPKISpC1t0HnSYnarYHIXjo8EMmxoIeVvFb+kEAEBk9pXc9QH/hGlAlM0Nft24ZDUBHNnHsCGfP4
Y0Bxm90UZGvgoE+s+c07Ck7DWb8UywCXt5mMvCBbTNlwtioxGeUwx+LWTDhC1vsugW6IHjrDOBTt
Jx035QagbzY5KbSqGC0AiA02qcOualAonuJpyYde4gM1umS0PUpbKtSU0DGlVvjMAbiiE6l1MRZJ
nDV4rAWdB1PrQekHs0TnVF2NAuhxgzOS9I8xFgKeDXdMMOim9ciUngyBbfgtR+veQWeB3ykqSeov
yNuc1atl8PiPdm7kqVHmCuktGyDZ3u6UG/1F9KpvCr/s2eUiJ2EQ+h+sG1ymInK8TrXiiZzC0bx3
WLvMmMUmI8TrGprefulgGlmjDE/3VUg6kQPVeqbZlTcoqWZOTLSyVCoZs6TfUfl61W03q4o9RfaQ
AT/eDWRZmMGcTuvo54GXsJWgMM+z3uxkkgFIES5HvFbrQC6Z8t/Icp9YEQyj1A7PfdSXO/szAveY
fkmgmOanOBUcenWgjAggKG9ccxsFdqH+yyjxZz4Ug30y7GDP9kaE0/48XNATvEk/UJ9XE9qCoSf7
IFLg0Ymu0u9HMtajJLCtIanWqdCRw/jX/yusJINr0nX+KSAxwPz4eLesXHazUchFC0kEMmyqmXdJ
uDrG3aFDL+PTsz05Rr3FuRCbGsc3fK9pyhx50QCQEmhEJ8vbaTP4n7ttkAJ/xYqrwuLf0XtQDI7g
KJDHNu2TiYn3deTN3PQlVcQBDpDByxqzcCjS0Kqad7/2pnm6DjZ9GFHpER6JJ7/SonQcN1NWNLJf
g11YCfXm14VF1YYDKOw/KiTH6dsn2UOWzSydQoG0KcUTOk19xKqIbkjOF2KyB4yUfiouYQKA2wAb
N+Ko5CqAjXKEmkOYzLjMldIKJRqlontK1AbeVeT7qHzC2nc0ABCLRY2BgCTb1nWSJpvtMxxqm/Fb
tzaetN2BjrAZnh+Zc5KfENFeiGhyCaIYlx7jVwSrWSllFNAL+setHFLJzb0laIalVItliH5cHzbd
Z0HuwbPoAmsduBjNSRilWYtxZGGmYJqNBdjeUtluL2gjH0YeLXFM2api+hFfJtpyh+7zfoY4urly
TZsw7AwvjDG6bAWlZ9Gm2Y0fa9/oCxRsym1A4tdt9ye9YcsojPJcsXdIXBedMXwXxKfo9/Fgc9G5
M9xgaHArJPtcohgcBajRTSNvhqxvDqd8SoiCVjB9XEsjHn0F92ZyaNJQQFgRmh8cYyHywfqV8n8F
y1OFkERqJFTJT8rJzRM+yCYNYvhFP6WzXIXOiBK1KOlyliuzvc7elJoD0njDugqS1BDvpiGAy2t0
HypKwlNKK3/hwAemoMOIpn5TE7vi641sX8QlD256PMLBPhpvPkPWvOENZ16ZCqKr7aoUodGAQRO4
+Hdt0OekZl5UfGQk4JKc3nQ+KQXr0036gMdn2xgEUMkpEJCXDCZDyGYEaGUcLWO1+N/0gehH6eYg
LnZi2HhyiKYhJH6uds4j95S9Cqf6VR//sTltnVoM8F/n8eqOeSa42sNKlM4NydAiOf48mywY26Ui
BXz4wrWux/kutjlKKj+Y3idq2KEcf0FBot7q1dMuOUOqyj/BB3V3ftxZzdhLdywHJKgMpXwgNg2Z
ChhiRvEOwvhvEVsMwqPNfX9Y3LQrrDBSaPWuFe8tbIvd8Y0Goh1osi2Z3yZAFDsUTCNms6fPIcgR
LOcUav6aeV9UXAnJGrGlFTjdRixRvwl9Xmr6oXwbiYD4r0g6OPJuIJJloyazqFKRTngGe1+5lWhn
6dZhhQzpnVZFa3kEprYsGGQFcxHRf+Rg7qqcTobWP7B4M4gBa9AjiJnZTa1djhayS+HvM7Q8dkXx
4B4+BLnPJTahlSD8Hq2n/2oV29TTa8T1Cm+2FdmoA14NTcyb6HZXetgC1VLZbb8QX7JV/cJzvfyB
1hTxYrN03o0b5SYgWbG/y/kwtmyIVKifWcUsayye8nLL16QteVlB8W2OtCf8dyVFJC0jMP4dpqIK
jriJEmYF4Hk/CvHKTfO1Oid2a2Q/AKmmoMF+JMwlq4hcr6yfFvsLBq4jAjSYOQnz1PLKho3nErDx
v7/nPrLNnhDWir2suS01hLe82RLMJe1eIqswYz86xwCzzaAqoAQtuDek3xU3FZJeCz4Xrfuz31KG
yiSMBbpLcKZknsBMsJG9qTQbP/e72rgPPjIITzsjtaHX0ghYXj0v7099iRy9R/yGAdLlJ7kHnxvZ
JQ6qB7YxEYLn/eaJi60P4ZsNughtZyw7YAjTpwt0efGO/cUaTlmO503hD9GVc0mK8F1tpx7QROCN
ajH/+teA+Uv4kIVCdMGkU0iiem1rI8nQS096tYo3ScRUQex4jgIl0y26R42KuD1BHCvvq2S1hzWy
PuPTxAMh/fq4ZMrzW3/B9oOmNPiCKyn01NjaLOojAIX2T3DIJoKfRIEAK18RrNXer/1+u4OreGw6
RzbiriVW/zvaUu2POUhoVFBqFgt+R167+3UXfE9jccRDfYVBfPwF8naLXNxwnNT9WxQogET0sA6a
JVqwoOItyXVSoxr5AxLhG/rrd2VkFfiNOIB2dWS2bALxv/E8yZ2p0NnDzsO+uHojp2IKfUQbOhg4
uZk4KSE1dcKwje1oyFD6EtXcixG8a0VA+5YeGViqYZriUrzAs9z/V6K4XibMc3XrbNylAzusQ6yv
az1wNzMwx0t6dF0fEhOi8+xdX566yQB/j1s2qOlnf9qOrMy/bAU9XM0H0l3ilnv9e6kfK9QfqAOk
WClNw2JAluCOdMvlHZor0iG987HF3go3u4GBZe4qa7GxsH+hNcRwwWVMDEeC07QNLgmpnrUYB3KG
PRumDFPp+oh9/IM6bA5mowhibCFbVZyoU+38YyUolRMJD/E5fPIz+vkCEpgfmuyGEjUJsVH0/E5Y
4tga/H9zIy/Bqh1czbSz0Gy2SSzYd+97D4jgqChZVDta3t8ouMCnCKPmYyo2IPzipr09EUXD6Z4+
NFXlEJQACgAUTrWS6MAicjds/LBSHYlG7LR4V3JJjyi+DiP2IzAqYz21PAc5+W/uyHhnglfyZCAw
uO6U3+h1+kPQOpnrZTdWZXDYnbfDTj+YMsWeqMX0HdqXEYVYR66mKR8Sv8kpnBk5OdMVG9i6Lb2v
FFn3ydG+KBzYMScZB/Ln470jp1ZavcmIgTz+5DLKFG/xNsQKvOzA1xth7pFsNy68hd8TrN4DZpKI
4C4oPUYDdPckDNXbE8Kt7YI3QtUfaNo4YxFLLrs16aJ4NIgB7F3KQ5ZRZ0fJklbhodGnqh834w0c
t7XQPUYAG1SmrVosrupJzJ4sWNq9jGbKW4hRiEsrn4Llp3AOz8vmaGVBaPmIUvBh9qARnzmYwOLb
h9oWT7dbUgtifXY8BDKAGhdhqymrR5PiJbBGB4vSS/V0Z1Vov2j6lPntaRpGlBk97ECyYA+UCas+
YdMg+QWJlS6tPfB4NkITX5NkNroKqFQ/32OphfBHsj04jkd4AFH304HYZfQqkk8Wyxz1wtZ03/Rj
IFWVoxrgMJkacBkEN+40NOACRQX8ftAahYWZcbd6OQVyO3B0wFrDe0rUPhoIBA04l34+TmRrMGGu
IH+grpcXzOCBtrynUChNUU6KkCKMM+8upch4K0GGn8jFiYapVEcEY1xS74TX4uTHWsYVRDi4vsW3
Lw5dsrJmMjdts/al/CG1yO8iADQEgrRm/ZuI8U+CqNfGIZwRObgRc1r0WvQAbxHyVcdcMOJvgUnx
7yhiVAHtWaLyMFghgefSvdB1Owrp5Qm18BYQvPUz9whtIUScdSuBxWYfZDZcsL7HCXXbvz30LICJ
S90ozBDR7zpsDz5C1jCZty2qQ8jOXTFeLw8G1+S+wo1OuKkrKHPfIs5uYq0sx5UXwlG/RFQTVhgP
QX80ubC2FohkhPXKap6AjBgNkAE6lR6U2NdiI4HUgP0ZBu48us6QzTFFvoR+SeIw1OUGy65Nei3t
OUgw7UA2BF0PP0g7MgRXqq3AZP0mZUfXSIzkqmVWeoCaQuk51e9gVwCuPN4EYTyP8Qnsdo/R7Msr
bEWYisxcupnikf5ty4GT0US5258lsO8dg73wVwZnPVk7wlUPSlxDfDrYd9RzL4pQ4FPK9oHXOOfH
KOyQO+yLCDFrHWibr9RaisrSQUQKY74OctGFTAxT5BR5HpN8+ziA/pMQvO/tSbsVhWu3tVRAe8Rn
8sGM4Soabi7Rl/MEHYI5GT/NKTFW0+z0isUvvlpuZ6Vy4zAgeJlVOb9anYCuF/uDQE269jsYcnc+
LpbqZsYV1WUvOd+rN0TFm7aqInVNbxPhCmojiLqvnPqpj2bOxNkNzG+Giln3yj+hUG4t9v413bu/
h2y4EZMnNq6Lo1k/GFjikd2V9rEo9g4UgHLzcUj6PIDK1bQGCTnlZF2OBQzaNSd+cvWrF+OuPP+f
/KWuhLMRWBpb7MQEKFKpUu640kh227mnqgs7HKf0JBf5NADg22T5+2G9kUGRbbxRu70Q2o1/5H3Z
cX/lSrafi9pwn5xXDHQRD+BCEgKe/lU85ODrQsqgpwVJVr6GiIDydC1aKXxGN4i+7ksxBnYZLt51
hBIpqP+57CNtYoiUbiAAwY76oc/FfiGDXBcGZavia4oOKS+B7lQYDERwLHUoaLXYlKrgbeaKzDdv
tvpHUacFrGvJrvqhlRtSzosBXAPUK76lbNUIZn2nco7wvsye1ln/1vf3XH5dm5tXEIj9jAmeK/ao
SeYy/OGyUrOSoAMcalXou6GZl3bAkIUjDabX6qTbDtKUAuOuxSFb0AISGosgCTxVx2bq5ZwspY4W
jf87oMUg75l3grdUgfPFW518APQ4s5H1+mbXy2GWkkCPT+veu1fvxB9ibCCWiHFod5E0xK3+hcg7
Z1lOpgaZDBfOkqe05Gk11bBmhuWbw1I9V7EhDLisJennA68n2mW2L5V85uLkdRnCdcs65LbqEJWL
6u2pMRudOcJKleH6vIZI33rb1lqxMvU2fkldJhcdmd+1NKctZxEFwku5dMz2kTd+mBuVUx9p5IcO
rWd+PKSiqZm/QUQCemJy2Amdw+SvyND3MVyHKPJ/PrJeIBwS+Lovqakfe3zXfKZNBIbaUyRZS8nq
O1A39C2VJXn460mGTV13/WsoGbO1MfVq2YJ7M9CHjJ7M5SM/kt174a2fLMG7aAk0yZjABuM75znT
dxr5jFVAfkCurNeaS8lvA8t2OUR6wiRfFHKaQq9krGlQkHhlcjmELRJBoMZ/EnFo6t0pHsGXH6GR
Q5K6SsUUQWA/RKSiuGb+2lF907fe25DU9vR/tYt4GVW75WfIgn3Yh7GCNCM4XrZ5muyer5j7AO6J
immF13j4dRjN0Veg7GHb0vM14Rijd6oPQpVKnKFZ6RSjIFfEDUNQ4fu3mf2KyOBmlRPFokr1WpyZ
O51OBOGqm2paM3FI3Y2tCRNl8Jtdqly3Lj81yufxepTZeP5qw4PFuyiDUV8ESQMZYHI9G+fgqzbd
xADSkOFCapYND5ii6QCj2SGGYtKTqBMNuWrSnOdFKCVj6faLSoZTYJQHjxrNWh9kFOv7OwX86LDT
FpqOPUCN6aPFEZQvXQUbN/81BGDrdfi8LiWfVEA0idW1LTuTYdPp+C5IxY72HGilI/cq7PW6jlXg
NIQOI7uvYCLKs0DLmkjtmTsGon+xlbJGmMn+I8TpQmz6ZiSET7ArrPU+amH3ZwjFCrNJc8vO7zWw
1LrCtYsi50tcUX+naLZcnwWHICYcCvCvOqiOw8Y46Hi/HlAAdVzmENlrO2rpFBQevM1B5YfDDag4
RqZmwJ3Kk2O6gWIHHMyenYEpObl9obWGQh/oVHvXyDA8OCUM+zEiD+5rLchvrBQi0A1RbiWNQ4f6
p6rweLCceRasjtH/Lo0uxTd1lpS34nM+sJTOG3rX1Zo+8JHqAT84tN1VUl8uiNvCcDMavOoH9ZYh
xwofLAX92cYYLKTJrLOIDijYFqYWCfhmo8jzMAj429u7d1ugKeO30h3y+D2V6XUbUSjF27OZQOyb
h94YpWzQs2QYp5mZXQHAGfradBey58ddlUOpQSqxnHun41p9Prk+xk/iX0vjneaMJBo5xWFp4N/x
pS/f2ai8tbq3j1GG2ebJhprgluvR5u+cChxCoWC77b3Gxmy1AdXTfGXCAJ09JwyWghMC24eupB5L
8xhrt9umdJ4w1bZWsoVv5eFlkjaFW3JuGztut2tjVXDR5YL6se/AsgFMIhWv5q3n0J8UyIi+/+Dj
cvD78jFpPOswyzvftkrF1quNXfXdPVVznF2AkrhHHTmfCBqLXiwRnyd/r5/pM8GFeeVDdzc17ye4
J6Hw8YWfSr9gx0IC8p7MGntJDWmT+FP74bwB2fGH7bk9XkAjGCBZPmZ5DBK4k3ff0+jW4O2Xxoo+
JFl9BuhKRp/aJZ7AtqytEUJYz3FkbTRW9jGh1Vr8q7wE7D/C7x7b2VFbWZzkrZrFQcahJ9ArBpF/
etYv2DFnf06lEJ1UEnsj/03iwRbmW6YQBfpo0cRJsLcAUfLRMjkxqSMoq378lD/doEY6+EJh78d6
Hw9D5kdUlE4Y2VvgGBnf0RDVpiZZkTBeYD6KrEVgBCohU7Imo3G6gIPE9dqQSugu/7yYubWN6UQX
bhz5qxKkkLxEIcZIlZXiEpktGQlSMC9LuR7nflWbAjSttw+eyuQZ+NN77sy/R38rgG9BE3BvGj6d
nfESDZc7H32EcMRFPz8Sn7snXA+nMJa35Tz4CJ2QclzmKa6Vmwn5yqans9s0G+Wlph8bmM/raFUb
70J8IPtDwblYeT4l1HqKanC8OLRWIOAMoU7Sz5QprTTPvD81syB3zjS19BMDZnn4oFFnl/41rbN8
v4u2ROY34t0UXGP8lqtDx4nxcOt+2pMmrTt9qCpLZHkHe9MPA3sH6EzqoPjhDoz7MhR1qMgPio3R
oB052oGRBesy5R0SLkYccns9VorMepiM1fl5OsslVtJq0p1bjBnn8KGP4338iu7HREeExbvwq7L6
D24F44cm7E7dDWldrEkaPJQWZi4utgeJge/g5Vmq6NUZ4WLOQFk31kDrVMf027W8DVUBsYQYJHSl
6YpvHMPreqFxvA/VdbFxBd1Gg+hrsyXQNEFxTWNBFUXH4ectdvE/OL8SDSso/xNAMffOhSD4jJaF
d8mdziNa8IRKm8UF0J5i6AfkEjgHMYu578v/NpMPNN5N28KIV5dPhB3D/+4t5JQ3b/gcQG+8dk1Q
HIPu8JmjLXhrw4Suid3HzHlbR2Hhnx1vQyhbRzoGJ7Cnza4On7VOHPT5ECgyatMmJMhEQJkhwKKH
ABcDa5cEoxfgpo/4pau+c1+6c/SIYDkiew6euMIq8jf/iIZp8xZvoL52IHUXHujHwvIBDDgwJ6OA
a54CHqI5nZZRq3m7fdBK2f0yb+9e/49mNJldr2um41HtNrdq11FE7bIoHufL0+VQabAvQ0YLlb3g
b9InuvC1/61pnGaAgueEBzQcDhwLN3tkOx8aqHf5v0bxr+wDO0tKAg4zk+G/2VMPmOQebeKtzHCy
BmEj7jyw5re0CNJ8/8pfd32C+BZb5HmOPthMUbUyNsanGQcFdY07oKG7k8PrWMKE8+J+MDRH0pro
IrCUcP89MMuQfasTHiVKYisuEusB5TjauyPXo47e3wIkaqwzJdRSPMYK++AtEl8iBaiZZvdg3HMY
PwaV4Ey9I56xptAkV74gvbpOx6gRcxitcjJYNpgR3qYAkLQPrCcdP4L9vaTQufrkMqPNfea8wu2o
T6JnM+ILcpMwmKY0y01ZHYHILwNEWGbhgTCRTBSndHJIaw3HadmVASkkSHb8Ni+6LQm24qtrpz8+
whSnAnBAzPxPtfK4WorB+2O8t9z+G0dkQSd1mz+tlXojLz3Ye8RmmYM/O7Oek3Kt9MecjNyKLYJb
IxKOuqni8mqXzKPH2wccUrkl4vctAYQxmMYIHEiCoY7/1IcxMNJ6tqxj0imRlcIwGv2KP/DVH3K1
X6o4lwoIkz1zX1gdND4ytD8C482+EmKGOO6yLrDBvJ1k1AOSZFvKPQ+vnzXQlrEAO3XB7DT/BEpa
ZmDn1Y9HQtsJhyShyRLSsf6ZpMbsGf/vYBKJQsx9SYuy9KXJp+6vv10rvEKRvRyUTNdmC205oTg1
zvH4EqjY5tYUg5X2+M8PsbUP54jLBqG6ou7Dmp1hZzf/6fnPgw9TCyAjz5g473LphrJRWiro+bU5
XOBLvJPX4xYkc2FLEiZ1VpUhwG+QgU438JnRt+vD21k9QuUs6jtw559xaV45ov4pOwfMDRMq1kEU
DckCZPx6pDenTRs65gHGOGbuFbtSFpTszAxoOKudQE6y7wUH80sQk4LJc8FwI8KAeaPtxYQQw+fb
8oCw0V9bGv5FvejaV+JohkaS518aWPDAUcQNIOr2XgaSDupy7onV7SS2Wl097aggEwIqRhJEDXKM
J4UMv4QrH4UT5aSNl4qFF4sboAxvJUMM7dUrqU8Ul6bvmo37MmeIMNbuOqQoWrnlRc6pyzRwsMW6
POYMpMaj5E6hxcdi4K3GwQq+9iJEvBfLLZ3M12gXbOeKP9Sv6lftngJoT+oxC6JW9mcXGIwrFlSA
vZ5MwklGgxhS+zGWg6L28baNSMeOLdJFsvrD+V7y2LXEHe5OK09lpN4l8DMZhoK0vD1vzKEFZYX9
DEP4NrrDgQb5bYTeUBVmV/QcxBXWtCfpweer4lkMDFzmpVWt07zkGN21nrKr1LaLVG8o28A62ag+
Un5iFxsVq+/3RTbLO+deVtuFHrVk2dNW7/KlMQmEnSzTgHm8NO53P8FAhJsjKQlZAEXWU8aO8XG7
aeJFlEu9BHUFxfzaWzBbid0vVglQqor+AY6lQCX3ct4IuZacJZypCAqijcL0YeJCZg2BxGV4bgwe
D16ljxrvHxzZFKcubotHjRQUbvXgK3/v9bdPUzgP8J0BW+WawrJOPzKzQVaLVoVDpb0tuNy148yv
IfeZAJ0m0ztuYUSdqblDTX3WGnSSkUnCTQUeKBCuse34txasZoNX1HOXa5dj+HSoFMWatjskMFgE
qnhB1MI0Rn1gStj9xTx7F7pSeq/6iZVXL9Bre9zrfk71PkH0i4Mkp9ogJOD61JPOT60T8N0Y4VZo
TttK53EGU51cD5iYDrs414vM2tDZXJL4mrSPE8/l3Gd1wdMr54Gbjk1yK7KK+eSeMldF9oRxTbzD
yeCCCOhI5Q9bGk9qo/UWUPMXhSZNAJ8e7/Z4DHx6J8Kz1yZMlYo+eTU0RHkEoQt9QK46hZKtGJj1
NofPm7br6MzBG6lNrlDndvHU/Skfvjmxp8pXAZqmrq3qPhy3vFVOU+i9MwMZu0BQqQpexfLodHlv
+3o2Ze/T68oo137uHKEwOfyDvolQjn6eZRXHBfui/ByugjpifGbzfyDMd2aChifQE8XZEbE3hMcY
ySBuOyI4T3a4vxdWqXKyM4oZ/9DWHdKBa2yjNI8jSg1o56vw1brKisDccFyii9fe6uosmfCYe+TN
CK6RdaDwWr/O10uqJTZBj+WosXri6cuONEt5lxlZD+GeQIdRGT19BQp8fktMcuOUaqfaybn3Js9H
OqVtApb2UqBL4F/J2CTjqMky/hg/MJz0nfV3KBSD25nuYZM75FsblQU2JLmlMYwRN3JpZ1m4pAt6
Z3Otj6eyUvY8Ry8Dgcz8G4cGM2b+HwwiMy2jhyS7qpkrIdTd7+8Ew1VWzAo7G8Fdl5miInGyVhpC
HQ/WyOIDyXqGNOuZR4yYplt2Vu8XH/76q/5RSxMyQfZM56OeQ9hYi6DDO0CpWjXosXlxTqAxVK2y
1Ttu2DuoSwTAbOVY2SMUIy4HezWLKhppEcqY8WtLycKIuyBGs/KrkTrbx05PnjifVTh0WRvL8i/O
InRKR0ggFMlvcWNTfEnRp4a8FnJNui1kvVQXw5EfLd3lif6ZVR5tqK9xpOCYCcrxfRGmcEqacwbi
sIrD0XMBw5kFMlV50DM3Vb+q7dJuF4zw+MoPnvm5RVXRwqWsxTJV8aF10QE4bb5pxRhWVMll5EFR
cD2LFgGi+zIIjuwFNaoAnvtpK0DSe1D7oLdrIRyTUTmvCaiRmCYN0mhBw5Kp7NUl3LmzShwtmuCl
82C4mBwx7c1M1IdI4mrzR1fPdtkkeg+HVFLVM2hBl4UJOFLqbF++eaYwkLlyhr7LYHvjyos8clKR
MQHrW9GjoZfzln1dz3PiTIiFfh3NCtQHNleUUqYZKTWhZg58EWVoC0fgDmiT7aU+uuw/jcfMtrbT
XhC4hYgs02BkrtgFhzoJ565VIOyC+pfwgDfOMGAIKbLBsmBEkIWxq8QgPm26Np7yt55RqcWRTjnP
vs5EC246Iq/yJOtgrKuPxVI+5vqO98eCdmMkUTkEtJUcKwuu9PVZslEya7LzjdIrFZNKVbRufPq5
Ref1iYc61mICHTSwBwroxacp+LGeptdgVpVgcRDQLeYtm8URxYaj9iaDv3LEMEbnvF5ea9Op1l9+
Z/3g1RjeQK5MXNYih0ibEGp6SrEgWxSqIB9GwrE2CndV/SYu5KNQNHzTl3PmTKndTe/LC2MHfUyo
WrjNwNxJ5Urch7mF8xOUXJeoONtkYnqjg+MAFLW8O61PQyGsXdH/ImT7LLWvAm/iGIu1IVacL8m4
GrQ4YxpGxZv6LqK+apz7uVt2WyQQ7nrS1yab4J6B8ACwb2MNJIWeu+TdblJwnUYEaB3pnyXFoDkA
+3Ff+DBghtETG3Lin+tP/4hZIEdZ1HBRP1sQjWtRPCtYpd7ciBfJ2NY2HqE+SwHy+EKEi1Ct5k3J
LZubU+Rvwr6zsYpuKS6OCPIhkK4qVwdRbRxb5j4GvjmXNnq8e01hKduIvirugtBUE1sK6zYiJ5AL
dFLPz2vN5tdIS/wRVF1L7gVL+jvWimQOPyQatTzlNaAhpix5IJLUZmviaedFB4VcJ9ZWZZHnmdxh
hGg/ba0pG8hSNF9tCNRHeNSofg1nMJLlN0Xp4/XooHqPw6+Y+en3moe7C/90LXp4AKa3ys6NHxBc
uRuK4/kuXiczrl1TMArKC2ZtS2jhOqDocOO8WhhA8wUeTLpkhZkAOQ/41sxh3RTGOPnDpi/P9LkM
fFv4tV91dZJ1W3pw0ukYWIUq2nxv5A66v+PqUBI7b4Mbw3zOJD+tAkua7O8V9CXHF2YbpgnPp/kw
Kb1lMAc9x4HpWb4nWtn1rYTCHj4hYJ2YjNWEMEX8qVUZqiJqghca4jnnvAqZM0HL4D49xwKS6eEu
VTEdwrdpckVoTV4ZzWls1LKLdnzH5Zl6Y8o20YLYtjDxK35UTwQehi+UOTQXKVBQJ9Sj3UWEE0UB
dD8OodtkJecSDYs6ohHDFAHZA7nw4/NpAdhWUYZ7w3YDs+2mVryv24apxZ6D7qTvz59SsTvw88vh
3dlmXuDaSHzKZyV5Ukd12uYyt3i+sOk2uub+ZR8VQL9Fsl+PzbJNVtMB4B9B2CCEihkZD1X2JvSh
5g0Mkr07OfRfBXovmq0xZ2eBhCoap6guMWPHe5BQtNNVZqbbPiFR/TymbL5g5gvqiSeJy+pMCoaq
jpO7mq1KrkyB5cGIWyceBHONthp3X6p7V0dxw1gwvGeFMsNgCe2IayADrLAZnDJG+oR5LyihgloV
AcGV3bZTsYG5C4bIvIqMDM6X7QT1GZzeGLuKUnkkxJ3CVpnaJfnjSpOPaeFM7UMu17QC4J2fhy81
KkjiX9E3TwysLPimj9HD/rh+aNNFFcqBrTt5h+FTmkafUrqY0OW65hxhGQzAMsEzVFAxlvlvNPjx
uRw8kjnOqWTeOYr9sttvF8IeO0YPPx60B/3rvZJF2XHEpWUuX/JtDckM5PpXlAGcF5IZ1c9e5uG5
CO5kN2sI/jrXpjKIBBwHqmz5fkK9KKGOGHeTY/QNPSMpfm7d2XEt5E4sWCaC8/0AYMp79q5CkUvf
oOiRdk8IeeDfoEugOLa8dt7qTavSA8jxxENuRHfs4R0MlHndL+1HX066EIDdQcdyVVUqBx2HKWhY
j4ppwM3mRhpH4+IHqzsc+367W6FO34GD7HIUqooHOgB/0u8aQEhrS4THXflX4CKS+qA4r/f/BkOr
nsOxxLGVF+OldBIi+RusTUTqm3eZ+ohYCgX6ctrBYkz7YijMk2Ls+nuYr+vbMlzxu4FLdovpbqWk
hctI1XjX05O+UISCP0lo/YskEBp3BctM/EPeBoQfwW5wV5ZzM3nFU3hQ9h/pAsSIWNwKNFFnmLdz
xwfM0KNxiN4tIq36FKlnCgljcy+jf6y3pzfkmsan5TFKo8TeGwG9WqSiQydJkzC0oxV/WjXwtXbT
wFBaL1EFw1VjqKZy+xs9mxTkUgyqwLIUFaWGjiYeZeN/Ui9HW135cigDAvm/WDQ7z8KuK4zMbC0e
ESEZ42FsvoQT3ugoUjBnzzzaej/hjeuwbv1Y/0T7dJDwemiwMka0k5hwDBQ04kcyRrzM8+e9YtVe
kXkEFKX+gPC8r/xNT/KreIjoidqTndUx964nmYahnUTXp6qu9peHu7sX/x/WrbnPgGD2LidgcoJ7
g6v9FQa50QR5yd4xRBVfntASmMrVe8/QAL0BdUaqCp6MzhdCewtqe+WuE2OkkFGsEWwbOzu3fDBC
+GdYAc0aHULGJWSasWQwPZuLH1tN3crY504fe8tiBvxUitlTZ7G/jGd1tPN574p9ulp3dUJ0YB61
MpX2xCFUHmICUhph6c9t+H8o6bGtVkVHXdNvVAgs7pqiKndEk/XGgUC919Pwsuvvtc44ABH/URiW
jtMU9+1yFnAyDPkQViirXHGx/DbFLMyvZm1UAVTjVaf0hCKD272yWSB7RyyFQEeL9gh9BfYWwSNU
W4TX+k0+XquBosTn7cyU34OIQG+j3C6zjvx2+/cXhQSjuEqOsVCYaRcdBDxI5EXz/20PcRYBYtlX
qbF6NeijV0S8WN5w3nPbfb7cFEj/AGVVzGV9CdkCEsafUUfzH8ksdsS6pKcJjszSEBL+fQbUKh/Y
44THWlQKHL8cGgPLu6q5oo5nBoLyPXxfRbgWoeLFvAAicHHGwqlCn5ooDsVZC5/xnoGcV4OfXm3Z
3zUcZshpluE4tU1zD+C+k6lB8OnxtF4lJwTcVOOWOmooB9CqarBb2PzsfgkMxWZ5kWc/3iXYRgtY
+f58tI8X7LeOB8rAmBB5LjOjc8GARBLLI254bUep3fyemq8Wv1Vq3eSmYSu95W2vekWZxMJVo4bM
yzgBwv6JmhjVD3uW+Xx+8iWVVyof/isJlO5j4L0Tx0nJXhmBbuq+95Yss470m6Z51lLu7Q9L73ip
CouuNSBFvv6OkZouawJvxMnUdE5/9umxZu1sNbYbSnyvTl3MTzuLxKmBDIZZt43WXdcA6ILytA1O
gL1wc3yeb3BWIy4AC1cEM83/C65cKgUEVrf+fbtp1mu59MCnPZpdGP/fANtNxiOIuXq6LnLyZrCe
wEgoIHWw8niL7zmmww6R3FOLQrQAQD6r05Io05fZCjUnWNzT9Tv0Lr+AJf45e+pYuCr17dBmQ74q
bcpWGQD8ueWo9HljESiHlJsQFSBfCHNE67MscrsLnJ+TZ9h4cSjaJV5XRV3ZfkPGMaVkyJkZi8CF
Z3TLg8oa/crFR6Ah1+ecEYRUeMJ92Z7L4/fHpBl2omjjBx/qJZsYEWUt/0snWL7BcKpD/x4HLACd
3KJIFefCAs0ZDWLRg1BpaDZ+5KY/E5nESGBa/l2NZCrxlWfKT2AdXXs0ECf5nU8/tug6cVDCG2Nd
7/sWL7OYcqGITF2PQbM+qP/3JctS4gSKzjZhWAj1VEm7IN9nB1QKKD1tzvCXr7AW+u+AeEzCLUtg
4pIuqICg5E7QEMvWV9/eja5EvmM6PEghzZHoCqkucjfeFQhjl6xlbLbjtQfADC7sgs8d+SzIoeSu
JpXO2gJwcjkpd8JollEdZufgOF7HETYPTTOxU7GK8fKd6iLMYeA3y1EjoTjVnxRxfKEiyh7P5iKx
mqbkGlRibXXBvXloniIEWFxuW9XCtRw1n8KNAGK/2WDqHIMMAphVVSZ21S1YR4fh3GT/NxPrg4pC
cY3subLQytBdEuR/IvOJZAw59GvHUW7gqLQeDSTrDzThbVhj1V78cq942XjucYQFhYIWmUMeWN4h
C4nSs/cj0ucYOFiI8GUlKeKA9bACXmWK7FTw7F0QCM7bgPd7DeuHdv8YeqW1oDHJ8d6J3fJetMgt
Bamv5e7KMbQU0IbH2QyUwdUKsIvzmBefWLJFOTGgTaX1WKphvoQ5IWFlcH0ovRMLsbdRvyYVuH1B
06PSSkvOUXFJkp9JyGbHB25RLooUq9Qh2eTEV/hBLU1QebnNY9hKL8bG7KdXPdj5Hc28TECdScAA
/bh2zjEwXNQBU76sA/u0NIe3k14wYg3KlRVeZRWGgVo4SYZf0R8chyBbBL9RAHAnv4ezdOGvYWjs
c41G2dxvwp3S/T2a/V4O21f9buxNz20v0M3mucrEs5ja+oCwF06Uw0EvXaOxOYRzIIg8KAILeyLG
5J4RsiK/iqcPXB9pkGiu/o1azIFVUeLCb053mnvDziXwpLor6O0Z1ok7r3cdiKK2KNninH4d45lB
mW5dNz9j2zyY9kpIiVYxbeUAL5HMQrhSFJWs4PQnwD8TC+zdHr9iWHK8JzAmIVwqlhWrpQoeiwnn
3FQYq9Wi9TdJSeIYY4r4JLv4Qj0LYrg76szxBYI5aV0UI+yYFdyP5DRdmfJn9c3DEWqCc4kxF0r4
mg2P2BdkKnSJnwtS0nVErvkkqVy9O9gXKWL5cP9XNql9FZOmauDfeIc6SoAGYfC6tfd/onr4MFmw
pjn7WtMna7ZOJkviPA7G69P+uP+y7Xas/eJ6ziJOXDZp3GosoU7XKhBGEcCoEspWFdhDs3MMXdYa
APh5qFtJtMVddJJhgOHd/neJD0XOS27G+0QAsdUep51r5OaRL1uIhM3U4CC5e+6Y+gU2evlKR0eK
L4AUJ1TDNUSvlDO8tZUh2on/YUX7kMk+F+scErjWe39Hh18rZqMUG/P1Qkwis0Z1F4r6qXjKbFe1
62yxYMi2f8meU70+JnPQAQtZT6df8hjggHhFhurzEMn/iPD4GMYNGeOmgzV6irVXFbgP3KS6oa1K
rJVpf1d8M/sEpDJud5LlCgebhsqEPKLhHu3C6DvotPJB34+nHHtSpVwXT2TzbA5FLIcvzHxm6xg1
3sdGQ9aBSr6w9lxwrH+ooDlSOEP9FYCZ70GfbcQL5cCd5M/nll+6HylilYHp5tnbFDgEj23uDREG
rHTAGqnMB7LwIhS1SaBScP2TrMlDKS67nGDHzBq+ldrobdsZ1CmmRHJ3G0DZW+nz4jZvdA0jUpMH
/hBNyIpqDkUcnvEM3jkjon3wMOGseRnto3k8dacVSB5b7xtdpCIC9L70HDSkO6kBwWsfA01VzB+B
eKbDw0ejuCmk7I4XDrYwyj7xbuZ7mrWW1IaedJyUSlg5Jwt0GxuyTWz2SVswv37YnDZc2p3EORb3
I3bzKljZIgh8PI+RsY2KjCM5kGMKnnGVeWvr9kPoXLwvJkdzWAR/Rn9GSuivko/njnKWkMJWlKPX
ahPFqnNY5uLibRfE7xFSjF7j564P7Pr4Zp6BWbk4RCqk5IMF2ZR0ny41AjjqiWXfO0i0JV7y+H+/
/8Nm43fo+wYffL9KGHpjjF1Ph7TRMSIBoYhajAT6jVRZQg814KZewZCu9ssRk4QKiFYFpcy4Ldh/
bnniV7qXOFpws7qX0lygcBo4hzoz6+tOITpVepIIXtojXsdvTyxg44/RQr09GA6NM+ObfHoCbXWK
Ubc1RaFLyTdkmuxE9jvWJQocMMNx/rexy6CC3zRWz1tWZzLmNMk3N8vDvTHQkY055DkjgQETHSiY
SLnTLKk26+R2UyhYWJSJElKf6YJR32Di6Bbng/iJftbF6+WihWLpFbpxhnbgdZgY4j/C7RBBE1ib
1H1f+1BLWSUzbBk5DUBn1ImJQs38gmNixqDMOBRs8qHSHBUp4lFIyQ9fA4rVBU+QWpfVdsCKcZdT
A68TMmO790TH8Ev9IFZP2J2bGNPJoZDlBJvd9TyWbKWLt+/3forne20uTValDP7itco11aw535vS
TU+8SL3yImYBz4C7LmaQzpWhLJn2LF52jCGmRfczUviMC91gkRd2/J0lr44W46eyBdcHOIjQWV6m
yqZpFoFUuof34hM9r6Ym3ZtzUc/lkqnh2WEdzSF5c34IEpi6VhGW5ShqwpzRf94zSUQtiJxhZuVL
jCRdRqdQD2exWk1Hh3lmn1FCp5GX/3fOMm422g+fvu6YIFN04tsZTy1EmuWopXgeaVbWg7R/Tbgq
wkrdyl9lzIxJBn+61m9elD6Mp+Yi4g4dYzWPYH5x/IXzs65LLIDWTUC7DfYM+k+xo0ZFyAn+yuIY
G/Q1C9RNiWVvOoSWioEpRCY20kvO0IVFZ3iz6JjCgLvEnG9D3k7M8vV8Fou7YDeFx9x/eoY4vJeg
D2tWp6rpIGg0QABdLQAzfvOrZhh8v010EByzjOTaiSlgalgdCoiAoKrUJ0hosnN9T0vXTEJotnFg
chTPlLXKkW74zM5CweVS2VR+3aJne4Qz+7AxWGztr1+rdPKGI+iOiFEvwJOgZ52SdGcwMY+GN2+1
fUIkimAqEBSJeavhSCrQr6Qc2TBzQb3jEzf2MzgZMSx9DiM3bjldvExW3d/6jASprxHPEoTZbmio
Uc4TRzH4M9AX+8s66xeZ6XS9w+AwdQUFB7Gmu8rEv5Zf0IvzpsRWlBv+QIejBDMaOrsFLSqTXA0u
qJhoxmK63NDzC9H182jzUn+qyUx3UU/GdpxZEE/i/x8a/FB4ZcKdEjvCPXbEFzDChFBnWSzn+UqW
snmcIsFYckdULN5xjk3E+zpRKyOUYzEpoc5iiu/evtLaePcezIOVhn9wy9uDOgM4dT7gKdT+W1ra
QU33d1u/95fPA543V9EFlLAGqYrHdycKVQ7lDK0VZxvcbqAoA1LTrAuryW9cSxCRQlIT37vX7Fuo
OyU7/kRG+1gApFe3KHbgovkzecmFx15LDDZIWr3sWjUYWzWi2BnTpCkJfpX8et3h70ae0DAzYOCn
WJBlu/FlvyUxlZdEQX1c3z4mmSInBEBFIguQOFN3h0HZFxokPws+al+VRna2bp1EbdYf2W+XpJ6y
jSmrBifRXp4tHyMHFgWs8N5NWtrr/Z4qe6E7NW5oGuQUj7o6wC0P1IEacOy6vjknAVTBL9djgOgQ
QHh+Je01wx4HobXFJGcmVzUkaBluk2HZzqjr2aKs4WXM3zSb1prqQ0Ybkz6JcerdSy4JTesnfQRr
Hf4xmahgvudYxdCB5HC4owTKSpKt2b6nCQSY4xR/bmicPNMjKbFmufVG2u2iJgqUVrHrx7koR1F3
x8IOxI2SLSUmlyPy2txhNJitw59xyLvcVb3U1MBXOPK+YLdCAPLNQqM88JlX1T+EqnUq+f4vf+2+
heagtTWicCJdRdd/k3xu9uP9zcWLalUMD3kf2Tw6Vqy3d9PUZ8Q8JnuBhDlQr9O0NIxO1xW3sGC0
9GTUAW9TkpgBelWr+jvgXrjlz0b9lw3VKvpwt5czKpQ8ced0F4nE7sLlwzI4YuIs1WgXOsQ4gRLT
hUVgiyVHNZrv8rz+7NfPnuDYyyATu7HeOFZbYJMb4qcQ/xDm1/FW0gn8gl3dBZwbZY+tmsPzmu+u
ruJzNYncYX5xPM1iNfr6Xcp6OqXrIvF4OQvTL8cbnxvftT7ujOq4z6rTcaoOnbJNmbZ0937KWamC
n7IpmmT8fIacciud9M6GQt+ShrUKBjm8kyew9DOkbSmBuElQYEK0Et03uU8BuMokKLKdl2N6r+P6
Vv3cAakBFdjqiPpnla+Cph4VRwyxBxOB+Ke6nuVCVQJ14FSRiyLNSk0aXAaUudR+HYeJn2w7SjZ4
FQOO0OwZzdZPphcWb2zZl7q0hZusuwz5px3f/KqJ1mKi7PR5/fAFfCYAH/hs/3p/kVEsJaPmyGWR
XaPC61siV1fHMeXu6NTZRHjLpRSMgqsRBw8GL4fQ+kCRx3A8Pb9jLiaozis/vkwZ7CBAuRTrEClx
h0/1ZMd8ie8Fo9tuyjt8Eya9C9kGnVNibWjMNuDAcQc7OEI49LY95xk437yrRvWFlJH+cYaZUujd
F+6LVQcaNcyV3JPVNv0cx7aZnEhrEmkZpVgCTNzd9i8HumLPFqMlihd1wA5/WkOSpZkFtZcAaVE6
4y2GMwlZOrcYoMZxxWWWK/EyJBpcobL7+Exak1cuKyEP/A5tMSH/CGlHewgC8qSX2HAI/jzv1gcb
mwpq9iRfgwFeppNIzkXvilJirzIWIWt1lxpbuOQRS1KtzSYjBoJUWRmzNEDUF42BNxZZqZ8C4ozT
VHm7xjTyHi1jpipWRS25fdG+mbsm7LDNtK4uXYDrQQEUHmp/ET0bQkaUxcrsou7nVr8RXXFWFxEi
R3/pSgkDjK1gGedAR//TbCUNcCKMQGd3rpPoIPEJWZyTSixv8R3U4lMgRPeTB+wvd+6RiX9m/1cM
pPHJszvFsMS9cW3ROPpfKwcqhcqWxruKcThWjQF5nSP2xGQcJWEAY+xle0IIgEH4g42zz74N4kfr
zuJXBk8/+bJ25SA5xM1XKPtp+/12S7Ei8/prrshm4R2cdlX9Fic36ygRBzZThVaaTxpad2bUaUqS
cxFdHQYtr/X2lOv8/IhJkomrJmfOqnGET+H0xAUga2qaEqDHveYozu3l1CI4W3Woa9kfXjL62t8H
o4ztdgp4/M+UksFqxeM9hzm83DBk3AEdr5MCGedCiHt6sELyDiv5rF0+bV0HC+0XQy6QB044tn3C
boUX3ntkCWflN7CnEV6HGNEY/L2IRSMH8oWmYr8z/yiVDcm4BN0ZJB4Wj2Ruxs1zZU4Aw4Aly71v
FowFHxgFJSg+VVqiSo5ZJDM5HknY2Bx7H2YZCVpIJoUwMUhpHx0cYDzd440SwucUD27wnR1G5ShK
vgy1TgoQbGDAY3IZ3Xrhnzppq1EZ0k7cyarnFECgsIyupLmM+Ev4KvddOwYwwM8G0ArtElLpZ5/R
LrmD48pyMgHwSsHpgphQXpx12uLidYSAdDeYxKIqeFbU1bFcIHbyLX+van88L1v0zfDhwHpYsxoI
x0TeMJ4rU18cK7nfmETav59gt7+t0jcwbg40Cyvl1hsGkPLtrSI3hBytVJAGmPzFYgCVet+Fwt4o
uIcfevdSOYztSC0H441n95FhlD2XRbyJX2DaVr5y0ol4VLkMwQzesqw9P4LEa8m3kZZ74l3a2Lr7
7Ds1n7O9KzqNxq6xzRrFIDppZB6hVzbJoC3ClYE+WiXJtd1YprWwPquycmLfS0+/zygnAElqQg3n
B5cyF5CJ2lmscs3N4F1fr+PpjtGrica1mAqMlVgP15VnqciqoQopBnCWwjzJxd0EABB6yn0p/Px9
GwVcqDru0lEOZcds08OFVM/3PeoBElfkEumfs9PUBEhGQhXgzqDkLjMdvTtQTGiTV3SQcvEZse5T
fBu4pLN8G0T0+pDy0p4uwdwQuLh7jGsKohPopB7/l4iJUre8hKWiYsQHCw1EejWmP+5YIv68jUbB
8U3Xa4tjHjWYXsGYih9SkiOpOyK/UOT3OJI4iCDwnKvCBh1URYAVWef627+2ndIVOJOdOQ+p9MrY
yJj9Omqj4BKXZMLO5zXh8YYoo6x9wOYiT8K6VQtRG0PGEIShqP5y+KnFDU6Wb5OOwIQJMyMYZjsb
kJBqQluJxtjwJl5EUPLotAtiAw6iHUFNwRlXpZpkHIsGJhPWTS7cJw0eIbak6pHv/IcCb+clQAJy
VfzYe5veefRsAKP52KvPVPvOkapUMLOfdAygAiuPReAvKvDaamKO/cW+Eksrp3hAaGQ7nmuuk+6a
7VqJz4jZdlo4Pm9xRwMCarquNQZvXmtRwvJTw08FFSCrA/Cvv4bqZvVOkKMostIoI91fQW1foQ7M
eJJGt9u7sX23GF01YFD9xGA7l+T/Nd/fBrILNxicgx95CUC+rNOO3Ou88oFU7tKrXS14dl8Mq48X
SstZezv4hZH8apHs7uHff7VxemqYfMqjtiFs2FPXD5X+Wu5TLaQ1ZGhGRlA9YJv9NuD9N6I6Z4j0
fPz4x1TTcab2C4PxoUxtFe0sponGV27RqQ5V0FatRfuZCv31nKLlI2vvfod4g2nMGaXxSXclzrOx
OsDhc5FLRTPL+Tsqlap1ZlN78EaXUhMu27E6vraQbUEhSvGgsh5yMAER7kGifMxEXsX9Gj9JAuno
enzo7irYxeYLALQaNe8ZsIQcKAmEBi7D7CoR1Mj6pd1WhyVQVK2JGrhWglslpHqt09Oq7ni1KKF8
SMCYbV+8/8xoAeaFg3JNgMtWXuMuj694onpr9yXl9+8Ivx2wnlKaFt7WayZe3rv9oRIeVHhlSt/i
0akneFx9+VV3ggpVMrGrWSTa2INTbsM7Pm7+LQlTuwuV7cJOwdT0W1Me8QE9I5qJV05hfxfMt+d2
1Q/HsdzBbMGymUxYbds43UF1euWdSJ5LTyXZSf+BIT7B4/LxBdii7whZQ6RqECxMbmXqG6h5rLm+
yTYuM0enrxZVJXOnprGe0+hTk9wiXH9OmWHB1175CvUp0IVnEzMTZQUe4SBCOqxAc+7464C6K91V
k06H8foZ8CjhiF8m260SzK3DITI09mo77f7Qo6zbv9USfeZE4SkCCjMS4/uXWFyVNYIkpxDyhgFJ
kUVjuoSz0SnNrJ41er9xCyApT4QrNTrN+by6eU+bvka5dntgs3TMkLnK6TGIP4uu83EHRDDt/5ro
WC+aMG/3WYn8/hwrXKYSSAsYQUSM7AomiQkSDQ5ODXrcMXE8n6nNCm9W1xpCN3ROHqvtby2O3VKf
qITER7Ddti6pKRE2P78N5vwRP0lBk2SMTrmfZNEf/Mzhqwo6YJJYCCnigXnL3FuZ3EtAK2Wd99pG
pbmZRtztZtTnL43TbjXUxFUnTV1cHVLxzVWuOF2m2PfVNx5iP0I+SqmhZYf2oYXmMt74DS+GOq9h
/wpiarj72A/BLlG3+pGOUWCRyOBA/Ar1vG/dH7frYWjmJY9Z3k87TMkUqKVP+n1F0Mm8KM8Y6CWN
5Vx4tVTvgv00HXMLh6BUGUvyftQiPJGFDWSLit9hpw/Trwk0gYpnshvniJPR9xa3c3FJWQ9LbFqI
4zuoQnss8LDS8YoOQA9Qq64+lOUN3LwSpJc2zUFROjsCmEI1x6kxPz1G3GhvnkTLVe8XI1CtsCXS
Bjn15Htqwm+J4prmrxmbXlDqpeeA8kennxKcPZaxf71ugZY9hPeF2SrzZiN1A0iSrHE6uKQVItcf
JoVSQ9ItFlChl5y98YTlqSXtcvDEUw42mJ9byi6Nf453jCXExKvCRMQALDZ5rTvJdD/YJtFSE/C+
V4XogADk2qS3o5vQ+9UdsVGDHNgcXdohvXkqwzP25MLwaPGaMUhOmwr7+uPNzqprRCrXIz/RwaPJ
bVCbI+fSdwPnfDJDOVayYFHAqnBaxm04N5Kdi2OcdcIwvnFa7WCPTf9IZBbfA32/NIOFTaAHIHmk
/WdUNUYwK8k73olFp8mY8FN8zGi+okRiCFmHLXChBnOQnAWbEeC0gSRxlI+YCrNSapfwex5rqtwl
IS413Zc+jMnoa6dy+GGARei6fLyjdAZqxGjac6ETbvIj7OdsTh2rRlmb4CJj/8A6OxwAUcWRS7eD
w1vEBJtr0HQu/V8QI7P4nJB0aB9xwF+sVEjEsY7Z0Xq6ll7el98UVRw3Qrk3nI6SuW3a1huFyHKr
eHREJYP/v8rq+Sn4uK8Y0f9KNaHXCeK+rd9MRtTXfVRPxqRqjQePvjYgUN5jpz2hDst8nxSBpNGu
94oYrlirjLr5CCc+gn3CzwYwvzgEPBzH5Z8Qnm+uv23tfhFCkOX7/TQWiMBMlxj44yoQI2hLjVLJ
qgXtiUrFOealsWWnPwDT4wzqOt9dCUqNEuEwHge+5Uc6J7lAkmJne6ZXouKdt0rgVHPrQ4XSJE66
TnuftWWvYYcT1CuP5Wu94/Q/IPQWuKEaYVCQwoMaOfxJBUKtVNIIzxteXCh2J7PI1gsOPLdhyeEj
z8O6vKZiZVqeb3qx14NOiuWmNJg7xcLIWLxe2U1WQYiYI3FXSLuAmorBnHExmjjnxS/vihqa2a1M
METD3Z/1PLclrGDPRdX/ege6GGivaAf2RZ+BUxMnu0jDH/O8fOdkK705cnavX2nc/7KvZZSTzJQV
pM0dqoOtdRQflxBY8bBV2QzZtzlvDJK6iRBJo6g9l3kxv9hZv5UAgeeOibpGyoYGjTJHbb5F+q5i
V1SNKTpJYpfgeLG0C2J29a4cXz4oPj2eKCfYbOoGK/QpouiXk290fKiOfKzucHhGSKkauDWR82xw
zysvglOkg12gRtge1m8n63qmynV/jf5UcrKumM/KLDrjbSB22b8/QYSmgiPSwLlgvHofHRmpYJW1
5uNulwphsx7Ya2KyEbcKvVpW88W/riTNLXcShKB3NsFSxNPiWQBS9fkSRxEyNm8MnYxS+c0PwuLa
9e94Qbvs51G5g5kXOm7yEjk28hp+D8nJBvCIb9cQ1FAILumjAdgSAfykjzYuMFQQpyCYiLbap8Ja
XNpENY0mEY4pPus3k6pCiVpH2U6aTON74B/obf+z7qJOGyiS5Xjeq6gjrwIKBgoc6rSLmBYiy2Rx
xmJiH6J4kf5SjPsC8LuNnhy+9jOWYrnu2TMcfxizIaCof0E3dEU3TH6e1wEnyPYrPj5HeY3t20XF
3pnzlHlYDw3P1Ofejnzo6MD98B4aoLbqnDzUDnAmqqYqbKVRnXRRiAY5ljAQhRDRRAuiDu8JNN4I
ctn6GKy8BHafEMIurytYz0igiE94nJdKZYTo277IMZvWivOR1qLZnW4kE8eIM1ioK9ypYfax9rTK
etPja1vgb8Ayp5HD6hU2TTbT8AHnlqsLjrkcb5S1jJUNdhAT32QNkqI8LXA+qO3O6P5QBh8Km5Gd
ASfqx4Ple5Ck6jJFWdFCeyS5br1hR/qaNCJo36aY9/XDAgqqsrvS+9KU9j0wpGMmgLskBY7VjXt3
ZmHRebadKLY+/6w9nBN/IgvP355qDgG7YiAyGh/A/CCqRMsNP3NV9cnKHrXscxmPqQiX62SYt31f
MLfZCx6uaNJtEIq3zTiZZ+ewMKka+kyRstM2GYtQW945AiQ3nTLagiaFsCSSSobzdPTTwHUyzhaX
W/Y9AWLqKzclBW4nzXzLnEwj4NyPscAF+ZRUt6B8qbDpkXpQSf1KSOzpm3VbNuLVTay1A5WzrSRY
FGsT2eXblbhzOqsET45mn1rJ5jx+kIaLytHb1dsBBKmxfJYFnRdpOj4ZuJNN4HyceMQUeJaahTAz
uFdrTmg0JMnWN58xJTLgphZ0xBIlPCpG5Y11T9xu/1BVm/wwWySyXcDpaKDuuG1bvu13DUzTl2Gm
/5m9D2WcZp32drqlGmb7Knvp2zKhAZBulPMxf0HXu31EtbSXotJ8dlZdYOqro7wbr4HKiYgmK090
c52utNggOT6JLCdcY2u8ScfNYkzgRBPpmJjzt0ZdZmBOIe1iCsLK/AZy/MVBw672rmwcNDoyUXon
79XaUlcgTQ/jlum0R6CCuOrXmN58icYctgO8Xzymp5iYMb98EYfQlDKdzWtkbT//zQ+jIdpotX83
EajXueyLatsgivLaCfqu3KHMLcdnTVAI5npHKbiKe1xmAwYZpmAplur5VsmOUs3nUZfcbCq1QJ+c
xVMbpXprKTm/6Xgi1h3Gnle6+sA8wAvgMw7rGrkUA8E3R6yGxpBM13UttTcOVzHrL/xAaJLU3QNm
i2x/4mUH72uqI7ScNHpJIjNEtH/a2cURDBWermQHK3u9yqTDQDzWuSMOuogh54jnZvlAGqcT3qXu
n5r8UIvS5XvpI/Y54Ag/WjQUTvdpx5qQ2UZ3Ec2F8+Rmen5J/MGwoEaSke6mEF3XPTgwCEr1veLz
Wb0C7pVQbilu05u1Ogc4NUnIKHyShZee49Un4XfndDFkDWBLpm3vWtGUpQNvgX/T+WAGvubG+fcM
sIBhRnK+5eyChu7/VfKMKYWPAuQGGabycI+g0YkkR6Mo/yIOwnQUUbiZuo9BvdiXTC1qLJsbhkj9
uF0a8CCgHewGTl3Mkgakm2/rSNJVv5TW/OGUEdCuzdytDq+JNlxyojqD1we4mJ5gld6768m4+qZo
b2SkHYfGl4ZXIBkelMjHAuDmtPRUhqF0n0/nm8ftwgzpiwlcru8LD62a6cKQ9zAOWE9qfEBNZKe3
S+8EHe2rDGy5yNYDfD8xLykWF46YIDW/19zNotUUY1MEgar7+S960AKOKfLAuuQ4pGtIoN4KucUg
ueO5w8153TEBUc8c4QMufJGIe6geQYdpmX+zLHnFJqMjDL8WRjgzB5a2O49rU954iEDiy1bIZK8y
1CObOSGyq4L/iayr50l0e/fBsLnECv1PxtgH5mM5aNFaivk52mlFtyPQFpGfAAJ7oGe01NHI77fH
bHwhAKdESnKV0RBeJ5uZrcGVrCWhps01iznPyflKyc8gZrBSfD3NZkc0+CPCD5d/qqkSgRS0pKef
pL5c4RtaPIINAwb9hLt0XtAJ12Xg+b2eNzA50gxDG9nRkYrISxzVlnG63uQalaVgBwehlMZDSPWH
PuF2IuhareKKODAZiwoOO3fT7EddgGBuBcDSAcS4PMVrrUulBEahoFvhk9NEtdyu4qmbdOuskzYm
EDKT9i9Kwz1skaSdpID8+qIRz+MWwj93NiF/QZpIjJiYaHE6ULM9q/9JpsGIWvdz04Glme/0808E
MVRojqOZXUY0UBnavtnRwBpt0Nn1X90uPKQKq9RfeeDZNbIyPg+ZDOLYfiVH/Zx9MrqUVJj4WVkW
LMRGL5192jDeBl8Kg1/dVqo4keFPaXN+NFBd3hmm3rcj8fXUzCC7Dgv8VK0pTREy6bvhpVdv2wZS
bqEXL5hXpplDRHuZY1cf5+rgSKiO0xWgYpZXwFtKih+YD/QKXRGHoSj1qXtWH4mtketkZ/a1H6wJ
kzzFTEeXPBk4fJIT+NBPjXJtS3l2uByoH5G/IjM7AAABa2ZKqpLd44PTcCft6/8hvCBn+mgpbV5I
h39otqnaD4JG+ZpE3woCFQp0JIeiGHJOKvs4F4qT4tslavXaJ6fVEWSvTsugMqtfxeXCXJTC8qNJ
m5CQCicN08T0Sevjpt1XAhagL+f7u+paIkpAuXRUrnL1RTAT0aiLShHULDWglwtZiaswtnzALxvQ
k9ZK95RuytwT461HrsI70lSpqFopvgqlKid476ZM1e9yXbMqqoTyba4cFUrWCBRFzDyX7YIkDUZI
Zj6ix89OeH0hPt13vEc/9bzy4CTNqc0qbuTxFAitiCmB6AS0EpnjVsQKwnY8fK11QWm8OMJ59bLR
SIlr0SbTE69VXv382EmW0se+Ghno7iIrqbUKKQA6E4wvKQWZbcneWg+a1V5CFsF16ML31IR2vT/9
IOWcCe9pHQkindWCm3EZICRiXegdpOcCMN7RYJYBNca7Fpv6D0iKUHTItIG/ouw5lB6uGvIfSaFp
ORo0B32/p95pDrm/Ls09r/th/FVkLoNYpKRwyFvq7DL/6JMFMvm8LYIhMgIpibccc7smV+GSeySM
HgMLiwnWyre8HIQJD0bKfmhU0MXr00QM1iJHFHHAXMpHVBmtg8d+7oZk5FOFIpNWyzol903QBdUn
+rbFSouTX0baSnyvjg6E8iYp1DE6KHeITeFKfqvcZb0LpIift/CyyXFo1PW20xYiER4aigbOgzPD
32Txje9meNa8Vq0iQ4zdExRC0Mz4+Y2PRzr4kQivBhq8lMjNjJvNarYuTdBc6ormtTlL8oGLQZf3
7AEVsHFor0oqq5nCye1M1HdY3I+zQCXgNcgfWOso7k0sTpaUmxgX5sVyCbHmggcd7m0/zxAcG4A/
iLJexuAoz6lAGEllF3DS/qRC5NV4ubWJV7xm47yGtlhcK+gb+jBrYSoC6sm7dv6pns/Hpur53k+D
W527+kqHrtCq0wzBU/Ic47EDz1CcBIdZ5Qk+xhihAyI6Rqc9dY5WpaZKvXI0bHFcn1dV7CL14qD+
5yBlH22epe1qCwRcd2U3ed79kWKJPxmK5i/8aau0QdPggJ4ftiWb0H7ox3wh7l9poJCGj45OTC5j
1HdUyhV3yKPU/NXEgJM0fyi9cgSBzC+fabvVgJ9HlXMwMLM1VKT7dd7Ce/CQLMw4adkNPgVflVwi
LNYLR+NTxGlPInITIDcMf1FU5p2ZDiPH6jDuGtSZTa01Id+lxmZUSzdN89xu3fa9c0E/nWFHDFQU
rVa0f8/RiZep/xxFyr0JmLqqa0NJ980fhtWOMg/uCu4L5Wu81uvUKDYGtNhKJ+JKCxjUFSfzRgwt
2HLcJOd/hWwTiWzOYNA16S5vgbuo2noM7vqt4QNkC5PdbtNVbI/+hQLcsd5JKFK/u2MfrYn78O2a
2kJ2y2m/YdxtYz39iyUV3nqaf4S2n+Vlz2+mjQPMJuThTcEZd4AqG7bWLidvWoQsxH4t9kH0iuxf
SGvdfvfcTrEmiSyd5U2Wd+3sAHM4TfL/CaIU+n0oCFuJQoB0XT6yLF/dDAQAvgzWd6ibcdTbFgKL
IdjD2xWinI0gieO3EcUx+IfJbbSji6yrR1wgMCsYCGPZe5LMFGG/XgtGbELCpThpm0M+909xcE75
WkG+4l3mlRhLa7ofBwmWdFmRyEzYISppL8MDLL09KCYf7zsGW6q8sxN3b7K3tAGtQ0ytq89Bh94Y
kxVfcW/xUp05uc35ZvN+LLicao0mdFOaiskdoY/y30KV8gi6yqU27v7OaZlRARUbPWTrwN4D+2Pr
cvUPHWW8V4WrpNmTsPNvUZRmMvcTcWMmLuNcv+Qka7VSIkBgFzt1n/V003LYC4S/WJRHMx7oBWNq
KjJSNGi7B9ArtfjafIlzKtVG46WRR/OfVy1TO3tUnbOazsUSA6lxRC9eDWYeB9NRilf09R6V/1Rm
UPcl2ghaqhhyn4YURcNJOUlE7d236fWy8Nk0Yi0zvEerH6AmegNOj1tDAEcjxnK//aSniJ7CuQpI
FJ8Z5ebzAsCzlpj6v6BiGxjMoWfxfDqImiR9+UbqiTW5l5i67spJiV3XBrtL+gnrvs02b+zVevX7
owPl0/TJqv/gix1n8Fw7wtLlZMuZkcYH/5Q/rOilRTJ4mjtD7vGSna0E0Npm6SZ29cPuT3w7NVzn
Dl94AzleORcCosycBiZtuHnTHkVqpQK2eBbiSfIGXXAVHjXBzRbxouI9GmvgDRkl8CllYUw1ZrGc
jsCqTsGw+wkmG0GrAuUmMDVHoGzP/ERd0Jpwx7g2/ktqMFRHsiqNL/Su/pJDVdX/ZPhKsTa5YoSn
kNo3WAnDQbgrRo+6x5RUv/ybncfUd2UoMxb7BKXrUx20CJPxCGCmLjI0G0hNnN/guBKbCkMBhYdq
hMe6xRi3vaOHYxSdARt+IDlfP3DoikUYn9lZIGLyqorcVv0n4AH0fOQuQRt7gyUF7Eh+d2XOy4iA
Q/XmLBE7nlc/Sp/Gy/bEWCI2ob9M16QNESDbyVz29/e1nh0h2vejs7Yxym8j3u9KPDS+96rAYGOe
8gNqQ32xjoplSZWC02z6ssIpycVdPlAg/S0Bn1cLblyfGKO/Csp86VnvnCMYpRFfFuxFLu6NWNIe
3x3LdbwqUhhAsNwEIvg55hOAxhp9N++dQc3k5BzGom/mN8HmT26UJz2g0J2Xho4C0vaPJbvwsc5t
D0SAJ0XA3tBor31cGBz3UplrKM+ZEfDhGS1TulgTj+Upuo3QmOXkUnxwq82xyJ4WOo9piAxt6IYw
zq9re9O4rnzObVtjIHCNSfUXv4hW/O8azk3KVzGI1eewTwMUdW5Nt7c6egEnyCBKgYhZJk0JJDxQ
E0Hq5RQh9Fu6qE47FnP4wBbqee6JMp9o1gvUHoQDnm9mxjLVrZEPH3xDuCpOSaJtbTI8axS0JzDJ
bHpAJuf3soz15yz0d2ji5yAKckxbt38ruV1KzpkFy5mNPaMd9ip9QghJnbWV4vYB57vbScIL5pRl
CVX4AyknIAQUlsM+rRUj5vbN43TO8fIY6/EFc7WjFXORZB9yCg8AMX6+jkQuzrVK8g1h8jLpj6o+
yjfi34d31uznJiH4njvLh4M8JmYv2xIcpaxo/llJYFz9tJmMbDPOaj0hsYfMTgLejPPEuwodoX2c
bb2hv6uvGT12Ikj5TuCMdOodkRaHqY3o9WCbwDfiE4IUuCZeqN7mnA59t0uhnGCATaSmVbTf2ObL
qllr6cVESc6QTia5Hrg0X8d4tsax+UkoNRwAiKApgk8mzF4+boTlWVSoxtiz0Oc06M4ooJzcEl5s
L2ZhI56LL02mtd2L84UOkoseMrmVBZSsNvxaLMzQvRXakPmt3ObO9+0Y/6cZGhhnt1taAfvNc31L
k2GoRfPGwN7zYOHnTuEt0+hW1DuXFOAdcqHqpyRWgpyysoCkQwQr6Gsq+Hj2iyhsN4zCLkTyfn6d
D65fShv+lxbcD3tIdfqOJZB1j0COKeClA2G+0htGbkZTwt81aq9eE2nZdr8FeCc7oToV2R5C2ynw
5+hQWZ/El8VWqJuETa4zD4439rGZuntxVLsEuiQZU/lJcOgDAbvhiwjG87/k/NptP6K/xQseTxCG
+SLi6slEx+bsabwebSqb+NvyZq+yBgjdGznetqDQCnlFfAlAesZ+l5zfGapGl9gqiM6iu7dBfCzP
ppPqyDjbKKANocPyuQrAQoJHSHXF8NndZz18CZigvjp7uoBzRdt/mDMZ6ioIbTC05vkJE3ChsPAA
cc8RVDZVz71XRIkV1iFqJwM3aZYs7mwe0K+KoNwSsBg3PrVzz7Z5jaudIXync1G4HQAnKcm5jJgY
e2jhCzTWXSTmGja9qYHV07H6vTfbITTVNfECaHMO5honSZ/cPXzYt7eRhcymJiMTbXEhoeIysDuc
FvIyGKLc5kmVDX2kCSEfK8YY3H5lZzU+uFNeJpP7grOUItlKtq7OcAFATZ4nIl7rRm7DngCcZUJO
lfh7rAEIMxLMXyemC9ZJI/OIVtOnfGg1cx9vZtg/7yqGWDvRST91ZpLdHE02xTdcDoZNk5mauFHr
xOGxpx2SQltQqcOizrRZRpkYh38t8KAuVQyfnpaIGvdtk6kjgVy2QyPSg4vtDjXkwflZChq9ZUNs
FLVlOcYpqo/HXuV9fJ7i2DVcpFEn6zPUNwM38M02W6gYNFlPQ5EoPU3/AhLG4E0qF/L2kzi45231
ae4AbVnUZVbNy5mtnNQsvkNBEr6DqjhWTeayjyOJzfMHtbxpvESLZ2RYSsh7Fu5jfSmEoCN/BVIz
ClkU1HL7m0svhTokU1ML8Xxs/F80wpGxwBfVuL+9VvOZdPBxn5CWfu34gN+iHXGZnzxX6xGaquGE
s2mnBQULBXfAE11bX0T8vXwLkqqyfCsztQd4YzCFBliEduIiJmeFtNJ0mpkPZhCQu9caVpvoD2+4
e0yujWtvWL+rsmYpd9GNVvSscMczlUBh4dZcEoS9vzzo9Ts92RJrMp10lkB9b1WK3Y33cFIwjNpS
OoJq6dRvVcfoVgpRCp7mZk0n6RO2lL7jR1yCGcHemSX4rgzp4R8OIUT5maevHNWLK0K068E3DrtM
CzH1OBc2Mm+54+cVcTkIDlyKLppNlt5aba1H8K07AsypwZZyhLzmjnf23B7F3gIu0HIbr/0NaYnr
wIfo30d0Jja4ZZ9hmV0q3xRFXZzVF/JzB96/d/tjrTmFVYLj5SbmDSsuSbMsAh0CZqy0v8R1YnMx
j2s4GKEmfdY0hlOQSx+e6HrPFKiG/KnpcbNUW0OsneNMRRX6L45AzN/+FjDNRRRK2L1tmRfMBmcA
2tkM0DPDVR7goZIpUOpEq6jl8lstQt537M5SYpMCpIGOAFgDbQmXyg0cdPrZAbW06uYSa9OztwHm
m7Lfig7caZZq2BbR0q3UijYhxvm56aGv1JBbWhdFGmRTNr/re9azBe1XIU6Cib4iFASgFWdp8/0M
2sricYx8cfHx36xheyVX1P9r+zoDEz9ig2u3pGQL3q1ZhdAL3Kxmh8lLLdymccisN+QAw/DJr+YM
qY1P+1vAJSvm4UdhB9eL11hbCs2xSQP2rk+98U2Z+RiRtHmZ/WkELBhxaj3Eqhoqqu1bfYfzIWNC
bcj+v50O3Bumc2mouu0UJM7iZibXlhIq90WSdD2mRotOzJ4y+xwzTfE459r0OhyCoU6WosxAJONx
IkqbtWrefFQUC9OdbwyunrikBGsEmv88QXp9EEhH3GMWVWyvam2d6atAFu2OvvXOGEhzw2iqUb1t
BypvZccz3NLwIuwodrHHtxhLkq1WvX9eHlOsLXBO/xyk3DURMMcJ9XJ9ilAXzcOAxaeVTzdDAHlG
A3kmDxGiwC/sNJXQOfpNVcQYJWPAUL2ZIAEtQAx8LyNxcESEnLqSuyq0KjZ28I/lhA4KEwX1JwJE
6QEleoFKEpaxryMkMT77ToWbxl9Fgj6hoDiqCgHK8upAsqjeHdxfwY7GJbx20bFUUlF/nOPkY7SS
W0p/kt9z4fzMNLp+o9B0ssDILjAybrDKH50DWouO2WRK7Rb0db9cG4j4nukF/uXZ6YLBHdVlrO+h
RxL2fIJ9lyFnZUcnbgguiszhDH4wy6TX7APtRZTq5MPPZT580jQY3xgVXXeifEmXs+f3mqufqoSB
yYf4hgFSSF+ltvPiZNIHdmnDTaMVliQ+ps6kfeogS60u4Arha4thajUyvRS5SEEMtwbrLyj1bIRN
H/z+Gv1NgYxfHHL/d07oJ1NvxmTzrHa7uZ1rbwute7PPD81jASPK2UtqDWa70MY6QtWj7ah75pHN
Q4pnWXx07KlHKUGJLi1vZI8Q2muK6v42UPHEXW8ijMriZ8XLurSiBgM7yAjLDGVhvaFHm0aojn4T
AwpfxwIbHA/XjKE3CHJ54tFDLyKd7inY6HEEkcY7/+erkxspnUfzV8/dSykxCdH+CoCWfIuY9jHl
fgl+p1PO1Yg6Uk3o82TMpR3GavJ8jOarr1vY8fybXyKaZ51uHj8EYHkhxHidUTrb13uP+g4fJIEr
Up/Ci25TeelVCHfNdX+DbpWlHkpBqsVWKvfxWZgfHWWJa9FCqSxgVYK7m7XGLo8yRcqAH8IucFlR
7FbDQLzRMwtX5XGQkYaue4tAxO9bxFQgMuWo41q0dbDPHFv3zarlwuzdharRrkxWX2oDgtznednV
43E5LHO3uOOt7ZXEEMUKwb1XLuGQp27fjzYyltQUxA7B5QDaW+6fck3Z1U9Bp6LNnSQdOyv59m2J
UIwVdqHZqZy5pEAfyOToUa8FyRLe0KBsUqUZiXtN0Mv0ay3KFXrxGJWx3vI/jYJRdL7abETQzV5C
72CwWWSEmBZVz0TPHF+jDMNf0tv3D+e13Qr7844MaRvv6dgQGfi4MImD4i3/Y+nZwcxGIOg4pjTL
N3E0vJ0iir++LEdNim6knxSuBNxy+hb5eKX2J3dzwkqO9ybVJ8PFFMDI0oZGAsLWzUNfqDeJoK6C
Ey4C2On+0kYR33R6/YD7clzftG+pBj9P+ceh2wyvXOpRBUpiv5vCo3O2/N2vfqh3xNuskklCck0P
7reNFsUPxnIqITqA4mUi9Gojwl0Ez7pQGj72vJofJLc9+uGlObY/Ndq6THhGb3nWWvNcW3GkPg5f
ivU5w1EK5MxkRRyIvd0xmGnezGMjUNiTuOgjD8U9RbplsRXHCSeG5C2BzMQCb7o2SN6tLQngCAVq
OS0tfureMi5bf22zhE53ZPE/TN0mlutHUY1dNXLScMy3Z3Hf3CPoHgEaoxw7AlV/L701yz4w/IaA
E/WZAZYKsjCBF30Ceu75Z3S6hwfBS/ZcuqaAHZdiC0xje5eQbkJo0izvAwlQJT+MRKkL1/E2M5o/
PWEwg7kzqgliRkVCVqfoKZ7p0EnED7fKacPJIx/0m0PI6zVsJh1Jv1kMc1/1uD+9gTQTzyOd0e3o
JcukJJ+6kXJtEKqCvOPZpFE5enPQpo8tJIb0cWIF5N5oWlXo2WO/S+X9xiFHyiWvxF5UclOvX75m
6mmCi2Mq3VrID8HAsMPSn4rTbly3XLpQ5gn5Y8HTsWfnKtaibQ9g3VTrH+tIZq3lmIRiUJgcdahi
BU4s9woF3IVUuk3JbSyPDG4yA7Z8Fzm0thpo/MHs7qVPoDk7J23GiIvj/KaMqOI/0pMxFKP4nT4v
k+FuucwYR7idh6Oy0AaJvoo0dHhbLUSzigc0Lo+412Ux0pHOVKnXsKW0haUh4x/CDK0gsZSRzxQ9
4zoBX1fzuLDyGis1QvhnZPnVWWFkwcsTyIkbMlPtRoiHv03R102UFZYy7pSMZqUwjt7DFeTh+NCu
/20bjo6+LyKhY6HoQPZcnLScLKzJMlX3aFiJAnfuq7l/nllFPUagvei3yYtkXBLIp+E2HQOe44yc
68gWnMVynT4zOYCLrFZBJ0VPvQP1GvlSNC04wFy9P+VlzyGpcfIPstGpy0QKcaKzLwKi1XZxJsjm
0wDOtjP/+3wzz5/u9MDxjDRqDLqwWX4vrLAjpfw5DaEVJljMFvo74RRvDnH4vTFSnPlFg3d3fbh4
P0uWjlHISg+RHSJqA7mPX9QH1ShElyVW1mt3k4vVTMyD8KSOUgyb85/zxzyX/jOyfuLPhtNL7gfH
WWJkMQeAHvqHHm3IbqJcMpkX/SW05DBbKXo8ghkwNh13U6pQ0TXKsyEnITIw3sPbY2y+wvUIZWBP
AAsSxiyOVYiLyx4tDX0p7jYg/MfnunHhyCwbxzUrwMFZpXl/hpE/PI08JvqxyJ2aEwkBML0ELwqX
a3US+DDKZP9PAwb0nyOVZK+N6mB2PcO4ymwha58GK+PcBFBqhsCx7f5QZUZRA3B4BjnIDBpsWShR
DGf7X7hIa10Q+P+Pdqbo7kYUEe8oGxoankuh9ESZ+MG0EyPQszfTAbVHRjE5N2Hk2kih79JU4+4m
cPVFzUrn3G6fsOpugxZGrm8cSO1DiwPU8Wmqdtb6rgvpJroirPJEbQn4GRCshy0OnBDAIw1RlAhe
HeslaJ68kMXHl6PL0J3S4rsUA35p2JAn7OPlRKVx/OigjlvnF+o+xd0+3N8BhhfVvn0O19DO+gqW
VB3ugKeH0g1a5wPr5ApNpeASzFed1Th4VdcUNKWCwwDqkY4r/+TmYVsIargbcA+g1KjlimMAOrHu
luBllEY3YnA9KDM+G/0o6NlVJOq1+0PDoNU28k13ZPqcBY92jeJAVOk3PJunXzjh2EfJPjTkrBBD
xUd58Mh4mwAGxGq79U3QGgK3/BKqiPrwZc9BW7HrFHrY/qqHzr7iotsuLKrJuC78TK7bfIE9Nwio
6pAki3ceSd8OzPvXT/k1lg6/3hUxCiIApC1gLpPczVKfiTBAOB0vcl2el64BkEMb2IV3Bj6/xxgJ
6kJRxrSgAMll5w65Kg30QUHWqk/caR5UqMWlQtOH4ZhcFaMVle9dr5r9eVzR7oWOZDl96/Fou9Af
32Kd1ACjgs1YtiVXWyLdAHK7tAbhit8LScscjwmG7PDqJD2ifFl3wUidNuWLH9feuyGPBDRkJC5g
j+mY2ILxl+zFeA0KnZnpzY2BSaVKySg1n2vOniBSzlEh/f+o+6Q7BrblyALLxKfiEI7D7id6uWZx
U/n+sl1LRbxgIURuN3wqJKX7egMC5kMJrnwngb8zs40inOrA3I+thdyV4DyNyNrjz9RU9Pj37hVZ
gcdwlqGcFXn3/X/vvS/JCdBYQoFzRA4MktcIhUL7aMAA2w0XP7mQS6EC2YEGLKYHjD837c4mqSdE
huttverubwhRaFAg2CAiiyz1kYER48YntVJgsrW9UWEJVEwVeiRrkvU9mSIqecIUszJtXoFf4I2R
KMxUDVigdd8qZarwHXCBW66BJ2NSkJ56ewVNUBH14ec9bhnznyT7ZLaaXt6sfYnZ1e3OvP6i9PSe
6Wo2XHmR9SoatSVqivfnjnrcPHEhSzeZkXANdlAK6nns+0ZIvgI3lmZDWTGjFj2/zYS5ayKW0IOf
I6V5HLoyy/lqrKD7pv3mZE3td4fPWV70RIkil53XEob+u39l/2P5JrNuplO7W1w2mQAnl5LJbuFc
KGMJu968j8y2vOyHyXg0nUs4TJhh4ZO2dgphBwlmFDoxRBJev9lt/b355hWmbbemPqK9B5Vwv0mI
R2/EK7X8eL/aHg0Q5IoWKuKomylxqEn95EsrRwcmC5B+cFO6Ao2V3bo0s0TmOGOdiFPCshBkSE84
Mtu4QsequdL9udB6TngdsdWvW8+KTHJL/pAoG52UkHIqzDBpfeluzoy+eHZdDbnAPXM2hh48G0oG
wh2nILx4SBgzT9JzjbA6bFh0h1eh98izTAV2aUJLO85qcR0aFJ4og1J+BaTOJfu5qNo5HEJuWhiP
YzG18+0yW+DaX1tKc0LCTBGCKo6ipiRHJR174P8g/2qjOsvi7BSE59/Jv4ZhZPhzBXVJtJ5lVBKC
xLeyRdnSvozhlOR8kQsnFX+tfFODqt+YwFRjjg9iTJr5BsSpIt3LZQDFRrIradkw3JASDTmm2JZW
oKhPq4UC1eutq6m8mZvGfuoXjEQYMuT6hMNgQl5fW89nSWNqApdWVjWAhiIiqzggyV6i27NnaAAg
524p+DiHzd6FcByfhMIG7hccKLlCexa4SYjAV3D/VQsAh5CbTS7Fbf7/8InK97cz+SXPFlAWiPiD
NxYu63wh4Nvs2/89haxibC0/m7glNMmfuMhlJWe3uKj0zIFMex7RXAomkr0EpDVGImnwfK565Z4j
qr4G9YunhQ3lFC9PgUpkwX5YS1EAsHcHtAv9aqXDWz15uA3HG6mBtADsb5ztSt9FxhWjLKDzkWO4
XUSAaf3VPqY4ivv8Rdiz/iFyXLUtW1HMIomWnOG2RAq71g+Ri/qcxmRvDT2XW3h8CJLTBJp6CrDI
E4GPcPzO5dwhc6SV8k1FSuI3+P5OUsNsm5EofOG9cqR/394w9jPTpg1r8KdbmdmMF2wVvPQFI9dQ
LKtX1tl/xvtPcJBRmqMFwhWAEyIw9jg/+dAWaIedldnD1UTFcqjMV8LMIH2Uhcccnn0VfzuSTTjG
NJ/TAl6SeR7mwAz2QzTVENURm6M2JU8DZ0GLkNkjlhWYf5UrVvuiVOYS55QVM5dhervbtDfyXUGu
suIo3IM1L7+FTIH5eOMjF/V+KOA6EpjLa6uA+XLGkr5R4/TY2yQmwxtEoRUCCj50sh9QKRw0u6PA
RhTjDeVT+cDKU4sqD5j66u7FCnv8Jm9E8EuaTXZMx82jLh06jOVZ8Lszz+f0wWHVAXZB28y7asQ5
G8X0qLExX8Vc+kgkZg3QD94khNxThTdd6aMCyGxu7/EEeufL9XmQh/O86vXYvsoMszjRy/AveZ88
r59A5lK/lW+mmQJgrov6kDhp/dGanAismwqOl8W5F1655ND/46bmZo7iA9rDR8Cj6YvjFU7RDvwE
Jf4GEl+ekyQ40VQh+4C3Q0uZi5pf2gqXDTPmAG8z5+4j8NSQNIm0476JBkqzoKk8RZMLWwiYdVym
UnHmvz88ATtu5CVVsxID6Npig6MFoQ9yWOfwLf9pTeJ9HgLGcW3Szu9tJREcZrPL/MRxalWenYq/
SR9wzqBOkDN+C2R3MF6+Gt9Z2rtX65mfT90BSPXinaB04e8WBNj0iz2Mex7NyPIAdnb9MpLUDyzu
QQ30DqFWCG/I0n2zIIvXeaIe4yLqZxBMLzrRTbs3DTqBcpZKx8dXoSUMFD270NzkVo1MJXHVL4r6
NsNQnbTWQirjv3An6RjBuXbEcqHGtAxNF6xuWxLxnPFITgVo3B1BHCikZ8KkBY7+v6curmmUj/ad
k2wTcURJcS20ML6gxi0aoKUqUCo1nqj+ARlCuPaKIepW4IPD8E9ZEk1OTY8kfzd8h7zCW8Okf7aU
XXSOls2w4TuUa12XwEC/5spM6Yzq9Stf4BIagP5Dz0U0OVDMph6vrpPo5EIR/dunI/40Xs9x8bI7
baXcaN2CaIhqjnOzGWm5qFooPr6vrcWK9gHUf4kDP5GvglyiRY7rmWZv4RPNE9bSSySUhGu+hA89
maQ8W3M5Au2PsMyV6OKIQeyI2hLpHbc7jL3E0TncOT53I7jfNEAwefavxESYsvHWmiTwSUBCLliD
bY3zpCFMmO5iFjpp7H6y2L8yAOTfls67ZFUaBzWxeR6xhaHZK/mUygiLVaBzlkTuwQcdA7X4WDk5
ArsoqiqlsicjIctb2iBz0MCDCqEwfmcxSz43GeKp9nQTsiKAeiYRZSQvNnvHxSvkayIojpYRRO6g
HVq7UkvBT3juuA5TOVmTAhxd9DLgoR33EyrL2CpHCK66eCDUxY7sNOtqUPJ8Tm530NoubUFZaNiu
egT9KFJCuG0TbhAF15kBiL/kY2cqb9ZRazmNcgZQ0kA7A613uynNNH8OYdJmJdQUBm137yaZPnTb
ixcfDcjlY/rq5NdecYVuCiVCmJFMMPZroi3Ol4EcGyzYwCV4lv5AQ3t3KBngk8X+FzEaChwqrbIR
pm6cbaoqdaZi8LIQ55MeTHwRrfPKhqUlOPlq4zXG3+EdcdWiIw15WrQ+25cW7PBLPBI5JRcqtR7r
9VO2vWRfcBauprGorvKvdr3TtVcsUMaMKVKgi6jcWKe3FsmjAtS1GKxDjsO5tE1jIsasRzavaeZ9
kSPJZssr7FRbuuMhnmwtgYGz9aG33TeU6QBCtsIrUOoyFsezlzaZCFZZVOtz82P4evAZJGF/E8S8
2RZm2rjydJAwvkV0OBKEaNNFPnmXGkfnrTk4AHsqTfpSzxLPrFaCmrDfDxUWuiRojmywd52CD9qR
UuMChDyyj8GkQFe9ujJ6v9YMxunhwD8lpYX1TkG+qcIPiXPD0aK6KHnJ69Sybx93Jgg7f8QKN14J
UOiAgrnq6bXb3hhKtNvD7Tcp9nqR7971cC0PXLUBB5rD4skdCUhWXUWL2A0o6FnauCutu4L/D8Ay
6A0cakVIWP2rWIKSAmeLD2ybDGTYDGch5yuKT4uaMjeGeu9HG13X0/Rx6fr0AX7a49qpSiYLGEqP
QH6kUy9GTgVTvyG+msV5uIFfH07DcTMT5DMLjd2DhycYSvxngoUFse+Ts78gsRV8a6PG5VaH6QB1
458NmnjR3p46U5uCC7w73PMXNlZNquMRtY3DlHjO7bRhOJxOR886cAxFSDw12cPy+cYnSpz14PHg
WS7ITj6sr5YNTDvIpBiVFVw/z6dlNsDjN/cet3YZcjw3vGQ71uRnqvORpKtfSAeqJHA0xNKEpNAA
fp5dkj2lGeMiNP4u/tAUOgoXfqzV82CNMBKdnOyIIqzqzrCJcgimZoolLGxOvYJcF305FPBK3oSh
0+sRsob+qm4r6z9vFB+RGkfrOzYCoX7RFuTNvAskDp3dpbLOKyIlSq0EU3cAh8ttFWgC9vNLc2Sf
reBtKq5JWk1YYC5zqRvfLuqnwuoJl428DqbjHXEhbmNub2DFAO2EhhUFGR6W08I+NzXo0RzDyilB
uAi6QGI7jze3SX/m5+eaQEmPNRsY1MNl31eHEd8L686uaH2cXzEt5ipUNGEWxLnzHuhLt7BsJQn/
S6zr+STZ7hnnbNai+SUbxwrXKXMF/oAXUNXQjiNDyw5F83JONf/4vtq1d4FbwIBlMy+F1P2kqaUt
Qg+LzHNit76KLKlQetMajJIx9sd3yHWbmJUjvczrb176hyNuBMTd9G/vgT7L5Z79Txdau2V3yqlD
voojz5EbCjimbC0G8bHe67m207K7H4O+aWp3XAZhCi1f6n1823p1Yln6d7zoB7p1Oy3Lbi//NduF
NIhPL32vOM6hdKIe9zL2adDKND8yTSUItea7Q0a6JA2Tr+6akdqbYA/9bKUsorE9sXVYif6CL0Um
dPZqSIek2CgslWYPatrXWAkLtIh4S0AQ2U3AR8qqc6FGmwBVnGMsM0eHeDhKmV7lQ8mXELBP/jtc
otQYV+3FkvRsoBAEmMD0W7ALjRPEywD3X/CSXjxlTkTnymfZFwM+lpb1c3EIJXc9NtMqQRhHnfFm
tRY5lLjO0SvPVdxxVmG3OuAt+x4e8JblJcprYPW+NcHkp3dye2FEBrSPfelo28ac/1RZxoSPqx3W
pnZTpG+oOR/2mXbIn2cTitqrYtqS3QEB6mU4tqSIwcqvFT1LHXmuqstdDV+VhhURGR7/BTCYBJAd
BuazLj3vtGEhWsqCdu7mbNf9WF4yLcGdURyKOB8G5eRtSunsDf5o6laUkUTRfuUjmR3TtBa4c6v4
hDxrwNJ01O7EdSX2lA9hnFSSP1Zc1LoG6Fs3p5dSo28ZeX7CaM+cTYMkbCwEcipsfEugpl7iF2q/
/0F9iLMzm0Qv/5MclIuk4j0twHBOIONfe+vya6dpHLR/4ou/6JUJLS2s01uwPGa7uwQNo0Ij4Zx4
89lQiM7MjT8q9NHSNyZ2vCt7UrTtdeL9QqCl+6Ct3cWQ0Wv9eJmwZ1ph0k2QLZbb3yJXHeL2WpBL
4SYH0wCDxXUdZYb9IJ331yEK/eBWnndU7uksJ/6GQRyLQAZydMfMEozEom2oesD44LODMRORGC8Z
OeOQlmho+xmZdviFw9BsCgbYFw1wFLQmyJZuZFAStp3uvQn5CFoDVAC8WZPIGmfe/H1HHuQgtEd/
Y5krSkz6/8MdA75HfWtDi0LAL6XFz+YjUvSvDeYRAGY2iBxfj0FD/kJ0N0qUiryl1S7Lb+KRyLf+
5ekGWUgMfThBCExwQa1/qylP5hO35Q3RNgjFgKVJW0krgo5k5A6Jxx6s0aZMIzplKC+3Mb5/EXQF
9e9Ge/TaFIxxtER0f2MwtZ8LlTES+aVbSMiETwdQB/u33vQUjMvIhAxbmdn4qI+d+Z+Vd9p6MBGJ
8qMF5hWdXeZhHpV8DcCZAkZ6JjJaDtFi/DWuKjJQP0PF+i06N8Hztvlh4qf98gLYZtrgWhE5MvnX
hdSIksHA2Lo+fLOriuZsPoJGlVBuvlngVaUm+W9bjlRBUKLSRAF4y5QyiybEseZHYfl6IW9220iC
7Sckt7jiLtsD+HprvfWap+7mGcMOGxqE/i7cSLvNocvL8L99enkLXzzgubcSKqXCrN0T/9dkWinl
GqPVUQjVb7rIJXUrDI/QZHg3z3TxcaNdYoD/nGwhJJ9q8eGekFUp7A+jgc/CK5qNt0Ue3S0CfXSH
mROHNmG4Vgp45aHOLxuHMU6JnDvB22T7M1sQNFdIbLVVYSEU+8uHZ8WGofRnY++xeg/PYnBr8WOr
7tvMjNo7hBe6Npu/Gz59uJezvp9NpCUhNbjL2nqTZwkOZH/yoqktNnzgqgR57qfud6pni+Cv1PEN
SvTFUsnv7sR9IqWwuDlZeO1w3SHIo5ur6bSfnl1LspP0MIimUK1+PU5KZb5jVkAGEp4hP1j5RnaJ
E2aIdmjVQYNB6wgy6kWganYvVkTNf5ATEItenwQfObXJgbk7GsL+vsUBMJVkLz/KiogYpGncfZJ9
UnffbSO2+dO/560docv8Z5q1CEQzDPXHnd1AlDlNWXGTybhcWBftJi/TNH38+54BQD9ADMWNygQl
VCHbesccyP0KGgwxry0yC/nqM5/sRKDlVpga3/mHjxw6ayHL2bbcBVkyYB4SHwUZ+UEbI/pF376W
d5hKRtgXXV2hPDChWIn1p7O0URQ0QyaTmcYCOkkiT6wHG9HsErEYTD7Mzk6nzcbjfcN89t1vUZJY
PlkjOenHASpVlWZGhaF0oDHPSAmF63FIRZtupPk5FuqfekzIdORdppn4MVWk+r54y80/Kh07AdP9
2Qm02vxEcvROH4W7leXQXQhbQjH7/e1dUEQ1x8omS1eTNcuvOPHxUoNe3F6eYvOH6/KaGf5tkEUx
vKrsP1LfGYcHyzAHTb1oq3v+mWP94prsIECftO0mfo7pKs9T1P+S4hW/tWsdFRKC79SO7ez5pi2H
zD+5+cgw5kvvCI9uExSF8vVHpLK3+M88fW55WTxKRZBnZ5HYlgeJHm/MVr4FeV223wUtFNdYumP4
wA7SieKH8V1HY8hZlfHDd4NuNRqAngX2mT2vjRW8+ii61a53ItSi7Vy5nfYCYVFI2FeNrUTF4vro
hYfvjn3hioYr2+ZPNXj2yVz7HDOBBjSqynFFz12KMN6NTKnP1cEEH4HpFTi08a97aLnE7Cg126tx
dlT7eNTFXnB/RHT1EuwpKJdKfnoV058VCEcUs8hoTNtcJObeypKWM5Gncu5NiiU9otnBCJ48FwTY
Uq7sW0XWxJ+vkxn7OOCWVrAixeTt2pWnTyNLGFg5Yl36q1VIZm/PTcrsvVEp4sutqfEk4pqvAUHf
n66O7UxPpP99fTLzUtLOoiq2DqR9pjKz/Yjb7iHC1DbuOgdcYri+0EEYyEaUV/e0tczcy/b3/sa9
E5740iIY7vVaORuOKytn+n1u+f+PgA4QbaculI6vpZxDonia57TrABYoB2MXtuKY2WKzwnSVHH2e
nDw3mICz4GuN1s48xP5D7BQVqz2QIfZI9NLgZi4RT2/oEUhtbqcBq8UT4tBCXRlUmeHKu+94nfpH
4ixlqkOWouVW3mJNjAkgRFtB1fsAQEWj4A7P2DpDTjxq7zy8aXeBmFpwVVCK5fRaWNVeD/zSlf88
tTXuSS6oaQiPcmdLNYkfmZD6qU1EV6HYwiD6AcNyeMJuNfb/c3lkx90Cs9stSGYeyNGJ4twjyHJu
be6yh8UsSe/Csl1bEngPaBAmPgKuzyxlBuS2Uw1f2E0AJI3GusudcaJruuRreq7M4GL23aPXRcMC
CFCmclYu5dSyV7yG8sgusNOz7CHOoemouyJIxNOsWIQ1SE/Cd/PHXS8+5C8dsTrQkYTsMyJ72zy0
EimWIE6xMrRJH1QJgBsXJBEkI4tswqWGQtuO7bnUiwKeLczb2XH7ypDw3eQOdvkMKSo8wnD2kUjG
nDBbQ+zcuIZrqFw3pSXiQ3Wwsb8c9itEwXUIjlGmOwKoL5j6tmot1XjCkW0r8DPE6DsG+HnKHkic
nwZrbB4PMZd79u0HAd4S39mckvZlP5fSwdkdferTewbWc+boGCIwePFm6dn/icR/qAfXgMJ2qRaG
JOVgv6Fh4XQwGC8dfK9CWesFPeD+LnN7sY/y3Vx/yTZ1mrdKUXpWzwdSmGrnVZbukCSA2005un6+
obZ2mfl4TVaDmTQexleJFwNUvXgIVRa/6RX3qwvUw7O1GL6r8U2QEOpxTNPMQKcl+7mg6ImUNfke
27Lj+Tu3h0bRLgrFf9a6DX8/vKacWB3ygyVZkLMiDbL4y6dQPDFcjfEaoicVEHnRL40qdlT7ETNL
SUphdm5ZC4Og/2Mz9MEFItiE3MLO3i+/JbqWgcy6xyqDdNO4kiJI3vSojKguytz8mY2Hsy3MnI3C
JcmBSgmYFAh4IsVIhg2uw4KihFzqEbbbY8gwgEncOzDR0GUyJL66L9bYdBT6rvrZOTFcZUoK31Y4
mKc2CAIYou0hOIvfeBwbd7ZggdSIjj1p+gGe0zN2IiCzjEEaAdool1sYNpaIw3xU46BII6npo8qC
qYxXKYZXEROuB9/r1iTPeEPSIiqtTNcvqwpoFCe8ImqTvxnMLKGLOZbkOppFlftavcsgSH47tMrx
MpdsUtR7IDdke7rWb+5YOJiAugQ0foNe0LxUkuifXAJeTWM9rqiCVqI4hwFezElz8YP5rOsaQ7Xo
xe7bIDXGWRgffZaax7eLiz5P96LealKQpvFamSR+P+MP/3TOIpcs/2/d2Kl6/XaPS9l4tQ/OB0eL
9Dqqr7LogYqelDxv0a7dzXm2Du8csJBgPMAJrYhhMttQBO0T89/m3XcWPuInGY1YVBXlzE/OCVIa
skkLdUaEKSvpRPmY5EM0NVD1OwiLaJZ18K7rMjDRr3ZrSy78uolmQEyekirC4TFEenVRSG3Xhn1T
y1xfbecYuhvP/KsBJIT3rs0g9hlK9fWIGZp95T9VfIjUMYcDiS668gPLIi1g3KKf8qqRv/PB/l8z
JgvW4JJQCHaMjgFD9U+c4RhIB/+5u94UvpaAxPa5SjmzRTad5UU/K0NgbWjXT6VzIjwUw1zDgV45
kHPs5UjiBdGYmG+OJUUzKST8Kde1dfG4W6AofaQ8JFdlE79OlxOL0t7DGm3mJl8KSjFHXowZshAs
apNOE6eSnrMdPk2osT5oh5DFM/rpdvqa0FENWqcvoAf6yFiOSXAk1YffgUFhOZih11qW/BUJNemr
+KVDJInrTC93szu2tG+aX0KV5u27214vuTgP5u1qvFNG7DvuqhF9kdmsMOMVw2ruXquCz7kUfprs
YXaehtLHp3v2IkcPLjH0VX1jZ3bhq1tH/mAxi+vO/TpgVBhQ4+a7mOCkgn/mDUSaJzUzfvEwgnyH
UPuYZsDyPrHci63jn8TY6opRWBVyTBAGzwZ5kiqaRrvdHWMB+dNtMni/sT4fjhAp5g/AuZhM/Q/z
2yt10sSNUc7YDTIQ1EO2h60cZ3lCelNsjJBwCn4hH3Bnk2WsuZRbJQj8tnOfhZLxSx78eEDcGShx
c99VxFiPPd5vpyzCyuBOwpP8LLpa3jILOzHOWHrK1pxzy8osxT4DRTOMOMV6Oc1cHDNLUryl/XMA
QDrKFtLBVW1ENuhsJsqNVEiOjkoN3G0GcjWIGaYv1jqzvkfqPauDDwRK/KfkHCzH+ZPE+9TWYNoQ
pOXXFFOCN4BnE+RBo1dsAoU9IHysFGv9J1zpY2kiZhRtHJYry/+E/k08zFrF3ilJLvKZ3HO7OhjI
sdgPPCNANGTAtjlHDRDKVFiyFwqVbc9SauR7kdnVra8AioSy8voNjrKpdrNDYdQBrv8I7JoH2MOR
7Y6JHxdFcbStHsPKOpXz2uraSdtoAeAj5erFi4nZJq/tgZOpd2UMLzSFJfv4qfLYhJFw4dpSsDf1
VapusQHLXKhvyy4y60x6MWM3On+6INFC6iyOvEh1MgwUw2k8VQL7QiKSJPtEZ4xzii5Md/VVKUo7
QaN+LDDASq8RYBw74Qq04FgRN9pkGQdeav/FrZAGLsGm99B/c236CFcLiAsEjru1cDm2lXOSepBr
KiKgzW9PdDq3QPWvjRt1g13huo+A12F3s2uYDP0tcztmLypw+EG+Ef15rsPyb3eUbwcR7BrF3pbi
ZTHDSPeM/M0DsFLCHCFPlwiJi3iSxjzy64mMuRdvO8xdZjwtRRAGV53s+UV5UIxTSQCyausPcRA2
A3f0+1YuEtVMnU6djpEo/791BpOo3oJWxccvMriiso/fabRXKsOzaE+93MHJCX9ZslAPolvUTt0Q
iW/kvlu4XBtclOeN5cToeW5Gf1ikxVvOD5IYR/MAQuLaiOPU/Gn9BS8THvrNmS0+hZIgrI5gzpUW
kMx3FyHQCh+/+8Pxo+ENT+kr0/Gs4/BaiM7VSZcdwVQmHS1FChcvHdUWhB82IJ/Ca4cCRuf5td5K
COIR03c3MdNjD3eCm42HPUenx2ra8bRmQp7Wy3X5Xd3cy+s4BKHVzFkqGvZpCq26Hv5qnOPf60o+
0BPI8zVx4wwaW9K1tG5o1pVgkMgp7Szj8t1hFcGYxNEjRbe8iiJ461gykIH0lP0JvSRTtTWSLeD9
bs+wnosITE6SzZa0B+K4QRujCCwLoqdeqMV52TB298f5MYD2zlqY5FSwd5wjRj1rEcX8hSrn5rUs
lhwnXLGXgvSThyK12v4UdGNyaw0w5UTAk+QZ2r4mkSVN661eYzdCAZyME0acQvSz1d8ynyGRLGWb
PolTJvDlnFF2sTePFaUIVKJRlk616E92vvJp1tHHdqqChkbhvWZKEN7Ql7HC0lXxlHOOwa11e4e2
oMj9pmBADqQ5i7eW85XUdSaVfYvOEZ/LotujC6s7Y5ycTVgmN3Fi7UO5y0IwlkgZ6lNJAzxGgquQ
q1pNUZMTIk0fQV95P8G2YQNW84PLpUePxylXQPQtRYMk4QujcYpfnxBWu0F9wzTHSu7Q13Ng3v24
YC4+OZIAcikTXT737bPY3sYQIz4JPSOULnqSKrVhrdySiTzUey5ROrxjOd9wHcm4WnoAbP3O593o
22vyDq1yGOzeFsHZpSL+X9eJ6BAGhQqYQZ09+LJVU3pFO5zREaJZPxN1/o8Gwd6JDU/ujssYYMsl
u+Fo+zVCpvCd9zUH0N8G1Cvux1SOXklOWXpkjGH3HqAhtqBHLyDaYVyVMGAuSJug+mstodVFEn3h
UcIRb1smLqhj9GMGfXkQYLq+iW6uBKul+grFkpsodp6N/SsJAk5rUOpDtZdVKHHrJad/xjfmZGNv
wve4qXDPteP5F2xikXAXOF3xo2n/M46gY/UTPf1dalrPyaT7xZY5bFHPI0/hK8piJVB2VMxSCNXt
+1JREbhi59ybUMUuMH/wa7R6a7rN86LZ6t2mTSDU/w18iSDQbslE5nnQHQr1Zkzmg/d0ZURqEG6n
sVMDRgty7O35tcQVnfY5LKH3hDO1nHq+DOUHVy3Og+rI9k/Ceqjytjqh1cAkdtn0/6e8Rzi1xf52
JC++BU5gJUicnahmQZuf/uWO/w5ucDfLqOgm/YOhMt+FGiJ1OneWAh9gqDekWyGAbt7jGm/aF7V/
ukN5oRf6CVAGrniftb0JQyBhyuHpCq/D3JsPRX8eG8Sf/XHDPIYTwT6sRJIofp3K8uujZZnQLoSi
2vZFXpxNduYHNlIcYqtCQKTD/efH70d/bIzf14+LgXeM/rqmFRMPXH5d/bJE1qREhnJK1q3BH+DA
0ULyBfUhL8eoeZxUNGsGNSLOhEineotPB+a9lIjWej8VS+Rfg9jaFqx3D4oE88n0WEwbZasAhQ9B
8KRKULtIM/rOn7W36JTgihN1rXnYpY8GcCSdr6uIlWO+VXeXrix6a3WuLQsafsQQ4DMdr4CjA7J+
vWAZnTogXEUhz9IthsHUT5Yq/F0nrZYEZsl3B5r03hIyvzE+zvHqUbtUi+YAINsk43CfEs/98JV0
yR1t1zbJsN6pKjDJxKmCnF/dX5ShCwxyqRYQJKZyGfzgEEz59YSOfH2psrbA8+CrSmvpFKk97pqZ
3brSzn7eui9wTOwSr0T/+TQZWk1cZX8SIfYGBd2wHRjFgCGXtwx8HZS+idI4+55ZMB/YbQLnuUYX
L1//iZ7/50VvoCi57fNWd7TIGk0PahPrtzSOxp/1bP8aTTLcwlFooFHsT1qJrnAERFele99mj0HD
rw5FUBVh27rOvvQ9aYCPhVjyvPCCoulnhHkOd5198+Afa/AzmJbTZ7nb6KVvqJ4WY5TxiTNB9kfO
swAcYAr3d3VkxlEvyVckBN1ruRGC+vXmKKBG0abpIR3q67BObuHYgp7Vfyf1+kIrdNDnnL4fzeje
10G94ss8CIrHpoVMVWb/jmS5u2yoe1PazLq0QP7GGRgJdKqwqNXDm+1+TxJVZ1LDSbLfefHM/JGb
VGucFUWo9PksmGNihf9n96bWxrRxu+KVjLjrQLjoU5nLgIgwGWCmRv1n3Q3RHFcgdg9RI6zyOf7B
o+S3fvCpkj/ULkjIBPTge3a0Ot9BQh4nicglO4VsnI5MjohLnOnGJX7XWqFMYyAL6E8QfKoP3gNj
eM6vsYDpoSHQlI4GOTrvp3AxwPfmROnH4rDTE+2hZV7PeOkcBI1eC3phaq1YYHpfliWrp+Lm4ATT
ruMbroq2HtEp4J4H+XUUc3bd2j49xpvO3RO10qdRiVdmdQFhdx1f0TAjOhcmh13QCWMvq+k7no/e
/QB/yl4v+tvJvuRkzfS1dQM3qKdXF57ypMqsvc0WQl6JEyaGUjAzIWNxZKWZcE0oXqHKcS0qZoCP
xnnkUXpd6690w39v2SMDzcN1U4ryQelnHur+qGAvJmeWY4hV5CobEw22Gej8M1ExAKxm0ndE7iLh
VvVvvXvvMR2QOMnVQjHJZFhbAJauBVzb8zArE5TBBQJj0tBxRqlo27XmvlifjHqaKsaLBmsMEyxa
rF2IKiXt0sbsuQb0az+KNTcYS+g9tQ+o+syVj3LppCw4DWOw60JAXlkz8xuqXqtEXftsfIjMopeb
62patxOf5V4WKhAR1tMEmFn6me7EewWnPSw59bceFfm0HK2MrjsZu9HKEC4CmX5oR5dVYAl8I8Ad
ajljbkCWIC/Zd9GNu1jcqkT4VQj/6erjznaZvUnYdmKnHug2FAf6k59rG1A5lUHkGGb/1XhJUbwq
Uxsr/kZbkF+5v1tridisxkqHEg94w6HHOWIxTNaZO+xorpkWdpuDPNIqaiXp52msZAqxQX9qLn7q
xim8xWmi1dsH0fKrzjyO9kkvEmMP/NTQIBH+E+THSVRFBN+IP9Du0uDnTcWmZdFf47FxEV4ABskB
2Mq3ODSyNkoAEpEQ6OccKpehgD9fWzIOqUeK3w1FoPbAmAdFWIl/P+PGd6AojYe8axqYi+oVdXT7
JsXMHeSfr6fEMra9oK6ulERN9/cmsISOuQGII4qXeGOlkoc8i8E5Uc7ue9430hhqVl5DYpFrsJy0
nJkrohBla1fHGhoU5F+FYvra9akrINAHbwVY+BBysPZHGORQ3KIa22DI6LAU6UBsE+vCSLPZChL9
kLs2imN0ZWAIxKUdXFqyXX0YkcjzsoX1zeFH9dWRw5wLo3pFr8vknRlHiRalQgXBcpkuFSqUseDG
FchSgGuYsz5U4zeL91qJDCx2fuxyA+HanCMW5REHVrOUMfLfkyFgjhuwz+IyYXM2UuZffUQXmrKN
hTT2zwPANfLVPe5dPUDykP/9k5dU/CmqUoKwRPqjZ47d4qdgAN/En+DeyFEd4+Of0YAn/zZCtrEi
oonhHyDGXvGLDXE15esQzNzAI93X7WhT9isnoIy9R3ppjDUmssKPXANEKrkpzcYvAfKM9wAp8wjV
eSMb/iU+qxh+SFZ9661n3yAlB1iRuECl8d5KdU1XBnkGH5kSHTXClYfBReSWUz0JqcL4hS4mvanb
wP+wAIrxNhqQnCT1wyO8OS8P4I90UN/HTyp/1hYUZV1a5IvHK5en7D5ydqzP/nh+dE10WKzYlhrM
WXA/Z/SneLBu2OAJYY8A4B0pkXqUgxTrvz6wLRLPVhQWH0iY30jxR4KuVq2kZXX526szKVmT8w+y
EaaNUHnpI2e/Dw/Lf+UH74O+BPg1UJMYwMGViwOPRb5t3gpKLHWV1welbSccWrf3XHpPNe72OD5O
dx4wSiRLMxGm2hDKNlXy9qbSnfTxZE2qkO3gWMSy9FrEOIS8qo/ujiuGEYhTZVnDw6/j5UUckAg1
sGsEEmY78Gcl8dFvkCw2FWgRKWDB84+Bnb3jggvbsB/HWtYhqgqoFAZiG82n6d3ByTpiPcmsNSIJ
I7Bt3R8WCw9s3XI479s6arabOSfAJrdZvlso8tNd3nwR+lGrDkWoDNBv8EH/nvKB2BFNEgNsZuZy
9r1ufX1VIyai7gjAIduY9JWNXZ4fMTIfEA878I9GGnorq6HeZ4ypJGXHbMA3NaBVUSAzo7a4oKbw
G2niq4hDg91r6DE/WkVL1a5dRkdG4PXr0ZoKfshjdVlA5Da/BBjhXGN0YrYDAo6I4TVxISqL0Ukc
dY1JKj3rNhjND+hufVBqbzHHJC76sU6qjrgcdbunC1Pv6XHleZfxX/sCjFpPIbDiPx7HJ6YHbWpK
m18qS+/VTIPiPDmrFi03pXr7YtHr/suiuLrV98GPNWszuqZEL6vDd3ZpJkAVhn9YM3JdEVYXnP1D
kv/tFkLdQwJiJClklWAD4BFUqAnZcsinWBvZiXtAqUpRrynr8i1Ny/7l9UgvHVqT0y3DRcPkderj
ndZiHm3metR2/CyKPH95xRzynHO8m2m03hFiJRchbDnbSrMKze1CpwaeGuMgog8eIobd3h/AiC3v
movgS5flZ/7+VnPF5VG7RNYZ7tQpuMKlGmPlzY/93TwiDRgpAli+5tXId1AIEVqg+I4qduJ9Qhub
I/ndONmilaun8+vj8HpFcWqVhCv4MZEvO29dO6tHNrJhj0hnV82Xi9PiKjw0mSOAffY7XRrkRRgC
mnnLn3HJiFdrBoUZQEfMGIvbEKmAQjE8DN6FSPfvyje8BV8Xmr8DI0IVKfrnfOIDsArdmOXvXhb5
QCA0lOd3bLeHkHm3Urr20o5dVwYVIhB7HlW5k/YlSwddVaRHyweD2HFBQEwzAF/asvRI2o8RuRFD
yobMjCSSHqCQHfrL0fo5irbCAL7j51mE3yfbz7G0/F4DZNATmbMvvLGkXbIomFhaB55ikSIV8X8L
5SminkoY7oMzhMKNi0xQF4h2dQbuBkb8FjcNCrCR+/52TATpu6W3viM8ruNOpifd6tnzN7rY1AlG
vXTjiktRD5IRjpgW0X7b0jUc3SiHGa6k/vHE++vnBOZQ9S0qVi0nX+yQE+PBqFCvE3uFLgTzbB/m
VUSVCWmOlUg9Y1QWwNxEvdT8a6s+U6E5PXd7/GEStpqTxi8ew+w4RokSE+3sBYdlhChWHNzEpJIn
pwrJLgl1irkbWC8m6ELb52byxQTxjxdLCaFGCotYl1XvnFMPIeUmHcnF9CbuzXrdpxGeS55eTSXl
m2vWqKA/x1Bk6ujAhUC51lAXsT1rGoW2FuZix7X+bIAAdc/4zskpsavE/Ff1eaZFEB2g+LNZJ2Wi
eOn8UGwMpy3Vu8FTFRezXP9A9TjfOwyJFXAdX7ewJ5wgDqXLc+sYf2RAAagauTz+2vuqZJ/KyVcS
WXF5ltWUxk/h+Ae5kzalIhLOCzLrogCHSlchyj+NJBIkw/hW9AzcgpW88jApwp6avsZz6ms8+oNd
PHa3aMumrZL38GfaCysRcdP4njwRiTk4ErzCsklCIYTVevu7VajP2nHSFMwK8/wdX0eIYO59Z46I
yb8o6zthy7nkvUj7rsERQh9B2XqV7uspVSGC4XFVge62UqjSNPcuBfcuBKJwxytC7Gkl/jcy3B4X
HOXUxtuqXWVYQ0r+mYIREjT0Q2q4TyvIMWOAak/P31yH8FejIVvJzCEOXVYfUd7yXenoWmcGnphq
SSYBX0/JKNLIThrpuBAoUf2CASs37H19ngWTp8pe3IcyRrsaHleeTdWZn9MC7qb5WCBZ8g9IGuBI
wJUNLjPMPz4+qdI3PbVcuLHJgoOzaS9cyqomO1zaTaqBH3Fqsz4Qt0M5+Gty+j2U6fdhPtLYVAIN
4aTEvo/cxHFoAkvZd0Sk8SIgHjrjRTgZYpae29wYltjW8f3iw3I8Az3GpYATc0OAL7wxssHGWovg
0v9YpJFHJBsKD+Ghep2o+QLdGLmMzyUyc50YuQ0Hwb7rttsXqR71luWdO3CMVwxv/JXBRjSnCmv8
l7PPdBP+YUpuUb87SP3+ke5bGPYvzDtD7F5H7Cy5YklP8VaKzwzVPv+d+dkfnEH0TJS9Jf+RUdOJ
5GYXu7UowLeoEI3TYnnYBU56unHwYfhMypeMY1Jvd/HtNtqxjdshk7TtArtqmF5m6wtPmnWbTViL
KyY/16Yk6sUXAyRdIv7w2y3z5T2jk2hRIsY4JQudpgD198wdOFCZnJeUCL6oZYlFmoE/JKJfxFfI
qNqKMRBDyHrD2IIduIuPXBZPMIFUU4Bt1cB8D7bNWetJyTWEP/Q6bZ2UtBk6TZKTqAdnzDg5GK4P
ffcnf2xpmkmj71zc28m+dLTpSVi2qLaDlPgMrUddLDV0i6evctInCnZ9kq0U/G6bPEvV8X6cQlRL
xIuMQMO82QaOanQrLpWHzdSYry03kdf59WkhXrj7+vz2wbpXHUXC+mQIGNSMHCBZhylBin5DPejZ
W6I+7F/O04T7aZ6BbTUgXTHHBia/1GlpwBxt6bm/1R4KFCNDP0NkxLmoOEj5D97HsbFJTNlxK8at
QUrjdzFjJp4CtHa7tHjgnPQQkGnPD6ZAOWrKA/rGc+SIkN/YlgPWz9rHjVkCOKoO2PpBIVJ715bU
1iabgMk+IVKu8ML0Lfs3J05Nks6XT26gqWcipuROD/66VvlIFc502OIRDKNNsw5yssSUyWjr8qTo
BCwdsMeQP9swI7D6XKbF0VUqn/4l0L6ooaElCWxx7Ma3lLJa3b1i2PPN+B27q5R42Ad3twWuBzcX
ala0lFnbBHMZEGLfCjP9JyxiRdXd3gWbpzBBWrgMgxsN884i1DB23m3sVhJwlwg3nkPUcD6vLUaG
hlXzQuDPRxZ6v3IhmAWVQ+xsufiLF+twPetlMdnzSdWKfs/GbxI/x1cS2E+UppEXny4dUHLuRTUJ
jHSup841BgYmryZHmcuC0v0Noi+dBv1JDpLbvBxSLKQvBO5ya/08QSN2ecBrNJF3ENZhjDf4BrOG
lp2YuvywsUCd/3nS89PotAZVsepyzuB8HNs4SgTW0ADbe8JJly+2b1fziI51o8fBzkXNkRD6Ls1p
ajLRYbbUmrkbKmXcqBETXE/4Fr/tajiWBndOfa0Ferss69HHLr+gxC2Klpr+SiQpy6nIKBbLOelo
Nc54PQ/LdbR/BLn+h1mg62H8/iZk5/QwYDLIp8n9EHMziEiX+MizmJfijCktXETNo8ynaZGIIJAQ
bOziz1pbCISKEsa7Jw21YHPK3/Oo39WnWwKfJwcp73yu8qHlomfslop2hvWpw3GROUte6d8OPk8y
NDnfXJDzwHXblkAek/2hVGrgbZ6JTcAqJXauqJtCA00iggVkum19qeDM1g3bpyE9CMc6GwNEtRJ+
gbbhkXxLmYeU2kN4EDMmameIgbJwnUZwDrrgcJNDZu3OEu94U3bilgkqMrT0dV4IHSIPY/qpX8C5
I+/f8LB583IzDt1NYxIcyva1ciu+Lw3noTUTh2fCB8sFRHjyP7C4JcgtNzXKaLXN6ha1gr9cSBZs
QvCQswttmVsac6eawOvs6w8sXIoRoNs8ZP+KITOs78LmyYBw4nqeJv/lHCiYccuC3suf/8RjTg3A
GQbtGcRTXyc6yH7GATWPzCCKn1ngHT/85NIO3POkV74Ee6jLV7Fchp9tn5+Ewtznktch8lEpo8+x
AcNodkq9tQRkUEWUSRT3hAYHLgDR4I96Rmk1up0btNaZEUehBu/QRogo7sabJ6QDB+g1fDEvqToJ
4FbeQ1vCBrUE3RrriLbsrZLdID/FlsqmR5t2C0llKTbpucytOjGNJQdbw7VDHjOcwHl4CRrsRE0/
bQhIcsciCKxzI+pjT6mdxjjXdhJCKY427uPxyy0tuZts9BEC3VFUvSjjamrUhuqgd41IuTzt1Lz5
DcpWc/IewCzZqFWF6KryilJcW7io4/7GvDHNWuKtUTDd5TFRrmfwlB1xuzUk0bCOR+Ez2pdNcelJ
61SDYSoD9lFII6DiXqynBWhZwgJzxSsPWoDAIF61baUT1LxfppYRQ0QIJWCEFoqMKyk7dhGj9OmZ
0hPCK8g+XVon8zGVtOXVCJklkcu8CM0swHMMNnXF2b7j26+XzGtSkx+RceRp38+wTRpW2LsLjmG2
QKr2Arj3lGmbnAHuRg693nmCpmzLg7KU/QBmDPfJwWmuqs7x5ma+uvB1mWDvev50AN8w/WIGP0p6
/6m9wKW94Ue93vqbL5xXTakcGGakTfuBxZsnV/ZvJiGXmJwCFHuOxY6Pag2bYJgh6ExIj4HKVua0
o5RPtYGPp/Bx6nG0BZ+5St5xLtAK+pjTC2oUK3qF+Y9QFXvXTlBA9aCaC6tLQOHxpweuL2i+FEr2
yEUCdgQBljO9Ez7pFrngbVcOaeo+Mhgab+hVshEm2vb6MKycUss9ApNhI27yzVTWaZp6Y3j3BGr6
NXIWQehqxGiMYblJIMmfFETbJUGMUI6lUBAIbBPPeK/KJcQXfsJORo8icvysyNeRHXIswIxtERKv
Nav3JeBTV6beZG5U3Ku6pdbAKRKU9yktsxg1xYb/ffTQ6PqSDDSgUzUetF89bn3AbytML3XXJXfp
Ee8tH8NXPA0lxrBmG4KPLZwvAoHb/xgRDSE/8/0ADBgL1uAZcE/tsXs56sYNs73GQePwAcfD/YAQ
xkMVFb/o0YbYWf2VljPwzVkoAXiphvDdbRLQAAGBlUX4s4j6PBgUGDmPImo8PWUI4WQpWNwDPHkB
YvJdTO9JTFA7p4RMzsc12FQPOl360lxDUNxyrWbNA3mrDM3bIx6/RpdAs/ZBTgtMD16mWYhAF9LE
RRvpyP/D/sjY+q0fwC5vtTS3ijXTvwHMwQZytUFTdclyxeQOJrEraHj9RvtO3G3REGyd4woy+6+F
D06g9hhbLvwdH2b/VHtwUifrAdOJHmqFkxORuzzMYPa7Ki095ASYmU7WvJe1LmFHiFL+0NpO6Z2S
yNStPWB34rCVc0Wv6J1PKvd+KGBJkQ0gBaCovfSF45t5OyDDeOuu9ye2u4hvnd5qqjIb/VWJW1Ir
m7EQFGwwm6x1bzkr/w9I5XEGmmk8dxBxCE2zynwN81sBLtEW05FUg0Lii/SobEVD1SnklwIVcKS0
SsDbdazb+TgiDhE+YXJDq8Wo3qRJbcoH3V6US/Yq2gNqMXR9SfB8q0Bnkw7Vwo7pByHI16xrAHaC
gnYVCQZh9jEVU+NiZ9R+WAdXTMnQtMTXiDzUKdrrlRLN7H8+9jOF6guqBFuvDjuCm/lHb7iwJI9U
oqkojAGpPS7sqfxVV7rLZOhhDELs75BG70MpG6Ky3mtAsDrBghKRJevF53Ssixybad7ME0mZhpZs
QFgoaSe2h9r8Fs+BMglHvWEE478VVAxvl/fNDnRw5UMwX8qAz1ouc8pEj+y+veSf2wk28bbhBc7A
9d49FNOUGCJ5peKdCQ2h86SKojPXel9iVuxJvN1aYmp/tDa/jjQquBjwTqkMh4HY0y4CEaG5zLUZ
QQIKPdlAQnvoTrpRzNs7MfEzRAQednOp87e2BgIvHq0ltWP7u83AfYZj/yZmnpLLIFUo8NGvhHoa
O9gJ09hTYLaOqbacGgjq3WxJHqWBY+Mksf57sXRHjHEnJUcYVLTTGjFEZUqdjVkd9lCkR9Ktw0SQ
7NEjv7mwWF3Hex3AmREhHM23ogpH5bs/cc0HEJzdJhMhRL4gFywiWylZRGei8ZaMjdX2gltXRhTV
MtSyLHmGEtNxCpsxWgPcPayyLagaWrt4YsFbi/gD9mEYPJyztlhGORjszzfnkoy7BndMXQpHc48y
2eFrWTM2YX/uKJ0L1r/SO/4KjRsNh5uUFPHG0wJAPTQWLbkk/OgnZDCKqeDX4WbY5U+uZfabXA0/
mAZazUoXog6qyxUCQONfeilD9pROkZsChc0oa33Dg4G6unqZm5EoyHPil8855UfBo7Bcvs5TSIVM
ToJ95FJNDr4IZdOjZXbaqUU5baAO65ggau5NXLsGKgfGPsBhVFVlkaKnUbZpfecNdJkn9C3jmu7A
/SHSh2Vw66hclKu9rTBKt9MJhgVwG/DhR54rCIFuyV1x4qu9EXJ4Rau9QzJ7r/B7Zgjqt8Uw3JWB
1bppdACF4rqwHBJ6YndxwR7SriJ9B7qMoBLR79HemIwAP/K887t1CA+sltH76oGI5/g4xGhZUWvd
6tH3AXUfBoDudLS40QL42WDx/S93UMZQ9j6rMdMof/xcZUV+i804kxKI1EgW4PmyQrQZJZxZf23H
mO5WzG4yI1uKe0FNVkk96bMZpSEzd2ewR59qHg96qRVGbWtzfyWAnUEM7qWXJf9Ft6LAMYqyI7Ov
68HVjIYzSjR5dfCw5EZYNNdVLYuk1pA64K+QMXZspcKB/lJL9S9W8jH/HHsDKDaHYv/SY1CK/ipF
ywXFMkGvbSmGpKZPpjcsN/f5NCUerS540YSD7Sy5m6zuf0SiIRVOLCSmlp5fx8flMTec92d5tk4f
bDHIFJIxOfOD19zFqoEq3Qc1Vs611yiuqBDR3Np4YbU7epZKUWlo5arotwX+CVnh7DGJpHNMdU17
dpbift4k5MTPU4s+OV1zf6wBR7rPtHojzxiZq+q7NXL56wUnhSYp/YOLKUkhfxwy0D4IcXzrS8UY
D0q9aRxEAmStVPu2nRh6d/y27sLeQ1q6oGz+phi0kCxM0EZV+z0HI7ApxNj6DfX6ELvVBvJb1QsS
pMFhxsapnYxbN1m5Q0vVKOhntfgApykpT5c3r0hOrgeH1GVtyZ1NnneP0L5w7ygkKW8Eb4nm4/cn
fIKD2StvSMrSTjCJaEo0vdzjw9hLD1dQbHKI3RAnaxRaBvGwuBs3mei3nM4XWGe1HE/fJL1TcTn/
6WwZDDJyKhiRYPw/+Fbz72m5EO1uefERlwOCwYyTAwfTL2tLme/UEaKDajgKyVVcN9zKE5Vc/O3J
yzs32Oyp0LNqe/2DsU0dfvKRAcicABcO1p04QMFpus7b3jd6cvi+KtmCb22+2SpjCvOW+JYcPVLy
CpJ1ikLZGVAZjAO8QBG0+HDRgIjQo03KTnPG1LGdsVFvX2f0rb1HSFNO/DWcO44j0uK8A3eCndsI
t2p1YRviD10QN1FztFQg1A2Z+epMelC9UEUqCob4cqWOf2b6nJfkLPirEmFZtoD/1k57gYEAZDb0
zPbuf3tOunL1esKS1NwtUOel4IyUWVNvsaP7iQG+eqBrYjoyTon6jw2AbeWSc61vaCaXIS0/JT2S
VMEi3d5n4J4u5jgfDBzJfEwjQzLD4YRz0j7TXLBjuCqCk+jVlw7wNGb/M52jk//t2ZybEmImbAab
Py0pUP3c+wNougPksDiiuw1UPmJaz0L7/3hXthL9pxUUWGalz1F67n5BKuJSRRXI1KcjFCLsVePD
FKucC7OXHDRwp5qsxL1uTjQBxDOafzVqPkNwAma/jlzwUFPaUYjI2XlM2Pe+rzLdFBN+G0adnm6i
UwFctjV0v62c2+sf2Jz4i4xVUUwA0Co3mf6Ryp0fENA+VfIStFPoWqeepwth6SosoghQi7A/QhQX
FKHSPbeCgSLnznmkL17pjMXx6Aqt7t341CcqqaeyhHqrbjPgkIeuA98wdt4pULJqDxWE77FhmQsh
yJxcYQ+9Al2pNJOpItfKs/qSnnokuq9p9kVcxLC3hey+0+3kEkM/yk+8KI86dvMX4dfd00qaZ10Q
9+BLHDA6mYPwzWPJ+0j6sXbMOlCzmjCnZlZeiqaO9flpeFVLxU8Ug8nFB10eymtx6CdK/HxSnryJ
nVzUSs+MSncXLx+85Ye0UPif5zC2d3RZyq/ojBORVnwEBg9QmvlAd5JLukWhmaa9WJrYeUeHRQn4
LHOsByOuR5mF2jjOBZrG+M0SmB4sdfvqPSsllk2tLJwgWg1y5AelrsmltSxULz5PokSRlZ2R+vJf
T4FBcTu4WnuqeHboyRdCUoYFmg4QOFvQkxt2kl/txukGwLt3uMopdaT7YHWqX9PdcLu54UQ54SqS
ZyoeCjszWyO6Os1vJX2jaoJoW4YTubS7YsURosEr2WhW379KfqTHpdi84syo282FZFT4kpZtY1Uz
X4M9vEStk9LSCM6FlcZ1aOfFlImqutTOVxMu9vafIMclzje6rU1bh4LxFV1HGWexMHKfd9/+egMX
HCcP57YJazVYp5al0QAbsd0PC8xMyAw4/0/+6Txc3uBysO/RSvyPVfL5gW82VC20Y8OsE84uwHPy
UKnST7lAzL0j1FZu7ty8NMqCvEERIaz9MkUKLrfyd+NxslaM0Vwo6fZ/d39S7WUBlyQM3oJn+RZZ
cVZvn4bsEEbK1x2TQiGa0aq5k0KRpDLWEpKquOp5sX5f7PaDkKKP0JgQWGPwoqywlwP2+JgjnXAV
vyHshXT7zcfGanf+8CAnSNsxhyUOZKV0okd62vKrQORtCw+YtWjBjHFyc30TdC3lG3WK62hVIMhO
sSdmGWJpKG8h6Vxu+MU2zAaMccOuD09svOOPdpsX7Kivh9id0JljgzrLZ7tRLmnnWoPbQTjnHrVT
+hCe3pYZV4V3NK8yL6/Er9eTOIrP83WwyJTvBNTRm3mmeyvQE078LqDHN/W97+X4vEXn+hWsj/8O
XWMoc/rYBllMeqgK6pGvx+WXsbgSPof8SX0l0F5O5tbKohGU/1BoHxGlSaHegcyLw6jh2gR1Q/8e
PrlqmyDKbTsG8oo5lIvxD31OawJ8jYFJdARJjgbVEVssSdcA8DGsYuJotnFr3LSIroDoN9JdZwTt
npUqZifAAl7XOkA1Tn0G8y7fITLwHsPCveGm5wnCQyr12oDDNDks6iwySM1YgQtdKeG+ASTuer8Y
2h83hELrvcjbYW1SWZAKbNxDhLAmBsQTFDiNCaiUESD+xwy0UyV8Yx7YnEkvQo6SKydOCryFq0ow
Lisj64AnrC7io2VcS9/9CM81IKnHX/x2NJs8jB6Q0HfeQwr52ZJoc7XeJX9jtP6Lkt7Smrjyko+d
vJ7NGbGvd2pqvNRW6/ySvKvE8O4ydvA9gprWvVUhNO8qQzEEaD55SE7ReR9Hg42Q4JWoRjOBDJ43
eFl9HIqQsQenTccKCJwHboVNxJu6wuSGKrBVVEZyILuWf58jW3qsunBGbiNEWEoIHyaC/IH2+wGe
4Ux6Zew+TQtJDYAJFzOy84L3bBm8WSckVeKQnLkZD70Ue9V4Sk9AMk3xTQDgMkOsL6Hkrbin9FTF
O4dTiyjiBPD3BiTt2c0UQBT+/qEFuTECwWbi8+0CMLMkZKC00iBL/n56i9oo1fhMbO6IccHsABG/
WjoTzoX5YPzwGiYB7kQtEgQ1FWWhI4pKnuKITLFW1Ei32pCJIlbWXb27AqYBRBNTUT3J5+V8Jlt9
bFCa0GogODxpAbdHHjCRxowxEh3gXLgoFjyUpFm3pnRC9aTVoglb18CUD1/KfPVPeAX+P7XGisX3
J+fRqdPpb8apVq6rvO8jvLe4/4FULB9DL+cyv8ZriKH9R/n3lagfsnddGiCC9S7rwLRqY7QYz4Nu
Ul1TNeZqhh3bGyvADK0tH93XjE1WZanGC0YZ9idnbvzKhZls4/f0sbrD0lIwdtGojMbUZmZM4moy
XY16GTRD9WXaaLBvuuK7m2YJnGSCca1Qzk/pjsc8MHmGQgAI76vDId5uH3mPi82OjaCaQSu10Nyk
aDMDrqOE4qbKoEBDuKtwUPWAH9pOCuG2C39ptdXrCNq1ozQYgP4ak3IR7+XpNA9zH3T4MEQlgvtZ
ozxYHFKP0VzXN8YDwN3k2qWDzTnfMrFbVulgCl14RiCMZ+jyAZJqGYJHjqk6/o/48wH3nZTEQ9Dv
I14ExO73/I2yqnUsIFuDYWJTzo89nX1voHXM/tRVGddyT+/2DxVlqOKPUBfLUQyqvR1HmIfbGYeS
84jlCWwwnVqic/DSrjrosLkcnAeaqcFEOhK5//n6wFBONvNAMyFuxyauIx4WaxmmfmKkHpsbxUuX
EhV6BD5Mk6rSiHh7883yvKJrD6s/ffc5e10/Iqxk+xGh3YocwZuH7k6wSwvwGpWtKGTV+tSHh1uR
mrFGqRGgKu2ALJ3uShqpLK/9YjyURTAJepvWsov7FeFn4Jm285E3LuP6LOMycclcSgf8qKwuPqyw
V5WBD1uicytEuVlhAA0Ld/GOMKmrKJGRPZ9fyFIYOcHamlljdtmDDMi8YydAILXrbGUvPrRXFk1F
o8FA9b82o3vRLJcJfyw7JPTRDcQNaTaruWebxPM18t32SksTM/7/2HkIwDxg/5m/oZJotO/xzXYB
VmW+9k8E+k8vcL1weWeoaT4d9UNb7ff4AMricst1JHpRn/kKjq5zYuv3qwG+wmLzIMkFOxLcbhZG
vdGuMA8gjRfdQLkkUOwC5A5uMdqJwadzx3Nuy20UQ+ohX8iJfrcMkesHAd7xD+cFydiyjpN5hW+t
DcPXDWTZnvaX8hGGm9VS+JAkJQjdNk32z3CMPe+q4UPTfD1RR7Go9mNugYGUYFLvr3mgfsL/kusn
FH7lfR9kgnbM8bf8VMKh0EmdrlkluAM8gTATkjW7ujrLIhgyIApYskciLKJ2tRL9HqeVPeQOxeNu
VoreH2uSKRawY0bAfHPZ+mtGg/UXt/h+uTNfHfJTEuuEm47Ap7fAgMltL3MkUEhyltUmQ+byCTxm
sN9WZXyg1YUcZIrdZWx4QVzG9+Y62C8dGF6SXE0ZxUkEp/zpW0oo7XqZKeShZx9zBk66bBH4nadS
W9IbL+VOi61uHOGNmHyvYbE/JOaZNZvggbz8Wytly4tLol2BkWPSxiLdvjvk9yAGtBKmj/NPudPh
UVCRxTEMx6mFZyJ1/tDeYMaq7uwyVt6Dj4isuaO7s9hSWdmqrmX27G1agq040LPIPqHtxTtOQMth
H5PyG/5L985JSdi5xaWQetkSzN9PwfxKR9ueBVH/0KDu5osq16PwGwDxxN3BftPZD8IJohmsmv2A
juCFyzS/DYs152XedBaiBKM76doCyeh9D4xPsS/deqGler8ZBgrNFybPEBhNnKLx4MPiXGFOnpYA
xyapzKgxy556zN4staxNWYOBk15XZROqoB/8PXeOQ1ZD/4M4XuZIo9opqOO46kkMT6Pawfxj+WWO
NXe3rJWWPJT5y9+JhAnsIX/OoO1ZaiLPaRiwRKXCySE17mVwiO7DAFIpoytR3PWSoTfQlxq8JpD4
UrwU5SbeYplFS4qJBKyVYYmK5dBDUo79uUEEqQXMAyQeMZ0QmNkuKkEWj+aDLbHb8sdJUJmwEh+Y
4RmNoH0U6ZMEj2Js7/sNCBWb6HIxOWXIpo4AGgnuJFGDpE3GrspDN2dTUdggO7Eb1GfW5/JU+Zp4
I5Oxb+8boRawM+9AgDE4SwuMoOlyWYrUJMB2uqwneeLp95oIqISrK7DQ6SARfZeZefoOGHL6XgwP
908mzTUjOUo6pUsuE6ypifH+MbkWn4poYMi0jhsga2iLBxaKKsATZ0lpExXYiNG36AczwiynP8MG
DcPD8FEdUw8F4BjdMOdqxiPVSZJ1KM0p/Y+p3JHA4vtQmWrLqODPr9YFhtcOh9siA3veJ3HtiCf6
z4SPmE7Duw1aLMrlTzgZrRgYig18iLL+NlldOVVlx0SWiEAZyF26BZmDFIDJup3RdDm5l/y7l+7f
PLXpqLiXkzJpQeUqYf6ryuKJpEhiKdqFebv317TmODL9+KTqUItWK/TfuzOtyvLWSwMkiH1uWoGO
wShvdyuZl6tJsJtVe3r98EnTegBBifFXhprOC9MzjcFQx9KYlDCENAYfZKm3BrBu30BWMLg9XBE6
RB6zOWPrX2HRKvj3GeHnX2XcjEwPFl2+4RZ61m+9Y4ZOu690cioanxsIYp8IrGWiDN3B9NpSC/D6
/j62ltrAkrtRbQRioNzPd43s6vFm9WxiGBWIxk0sYEbG2TFDDYW6c7opLiaEeWQjr+TSBv/Xxtym
7NZzwWWPh/GQfD/7ZLIAJ6Gisa76bzJG9ZN55RoyVRyc+NE1d5z4Ja/6usCtdT15hC7m3UOvdxFt
aDmq1OJYfaJDfOWpNTca9Fty3UAibC7teH40YzG+/H6LPxXUdNYxrVY1zLj+bQ/5dyjQr3Q/L4/6
yp6RQ7MITIK45obGs64YyOIR3corfo4QIZKJhcQlZTfhdQyiWotXmMA9DCYq+CdWvCzM7SBSZXRQ
yWezbA+o9OVK3MXv07LSgswz9QCG8Keod81xvEaEDY1nMkqlSzv38wR0HjIJF0qqb9efdm2H6AP6
7G4o7sJ2YMtU55Iey4KkmPfO4wjGI60OhY4lM8HQx7UXZ98Cs4Q7C/IrNjAFJcac+pse9QHuLTSP
djPQWr+WG7T9jyVNMRmVBySidaxwN57vmsQwpDzCq/1AmLmnM+ssW7U8kTBEyyfuSokWkVugzXY1
7GN0gO+m/7r1RPdrsDDEfkDf1r16X6SeDbRgKjUuO+g01IPDHu9AKYfJByiUQrPYoHHDH1axpqv5
cWbGoMCeidB9pftZBJi/ROuwbEJcZ2ywCjhlV5mQlURQYHhUqsc6QCyo/TFFNJxJuf6LEMKx/lcg
JnBxWCxNf4qvYTAGxAHlR26zJVn9+HDNVSbweAEsJy4GfkZ8q3sygUjiCEkvaUNbneKM73g+m45i
v+AxIJ/Pfvm7iY15XtZD6bx1dp8q3V/1PvfzybCLwubiAQptcidHmwWqq++b06HtAx3L5uUzvam6
0TXM/QX2wiYbg8KQ+SZw6cwWxByrLcsm50k1r7V9fVZXrqdGym7Ba0MmZd7eUsT1tceoBllxK3O8
SJNBtU/bnCIpEc4KFp0zVHqwxoS6IHNmJXMs86ibgiVFJtk99L3jNvOVDNL0PJwxNmDsniVffWUe
DuZTsQ3jIq6Jp3lqh44bF50SCtHBsVobxsO+URVYyk4PZK49m+LhDDjZ5ZiHwZLLfNkBKKeHPX5Z
qarA1GnTHD56O0jjO95KaOxEZWIbODw1mX1MO8vVH45JtypaCKOvwzUR4/+bp6u5d1gVCJylQ9Hd
JJp9cRF+gWMZtZEha5STc2UvTxKEzdRItnLl3SnWlFPCGTez6lWEjQz4P/TQie8jcUCoiwrbHVyu
hDbmHT6ZFhM25HfkgISOLZ6O7z1PEB+uoAbfXD9lLBpnHlgSaMotaSFgCrkULQW2oLx31f+0HOu0
NhQLiLSmY/DJZYLVXnqD6DH0AeF5ydt8Ct/8iRZWMLBuI4/ooqJd/jUuRC/a4zjz7CCOFblkElW1
lOxh+TwRIhjstOd0UmkKUWjXAv1oV0mqHMGC0lstiTFo7moLRhrcaiMJM+ajBGMh5qYgfXxF4/qc
Qkf7wcILR3SoF70JAwO9X8BLUAHQX0cmKrVS4DPUVQm6sC6JXvOYRnpjkg+5qjkzdVVoBbEEakHu
53whIeORNNEtQMWV2svUysurP6CuLekpZhOf25z+u7y2CUFjHT48IUFNpU2xLMINRdWnNBCfrFQQ
UQFPvSHunLIRcQ2NyTzyGrQf//0uZ+5xjdTCgokC+8yeLC1cBmue/21ubaeJ8xDXGO6jfTi1AL8R
rWMXtVSy6V/vOPmUefRGO1g3KrJOQ7bytrKEFHBSrp+TXW9VbxHECF49ynTDtfm9vCxvgXXBuYZ8
BBeKPXMA/bvQVZreA5qyf5lE0H9Tqg2ahxVPahZO6IFF//ApwBS8+UUn48bhDfilTJpnkGfp3HhH
VIT7qPQk07uZwdvk7bI5u3CGqC631zzn2FWwv6i9vn5HDVlwoZg/Kheuo0lVZ9JV19x/Yn9uIr1S
nUxOJ4VNlCQ3b+ZWNvJwb/s9m5qWBbBpIt6ot6maqAx90VS/uR3AGWS1yPxcLweLxYxlmtIpB73Y
QkE7NVFC8iJ5vV7JiEUh5CCxuml0xv1wEdX9bDemqhG2sifqj0eepX/Q8yxaTIzybX4QsU4pcIhT
zD0D6YxVafIM/X1GB90m+IGXH76muuEGy50n6K5qHrCCf2h26o9q7LeCey2CUiac4jU7JOBwCu7N
55gvtgog2tNKAmltlijeHcL+TIlQnJQJE/qWCls7fM/iJnrY+TpL+QdIKbD6HvK8pmmIWvXBiDBv
Uj/K50t02u9nfo+DXlLmknhtXwwYHvf38OQDslZvn64QhzefMjnWsDSVmaQCuG5fvU7e7/DZaVCT
YR8mv1Y1kf9ycjoHf57VukMUV0ouX1mAbOy1qODocG+jm6rI6SdgyLl3mJ1fJa/UsycdaaDiLI6E
Gp2LcXC2Wcis/7HrxEa/TOQkYDjsQW6bd7bQrJTIbcJLBHz9dCVcNrI8Zrun2Ha0D1MCWYglZ940
R7e7KENGiOR2B0onu0p/drjYOuMlplxU5/RaP6nzau5v26RSKkmkqVRB9Bor8c24oSLkVe7+pRgf
BkJOIdsrj+Dvz8Coxk5xzIzC0pkZQIC/MAHoTgaD8KcOTdJapHEOdcxXeriCFjA4xZGAI97BT889
3oNNCd1y+E5qz/MKRVpoJlk9Wja6s9XwDn/FPJGVhLr62AEn0jJTH9DoTwNiz1s1IKERDIJPc/YD
4itkObGBU40dKry5vdF9vYayp9kJWjF0mhQZtRb9VcxtwRbh2LT3P0awzzB5rbaXLu6yjubctR+s
fKKVY8BkCxS0I1IK9TPr8mEAdgcb8G4KTCQqccs4c3V6p6Aw5NK0D+lqio87vIEIh6MVxFmXUE2P
SVnSKxepOeoXNqttQ3Lt70YTF3ufWMo9lDZT0i7Mp3aqWLPEcgHjoKb1Qu0A0gey7BZjJCFtdpN7
8qk2K1snLaHRgkASlYCXgasEvUqDgdwrvYPvw39OJTH1P8EQEotzrqH7EgyNoLIU9Om4I5417p4q
FfyWzKuVgvaVfwd2UjS6ICqBj4xMyiVz3fgvkCVyUrXYWccgoLDUBx7Ro329LhOBEKHzEzg+Dr6o
JMVRVDoZe9yUZiIiqbbIqjw40hb09MCLy1XY+XQCf01ZRjTktCXfaEv+VDtWlja8J7NFTBN9MgFe
IIfUSwN27P08GTSXkrTq5io9riShLMB/iTWaq+VOzAaEY1lHNYLHFXImXAJcZr8XD7j8+GVhqAEX
XceyeWI7i/B6pRuAAv7IyiH85CTtnPiwoTdFfkxu3zMPgYI7rQAh5hAIa+OhKtGnSqBRYWchGsKL
+VjKDVqIv/gtczG6DkJhFtiefD7G57topGp4XTHGz4wREs8CIg6brdaM4T6Adwxu2iLE5VRURmUT
QKaA9CD7/6TQbpvFqRUtUF65n5mDh0PpHN9aqFTvV45GkwGujctjDHS+c8eujumJCmAkIx76INJw
3SccOGwjW+zC9/JXUeo1yg+kMtlXmAjPAxh9EW8nn2oOBcfdzkzSJYKp6hlXMNB4o6jcpBtQuE4Q
m37zaunavwn2IWdFC/s71PiJwilSFcx2frxOB0+3ZMHtxwqc4+Krk4lEAegXQ9yjn6zXb3uKXGGN
QDwuH/7VoG1YB2+uNpVixZN/+C71MgDZ7GcCUfPKAiYNTfxQ+yRcuAX1PEFYU4uD3knT/Thb66nI
TheVAtIXqeHo6vcbO8AsgTnvEP0NhyGxLNT9X+Wh0NNRSX5n4wDC5pS0yjx4vY3apqsBq5oxZ77G
6aNSRy6dcfg72e0q95U75waC1N1EKGVKjCBat9QZYa8q1LNUAy1QOqWjFcaaeGTM3Z7Gtce0HrT8
0IXzHOp68Y999XALhNFMrKkqVMFyGEKm+zmDiAcfnPPT82MYB4dv9S140YY35fv7+XG6Zo36gaG6
tbTnT01WPa7d4e4jI3lIHSayn7HvTNqM+E72XfNzzJ1/s2BYcwxf3ZEqw7913s10cqnzAgHxNkeP
xLYZk92Nxu6yVer9bIc4HmxZOUvho6boJd9dwVa/rnun+wGf5hH4JBXOnd2wwVDUK8gaC1hrLG/n
xtEUvQL6rT6tNwR/Rg2s9RjyQgL6N1kfMAlHPrwBTdY8yQ9maTkNeiM9GaQvx2rPBoZ20zUvUlY3
6YgpVw5bQn2ISKJ/ItGh8mxv9vJ0yaInYlBztyoVKm+jDi+npOVDP8+bZTPJny+Av6IkhAUQX/4W
v0sdmvlBlOvsVmr6mlFiSym37iTqshlD0AAtadd5pHHMm9BlW7/LQMr/E9+kEcT2yqdiTIzj1Mnr
QRSB/D6k4lnn8B6f18+XIY0xrewcST0nRd3uPHXActbbCdQqlEzW+C87juZH6X01sEQyoLWIkFJp
C0YuXuBSR1vsWVoyfSmaz+YIi6zshYyQkxxliE7KHpv5QPe/7H6/cXbeOZ/9BAEfeAUtaM3MOhvU
GkB/jB6Rjv8ZbJbvrCYys+HHECGxwH6V8bpaHEGRxmj6a+D10/K4i0/BpP6FdtVdvP9x/eaEi/ZQ
Ch8AHSD4E0BrPS8zDAR9sZ3x3dAChQ2umEz/rAa80OOR2gsEinyl3XoJC4zFYQHWPiLSs1UFefAy
cY6a1aimtzJTUBXtiQ8+rNsStQGVK3dUrVTv4hmGo0ZdX0GJH7bBZ1KPDfqQraiXnkDW5xf7lvVN
G4wP7qusMO8E9iw9UcsUts1tYUi8UdkJXS9bdyNTQSqwMcKzKaRTd/H3MSWt75LTLX7UZFum/F6W
ICiSW1x79WwFZVGJ7b5y87idKtzN1ympVHymg2iyDB7GZnhSkvdjVJH+HT+48U0JYidBi6yoZJDc
qHCyFvIsGP67zNgcG/sZ+TIdlbC4Ump6pbbek/0jitfuB/lq/6TXueJDtMbE9dV7TaEJ5VClZ72t
45a11wkm4jGSzytQPYbl9KPLxuSRIVC6SFF//5zkYpb5Dvw3zz+ds8ovQxYp25pbW5+zKHdODStY
yysHH+YgK7fo3v1ccto2emqTUbpVZeEsdzBNgiCFTlMC6L5xohkzee2zZlVzcOPTCPFCk6nYyMsE
O+eqDcKJIpeVjc02Eic9Jktm4CZnA6hiUYWJ2pR8H8p89Ijn7BMr/M/yixJuIx/VkDxnTpNmE7cX
osOy57UmKcu/o52cswaP5H/lxU8nPaMc+bPQ/SqyPskmVJaPLakvY95g/m9zHlnVQWDGhOmuHduh
6Dlvi+hqSUAgY9/+bkKeUddK69xoKiNs/jG6bgBolwx9u1hRwHK4N0Q33dhqk8Tiscfv5XtvY4yV
AshXiMpao83v23zxOQqJSytu9qsyr9AsCWpEOJHwJpZOsdswIsPzvaElu5YE/5GmYnstyjwbD27i
ymMbe0Kep4jU3+UQaqMshDnVA7Gv7PjK6SbR56g+lL6qAgo8fT4iNH8ROzNprr4HqCofMB0tSQnc
OUnRbDRioP5vuMYO1I4kV27o+BUnAA1vLethgztIG6aZC+llg1XbHscVpkjD4Pl9pwhax2NuwDbE
nPwDgOnuPLKcfRC3XBQ4nV+Fb5l7/kSos5+Nqwr31pIvIWcH1iaL0QLcvAM1QxCVLhMihJ+/WRM9
On3Rpu4LuFY7FvYfRiXbiYnbUG+1AIgs2yfOtWyK2FC2yY472f4Rw8sotSa9AVMyDemhNU3peooh
IsHt5T2fCHXlCH/FQ1B9r5xxQsfOzBrEg/nVRsi02gDksT6NrcerXeBZYnFn80MPcEWVyvrOeQJg
zNyKoRXkinLHW7CESNcEfa601SAJ34ZX0w5dd55ytUwrVv4V091uolfoY5YD6MYiVGysl8rotLSn
UkPRwfw/VJwZ7g4CY4vAb43lufMqL8FtqypX5UsfoBVz80juBe2jl+GpTJ/8Jhk/SY0G31EyrRfv
eKKf3jIouDvdFTW8nHrraiFhxj8iD4+AoNp+hJClG/7YBNDaYXfeFhzH7usABGL30lTppjdb8gm/
swhqZe746rcutE5IiWbF5nfrQBYnfrRMsnb11pNqioMlGEDq0tSURcY0QnAvyzBkyrrosNBQ0H3u
JUu9a2luEhDN1Z4BCUgWA+jXtgvF03lL1mttGLKpnExHrAwCML+EqzVax/dUw5xIjDyY2oHacT8m
4Z6JoRVvNNYkAhr1dHaNnl0wMQnr6E1FQTjQhqG+OmUNbmNZ6TvG31GMc+b9hgpb3N8uYazaoYRB
qazDs2wKowv+At92/SXILHe/NoN8p9yQPzTsE6uAklMle+J57Jo+FECHAJzVlTDbZQeuzQzOG8I6
zP1yeOPvC2XYgwcPI4EanD1EZbPRSfmOYzp/x1ZuIy38ooj158fQsRyUSVCBhBKQgooq7qd8jdCI
d53FBtBbZHF4S2UDjjwPp5ZDBbulg5L0V0usElm6sGtvGqoSQSQfv1tA9Sb3OfzSljcOTq2pGbiJ
VZLC0g7JK3rvhVmlOJtp5dEgIhq30x/++fKQ1cDl8s1kvGzJ59IO0k6pum1Dr/Tav0U5AXhwb9Cg
tZKe3cDYF1xuD/DCrkHxlAZI90Nue4xJ1HWdreXT1qjS9jbV3RiPypFX+OAGZt0SGP6G9gFR4KVV
UhJcOowVL2T9XEB+IiUBV65VX8vpvCMeCubIjYNs392Sfd5kRBttf6JWxOqJx2VG9Tx6EYM2VRIo
Gn2X6GNWXEDRhZ5BuRe45W6Y3/ccwlN6zfpqz3DJ/aIN89yrwtrqavDbi3vTPktXQvejlSpwQ1KC
os4qeT3KMJRtFCNAqLbB/fRTEJHOSX0stuQETDQmSrZvyPJtQDktM35Jke/nP0XUj9/bhSdVAVnC
avmNFHzG4kcomqurcTRSZCkDcONY8fUr7Iq5H8eHfU3rcn99jWpX94iuiV+/0EghfhMRFAASC6GI
E+s6SI4UT7Cos6JVuJRMj1HtpNYyWvqIYqWYC+fuVP1d7M2zBi2m2P7qmVuBEHwWIrukhMtnO4fb
JBweFW7lUbcFRGrMulIy7sA4tGkPfV4SDBMTPcR7e1H4uEeEea1WPYJkhnZtClAnbSIxpSVUq7c1
7X02sqcZEe/ZlrjKESISOZMQ+tuHjfk9fKCLqAgichHqoHqvIro41tUy+06CCyR8sw5bzsZG3d73
zsDbxtwrL9W5uf819aBuR26dmnerejeKmrQE5d4MwMwgVIcq5jgaHWYPfJf29iO5kYmVVg1us3sn
1XBed1XAX2Np2f2iTuEM8qPoUpozc9HqutJWEzY3ntc3+xvLyhkoEadGYlhHL0s9lqkvG2RAYIDm
6vuQa41HDIUhGUBP2fwk7SyRCUIFjezCcUVFi/kC/0S6GYClZwmKqO34oUa4JpyKDx91xEdWl6pY
3Aa53xqkIjEr1ufzMpGbQtgbRQIy47adFYrcshHkPVu+tpOxu4iMFg7HkyCgb/pCWek0DIihrT5p
gVsPDEm8zZvSCQHRGuR4BQWc9T4K7HoJ6+bkKTM4hFs0usXs/ztBZxujo5NAej/+MP+dq/fq0w5L
z56JxJtYeOD+oD5Qux24aJsO/qRbDzsBCEDzVsM2YPNgHKszWMo9YS0xyYEZk8tsGv6qEqiJ7XgL
0dKyU9lJCIOz1vmhn+L2Ww3DCjzYle21H01aaNd26vsl0mnFKwDJcI35JGxKJk0wezewqeKc+R2Q
Psljm2zXRzEDHCjaUjOG29UaAfta4hb6IqxF/WNGvErKT/ERyeKowf4b2hkIvcg2WLq8oa1YEsGr
9vYcYVgdz+Pq6vfTmaiHY47r1SatVSTA4L2FT0r7/sII7SWfdSa27f9wfyP5SLwc3m8Hn3gdN8Pr
eU0BGFojWml4HcoWeXAR0WHGyt5dVSplEQhS0CF2K1yFMEbV6lXQBgTD64I16TcoXwQmLpeN00Ma
R2O/jmzmKDwpADmtf6cFyptiRxlZN1NMIs5DkeYAz5Ar0eSVfWueeGim0SbnZFB6Y+cVOL7Birzf
elAmCo8MSonx6kIO1Z9CblsosP//OJynj/inpK0lx6HP1JmPGXMKs2UbepMXl269d9pGh/5SNKqr
cuX1FW+6oJk6zpjuHfWO2CL/AljJ1D8q1tZADo4F3A68Mv8vk1HDa4n4fHucbyrENtSmHhIX13nm
4xFHGu1EfmZR9AaQRoV0REuHuGoSVzw9NQFkjVfyoGCv8JYeWokhBgWL6F8UmF2t7ntYX7y97K7u
AcwMOm6mpVS9SRO3iYUHmPgpDJMCYSiESR9EcixE5QTQrGMhEEzYu7wDlWnMp4T+hlDrkwaaG4br
bTEpn8umw7qvGvA1WjtdgjcqA2GvuYfMQwiF0YV0PihcK9LaD3syID0n3PDPiTqGALYrMysD6VlH
sDzK1BFw3kQHWs4EypaoKMcgIapNTzqTMS/7upA9DiF25Jaf8tlyP99CyQ33KL1h3feDgp2CMqq8
3t5XdAaBb0svki454zbte8MNxtMIZU4Q0shOzpdlbe8Hh9LpDsKLTXdHFrrz/w4bjXf53UEKY62i
C1mbbBEGND23P4W+L4u+0eXILy0wb95z72ro8wVVq3ab8xVYReAao3gNFMYQ9XyWx9hwzrtf/+SJ
qyFLXRkq4LcQs2noSPW+ntezPf9vp2DTDi1nTKBtdE6eOfzXhx9kYbbcaiFL1yhAJTjMVVR4bBLG
kyWTDE/xOcRGdBkwXpdTPYm2A8NKliG8IrCZIpmihqYky0NZuaHPmroNt7YezxbLWiDndSZ8vlu6
yZ/txKLOkz7OewATKaqs7c04g3h/5myEG1hu7hb+NB2J/t2Bm4yWHpWeZM6gtA6qUQ81y4Uct3SN
InE8yZ1A3SSsFfcEeXuWwtzxMnpiWnDQHr0wknJbEk6VnbOh8CjyInp9s59AfPxIsIgjyIFWX4t2
lQwVfe5X4EzkAcAd2sdhp1tc/5QbxF3J9y87VjD91uXd5Er1AasO6MCoGZzf9/mDVBW5pqtNiHRy
/y5WVKTVF72MpVbCtCrPQ4m5JHAUDWwciPJIEU3345XxTdwTYAHHzyVUfps0us9DWURJy6d1K3Hi
4qxeNN5L18acsZZyBKhJcIhOl1Ui2PJhtdkzJv0J5W+4vjKrDzpzIEdF9KpKfRZHN3ziRE9zpqNV
+DsuMIen6rGixGjVi8gWuvEI6rrbBIbuxhg07ln8D0BNb1yHmDFB6VrLl64Hs+DWRY5JfLMRylLE
bULIqBl7ktOfHuJ7MiZg/drKStAfisab7Px0fp6eCrb+NK3Q6VMLBaym1RQOSuSJMdI9qBVMlPhR
9WfPwvU3QPRf1wun28E8Sqd8VQ+1yVwaIP8dfYvaMp3QjoXJ0hwjsjvhRxhfJCCTT1NxoHQT61Qx
EBx7ijHUzznQiDGSfbulQspM7ChK6XYXdmf+U04nyeO1jGP58jqcVhSS3FSE09afUJdgeSalrzoo
PiZ/YZx0rltyIkwg4wgsXRsUiNYxRcoGPd+6Tk+DaHWgRb7MrO+ptF+fYEzdqwUqWftEwW+mwPGN
Yu2zK77qZ2MTh+INuPukMiebVj2DY50sMlevl/F9xtttBr1FY7aLOzzy1Lm7hazsV4vXgkkqojfK
RAORpHg8WF9gZJ297gOdkWC+lbbB4ngc2msj0roBqoTZ3+e6Rp2hYXbPJ00D4RZVEhswHRz7m2/u
hj9Kx7WYEjh/HvSedsE13g5u6p18VOdaj5O2jfD4obBRNMSA4Nv31Z/tRJ6XFZYQO4MLh2NrZyIh
T72+VAHLaZTqfFIlbc28kDDJxcTLQtQ3glapxWehxUhgXNOo6GhtiG6w9w3dtY6S/7NkBC53UfRD
iB0IHi1UI0SZ0Vjc6dlNC0C0iDgayqal48MQqlOnObrdJAunfO130gKcx6r6SqhMYa7zZGKUnJvb
Uhku2vMpjGt6mIOl0jSB7II0/BwqCEjOUt1X/fUsdcWTJQqFynN29WB16x4EgsE7ENYhJY2Dncqs
i1JV0jPzkCuQoBQkHp/DKMqsquLHauX8v+5HkPP36T9XIHuzQBj4PLOi+DRzPW21fIIEEreAxGPk
ZDwJGV4AWTmTOiIZnQfjCISrSXkazfCqvpZWlOJ5LgNy3mltXBQuyfo1xJQEs16bMX/wngptKN+l
Tg55SiECjAyKOskzw2G68wVuK4AWHrpzftdLh3i7D+2SlJZvcuVUIjEEuhmHmAq6GzOg3v6xlqJD
XumkNnjXoKmHPmODjxuDw7YASm4HdkT7JpKBZ+Yp1Q2nfpKnkLAxBEHlvF9KKbHwttoGvuD54xBx
FxLTsXruwLWj3naTnuMK3L4dL20FKbQzqfabkLb+VLmLGL1dWnEBMT7UaUlOVU+gw2w0OAc2kbsX
OWvj4v8XCZP7PgIYTliKhL3WbA6i2Bt6aS4aiALfOsTbFpeFuoMz9JvyzP/l0M9upZENr2K/0Ii3
n1mVYoZcoo4eK5485ovJwdXn34fM30X6AJOkLr8h4PI1VnX4evZcFB02eynj3LwN+AuHoeHNf3XF
rv5T6QJQyK3dzJHNLgbkD0sTOeZEm1njuZvuEh0JnN/rKw1TLQABzl07J0htCvszTeunwCQS42Yv
CT1lYBuYGo+65SJHWYXe4l23y4ZSXSu6UjVQHS53xfCxzNBYbIy0t4ytqUemX7b0faHBS0Ljcu20
T1Ru+9cohq4tMlfUgW11zgrxjgqRhoTX628IjzlYJxBLOgJJ/rIwEH2dm0NBH8mnn8O5YlYl53ra
W0Bpbw4kJk8EM8m3Et/daSzgfBBbDhiyPw5iqNHvSWbGWBm3Eo/jCwT1kh5WW56rzuxGD1IVlhd+
efvoQCRVsS0BiyiBa6gg1KwYwO0GRtsuw1SjaHU5rH/aCVKBqbfqL4mRQXsXHdyRouC03vYp+CMS
jazJt4ZN3PqgTYes6eYxY2LVlM0H8Tp3yBZJCatF6GJ9ImxIck0YCwYxKy8hIG0ZM609ooQF7Oi7
CsH04cl7gkTf5UxSClus+xO2BbIoqf9E8IdpKizYPQM0qHYKvQeIY17tQ/+H6SqWxyIZPwaBoEGc
keZrJTiAweh3+F/wds8iTO7uzUV/wtFn0Q3Dhz5meo+X7Y59Nzp68tSZ0m6YJHd8JYHz9QLpe1q8
Ao8lK2FMnC0BDdGnpbCCWTzlp7EVUyySXzmeIS9Uta6CkfKoHftF7nOqpTRbrcVERa8pTGg0yUZK
u3w164kavxzQ7XsimewrDiLL5ZXQiGTm4CmFri4AJuLV/prgZXEn9At6gfS7X51+y1lASkokloyd
EB6yfu4/Xdwpum2gfECHawIyGf1/Ngwwt5bjhD/d3fH0e012dj0xNPIZURGx+aIeAJKLlhKrTtam
Qz0wUOVmFgByfa/BPjNl9F6/dFosrNrOugLTCncK0G9hoRJAgeVUlSaDo5aK1HqKqPq/FdVhAliu
efVsSbJeGvdalOn1waGPsSOJYbno5ll03t2fwNNH85+E9rVgdFqfqd0HHgz7z5/K9HPKdSO9KmDS
kPCTKh8RprsT5SHoZ/QAqSS/AaOUu310NWu6heLH3mcxBtGsMP17Pra4+/0syZGtM1IOhz1eFWrq
21U2yNGMS0dWAHbHUN6wXsXuP3o/UX0pf2F69pX20JyQJZE2Dz+BONfVv7+g8wHQkrBkEU3J8vUt
IOtL7W0q+yx/ffRHH3Qc59yWogA8vRvqkJ8EMYRRYyMcv24QA7E4K1B61SVpzP2u0EutS9MWCjdz
SYiRcr9fUpYLF52tOp7PQUOpJqdMpohFd8mk8K6PExToUNh//Ouov6NeOVzyLRVCWv5R0kdR1gXy
vHxdD/pAAWWJzWxdR7J6wJwp4WkUwB9kmCtS6zRQu7OR73AhnUGktUbPRgEsUlnPYMEv9K57kB/e
xBrwC0xjMHSsZq+TdLMtQ1vg9q4rACK/mcoDHg/WBIDpjBsuYLPPSMqg46+GOg1tM4Ysh3PnvJlP
A0M0yfU0pvBBRxn897DcWN1L23G2L/4Lctm6pzkbBRXESC+A02O+XXcHMzUK96V9J6X8gheMSG67
/+vtJiOvY9+nfNnX5v0Hn4/Cxlb/tohqpHUog2zYoXAkA3tIm9ISrsNFnC+32Cs/+loY/nENbA25
ke4Mc0w0TLAH44frMdwa8eY+RV+Dv2d7P7Pwk+QS3kMBehzA70mFCRLehS+B+It9ldPxYQ7k7oFc
1X0X4utMdj4kTHpfqsWN6s9XRzondx/h1PfBZQFwANMwRk0Y6X40rb2Y2kiwPmC/yMdW8aa7D4PR
GIy/EMYk31sRlA9U3wyKj+Fizs7OLa+zyHgrV5Fm0sGcoFulk55dLBI6tL0YF35zF7q4LnBN9hzL
g6RlbcqPqDp1maiF1J3tvz89aRXSNNZ0iz3MvnrQLK877SWxcoQxnZklnRnrrYIE5+hzXAy6+iK+
PtKUW1szPnPmpIHJJolUSKg+W6x8wEhg7Wv8Jf08qVYp2Kg1XOVb3gUSZ5BauhOVeFOt2Dgow9Jj
GFruGxogUIublTxgVDA7z0mNBRXlgKgRFjRCMaPi0EIc1ysB+CCGg1BBoJ1RriITzB3ZjsvkgkJf
YSsz49utQGEsAS/YCYZO326sbC5zUrzviyZ8ssH8XkiiQLY1m18a3KHfPb8TUr2TQiQCwve1JJE/
+MYu1nuG8KKSn/JrN9nHV+vMYZCaixuCWdJNGghJKJR39yrRoQ8N+dNZw3YW+/wuY4pjE/bIuJB8
Cxz751JY6H3koXSv03PBZgEhTpyXCNK9wY86308KV+Iu21AAZmHYNdbsxxJGrBv7DMzXBFruyqRs
D9bm6OIKCyNeCsgLLWBZWQi4leNaSI9eSsFvNi5OcYCJd6ETo2hYL2zt3YsMILtskWN9YkS/DqNW
xoMq3KcxmD+EsD7wyY8OpFjdnI1vcJsMTmZEnrEX+UAQtGrA/g0vkex5zroYoGqiyZUV46WJWyGf
wAf/7a8qjfMW/nkFzILR4aac/AelFHbYY9alA7JI6YUGinhGpILE01VEY62KPAFKHYzKpi37BMfz
er+OXI/xTy9DhYE8JqGaH+ZwDGarCvMCXKfJetECrk2MMh8N8zYHxCKCuW1BpUZZWFPjJEmhpAal
xKqp1OWsAr/d2ORQTYaGnQGESr0atswfVJ13yCKpwLLl7YzgkbjFBszXJuzpzsZS8SjX3um/fK0G
ThP2J4ymUemJNN8xodfgJecNJjWqWN5BN49Kyhn3b7s6JMXb6fQ3YCq4woism+1NROqhwNWHh5Iw
EH0GGWIrP4686+shpqkqVA2S4TFShWJSe6UCrJW4yEwnVme5U2FIsADeXC7dT1VlRhtw79dkbQvf
lE9kIHOs05tdo8vm3YN7a/U0v0RC9jSACXATc8CgbIQslODH9+QhWIv3S12UOqVSepAl2vxs5KSL
LPMixeCYsRnZvQWFSkTZTz0GbWIHCieMW2TIcrwQTdW0RQOqLPV8kHXYiHmJMGrOSQW4YhoslNdt
RzQ6/pIZLTyT9utAtFPzXvrAKK/GhoDWX7yxlV2w9yQzRx07T8z5fHrTqbJwkqQzD+akscTilNfQ
f+u+7Pm5TOAui9Y4SI8w5Mov+pRKOJe2bWh/lW49fpeW2JJLQ4Eax3nMT/kk17ZmLLdcTe9naWmY
NteInm3TSz9VNH2k8O9RBJRqASgbXrhceC1s/tZ1wsGUmCKn2Zct/RnokxtqsYDnSjqvDb/qknwH
JORmUEun0PaUpI4LrAmp1F36z2NEhmPPuMxpj+ezrx3mDOyBECEoC6Zkx4SAeMZLZN1Of4vW0wLB
D5waPBByNV6t4xv4tQjIs4h8ib+58hrCkrVxQCIiLps65PjwheDEyC1r1e6hT1xatWOgpP4zReaK
yoO3c85OOQ1G7DMQdd2x5K19GO9TkAg3Q9WZ54rEcBWRM3YvkUnJ5J8RwUMzsiprs012+IbvWShx
/1kkouHIiA0GLlMMNhqk+63X2bXqMn/r962X+FMlBMDMtJXGEnwO4NG7Zjxc46aWcVEKCwDY+iRp
PK+9awf0HsADCrQ4nsuoDAOWWcbY+B0CD0COED1nZXeAoRfYZ6neNkQrxm/pZNS/L50aGCidLFLw
u+L+oCJLdd+MkUVhTrfOEk/8Ag+gOdPOESlpsmtwb2YVWdQKfbudmBg1bxWazHLJHhjafYwdrAyW
PJXp17LXrv2XXV9YzG3wsNc4NGK+eBfUG6JtVC5kxFzwkXF5Js6X1ea702TGSBnuqUeQFNQCFOe6
HJ2Ba8PRitPWj4jxJjEXPRZj9sYV8smVo6NCHVHcFGmOQBSbbS/zDeOMFnLwjx4tJ4wquc5px/Zn
JtDHCZlfK6qtb6W4iig71wIXUanRg1PXPV+Pk9zKMKwazN4gixmEJu3eIKAKiN1/wu9mfmDhtKeJ
jHiPuQUoETOslYvS6OvIwVmtsnODe7+0WoReKEXWDZrViOmDOxo1MapC7FE/Bfypppj4zRVnPG4B
D7Iu8TedO29ZPCk0p1Vg4Pa97FShrPjk9+wOrqVPfcnrFe8rU2FRJpv99ih1gxKH3OUZ/VoPD+JC
TYUAWpDXfgNWAf4fK5jq3juHzqGZfio1bg5MuL5uRUil0xu/oCHL0DS0qBsFgH3w7ZPdWuG4fvQz
tXUGFCVZuOpO3XZveIF86w7zTGLkEa4YydU7nwpoY0KO0QI1TCdr+JdlhdpcYHC2R7CNgTctF8jl
jY2+Bf/Oxwm//FeNK8NzFU0yNEBAm79TfeLriv73WfFRK2H/GKs3weXwA8jmMYrb0CjFqkaPbYIX
kFOPGmSJNucJfL9q3ZeoZ9k3VSSDf9DETzS/9dEcvcqvOFIu2NrLM9rioiVlZUUQoMfYCBtZyEG+
gPLOdRjfe45SRIY2SlxErA6ZMw9XjOBJ9RkviaP3Fm1h5p1/5iuO3x9NDe2kLhP4EeskH1r5Ergk
VJ9CDLoB9hDpo8ovnz6Juybjn+jWxmjyuIAVL98nGbOy5jyf5omnIu0mAQaUN8uFStl8D7U3cKQ3
Iyfg2Ul9/pFU1YUtyNsXvr2mp/CUfZvwcxjJrilJqaukq5XVxgu90KEsJ9VY/UTkbU7lo51Zq7L5
1v4ZZT6GJ/o00ImgVB2aXX5NHS9ubS9CZU1et3E5hQDRsX+s5dFwuZKLcbu26SiGIVYwoT7j2R54
oTEoGU2/zPLDlFyz16DmnmRGsCyFUS4RZ5rLTr269iw6kO9+6X9joTum0bXleU3Fq5iGhlYHtUoF
cfuTgdV9Txoa3ntnBUpWt1cHQK4tnXngf1BEXuFjYjO1mAR0Q/HC2oZ6HYLsihcfhgi5kcjLH5Go
Phl8fjh7hrDktulP0wv+15a6F8oLK+ROUIlKRRRV+H6vZZGwduUdhOVGpXhgvuOBTor1A+RBBI4j
XUuFQkWDEdLKgLmuSCemS2S/qxgv1dOi7u2L9XHuzjAisinJGEARcydvpsJfZQeB143WO/SLVUF0
fpaaDVEzdYYDHVbP5gG+z9E/kwxyL/vfqctvj6UN/enQVTrmJc9I+N0Q0YHzgZ8OmfqrwCcn6s6Q
wZvLvE82nPOfaPnorPAVZZSfbUEry2XDOH+x3RIJm61ggrPH1R8DdL03R4qmoWzvcw308n7W2gqw
zKaSH8y+ihNT/FJI+6mwihKX5iTwJ35DhmX6N9F5i72scw//FWcJsg1HuLT2/Zh/cvCz5ltMfybS
4/XYYl9zugVQWVkd6wOKtmc8jQgrirp8Lqd5MSOD1q6HAE2bqcVUy83rphbeIBbiuSnWpWHR9mi7
42l1/kJaAESJt5FwJEYziFuDN27CSYK5KsYZjj6mILsUGaH9ON8TxbbT+Xn7GsmIe/M7B8lMRI2T
RCoooGSNnl6WjGCEPLeoeWl83fau1jmxRDlqfpUNw0wpLMLIOQPbHS9lfr28h0Xy4x1nz4mf400O
lmqGkPvnTE4/X1uZ8q1NO6B/4dUN9o7UsgL8xCNDbAv+hvCoJ+6OoqftV25owxPdpT31tJYNbBKo
3r8btdmm0abWNOZF7dxAxkxRcDFUpU7LXBtoIE5mcfg+5987GVjvAvSEHdezKUda9BPOIbABiTk0
pLh0MoLWg+DNjNH6tGnNlz7gG7dTq+eNZVLT+m09YJ3EmJypCp2TzhL5aEo1y3rbOGJe2xD1wXRC
UDvaUdPr4AKvn4khGKi1eksE0IUlc2QBChUJosP7Rr6dk8d8kPMWfD5dfql9Cduz5JXSM4l7EjAz
IzCTfWHwwSEi7SA7wp+jmLJnZ3/6yGeCLVXkp5WtXf1t6c5s/STWOjhVlhK5nYJw3DNAWuXJ5EBo
aMArm9yYcsPOqGpWP+v+m5mbVR4pfwTM/2RFHkqOSK0dmIEkagoWRBHzWRnLjhe8YYwzTzl1/Q1z
xFTRQot56d7ZmNZdJDGmi8H5p9es37H4l3t6gO4FbUAWbE5g72lulGV1NPAbGDawoWkzxFwcGmOy
u2VQGAgpwWp3ZjwuYfYmNeIMwi1K3nVSrMWGXMV3xJyXig57IsFFSF1I8ud3lf9w/WRG/XHH3eWa
ecTZ7d1KEvLmPUbYkqZuSWF/EEj1LVVHIvmp3nAa2TmEa0smiR+jL4Iz67rrLfDEiUw12XzRzKF3
eIb7PnTDjQNvqdx8Be8KmzTBmD2vwzjjius+N2fjd8p0cLDG3tGtpfCNhwywExPxAwABSizc2Ivc
nmoBFdb2d65n/8JOUKWVZWbt5bs7XYW1Ir85HqH3cFtB4q3Fp1+DUIZJE4kV7gLvoN8xn63os3f2
jCrDuOeZBoCeVK0RxrZfiaxK9dNR1w0sA5DNBVDSKvzZbxY71XwgRqvGEBWqiSK+7msJMBN/63Yt
t/mX8eOE24Mc6WQ4sWnvTl2czqE3il/b5h92n56PkVbpi/VjRkT2b5TsrUkcDMFqB35M/DjZdLpK
7GjmyMQUPgB3dI+nnzVQpHPB9gfMeZg0VnUlKaFegA7F1kNT72510dxMuTrds523k0vLLjh3IfzW
unpTCuh6znFzk5BonNcq089W4ThnXoRi/TEP/XjD68hoxzEwrx5flsiBI7k3c6ZTztq+cYqzaXer
NazzUIZSTjgsu2RLYzTk6jrKIYpyHpv670R8lH5SKCqLLIXnEdk2H8DC+mHkA93bBIHMOziiptSB
PjkoKSXdAku8FtphwlksjsS7z0krJhyxClN/L5CRI5ZvSoQLlppYw1huyRXm0/XXf5RdJcHtiMEO
nZso/ap1vmgy6Ffyuo3pDfQgmDWt48hcS7M0tr+yn+ftfDOViaP3okYEF5dZkwlnHI1Dr3P6Y9Ok
wShkfvT0HU8PUDhCErBUwZWipYytWTEcTOwZu/zwAJUBBPv05l3UBP18x2EUH5pQJ2TeOmmklmvW
HlkDGdSQ4JxYRHqv2022sC1Da5+4rMyF62O3ReFt1ZxMRVvQ3mkM+NHL6XQENfSarm8D/EpZjF1h
EztO3plQbirVv67jdo8eOvwm3Y4NUPous5WqGG0+bCnw4N2u7tr4ulWEV51zBQtfdUL64afIqSr5
2bdBz96vbEMx2xvLjk1XvvLj1B30ZxeuJR6f9sWxYqfFxFys3I92VNOhqYx3S+OXo0Our1x+y005
8ZsiyfbYygH6kwxYZGKaoK6J80BQ3UJLcfBQCiLI+sGndYebu5IdZFnrvDpl0fMdB0CzH6XxvURK
f6zxBAjQFJgzyT+jZqBvujQnoc7nAkpQPKJRyxI1cde2RnRFNarEOEIjd0Nc2Drr/bq4Iy8uKQxQ
5oPMgCnZkpdGMiZsx3HkJPtv82EOvDxdp72l06yrMTK9xGRNQh4td1e1FYSckA42aMt7fcU2IE6T
zHMPxHXNlitHvez2EAnGHiSw7G4skFe3N1O6Tfxw3YGZk6kvVvPRI0WjQMxpk7mWcPDTkgOJLUHq
kDIu5Q3kjhdiF+5ExZqsyUQUE70yHU8lCxlpteppsXe57ZvI69wcqV2N15c9hzKjNJWV01AHppmE
vB7ZmeXhdVEjcY6GtT/wPQfX+bHBL866J7B1MV7D4YHLr5dutynU4yiIkIjnovte18ePbDK/327A
oWfiwsEa+7UQauMcIC2I7Z+Oci/oLeyIkNNSEujAe6REyScINz9lId0qJ+ZsBOgt71w0pedRGX7k
SQdqeRSGXKo+Dq6p9u5idn9ov8c4jw/m6tXCRY7oK3ER+cWCKgsQPYHEXfkrv5owy3AjqUs3dFNu
EJtcnXaGU6Q/mHGVrpo6viLj6A2h9LI6ey4ra99RRIzfGk27SbOH7KG7K2kKsgavEyCxSV2EKu7h
DvC2rdsp3eMgitv295xv5JjkwzPdj8QwjlTs/mWHVEuxwpUQWh1USUUVtBrNUQbellpex9eaKqPc
FxJFuthlxdwvxBgYl886vaHJAqSXpgfUsTsO7M/QMxDtdaN//XOEdVGfGqzFl1jLjGUbmAcKTd25
mY0fSRis51A6vulegE47hBTEf/5iMknKezQ3886rwb8zdZgPEZ5017TtTHJpNZkpd4klHK/4VP15
cIsjjbg1DjdcwU9lvFk9r97D/HvzqtF5fcpGk6IjJtx35aeL42FwTByHfTdjRFtsk54BF9Opxj2G
H6V4QorcUxDUrVwW4ntwea/lEEAn9PyimnZz+Dp/NpiQHgwX5IL1Wg7uddtKD8TChZts0q44IIFn
kWmU7SCBaYO8UFBK9WVDn9DKcq/IhmG6kuyWG+YvLhucnXCedEmbIIqAVuDYmFPOuasQHbthV/VO
285yg/oMlPcPghnoQaqx6tYjrX1+/FYOmpqc+9ue8si51F/dlZQYfkMjoVRULc/6j6+fKb+Ioq18
cnTAMpFLtaLPF8goKk9Lt1gtYxxnByiTvPEEVV2w667SsbDo1DmsAVoT2OiVYSMjQKXMYnSs5u38
P0wBq0qokuBx++GlPWboI+a4Loe04h1Vo7pbcIOOUVpNtJRG9hxOVkw4whAEVb/s2yxXGLIMVITQ
v2Vv6nhlHolYKvsZX8sIonBywX3T7NqgDctJxVbScV9E6q10G4GBTcfXADM4hgCx60iN60BX3UlT
qeo3IKdIcLQH3I6jtqVYnaMNF0JtfRPAEhbUBnJwKpAalJKGe9YuMgjQXmuoFQDW5P3qH7VtIYx8
oDWGqa6ozMJHBL6dwpbHaws69GWLAX3WGv4rx06nAZQFGhHG0v3Fu7uWingNbKT+cs7F64pcGETH
TJOvkhOJ+Q5wV3d4meHc+Q4rzb6ELQOKfryXqhE/M6LaY1zf6LNXuPMVLrpiTBFQVgirSE4HEi8L
Uvh+3LD5MT2ar0oDIcRWt8LX5LSG8S5gkTYr7yT5ddDxa3vrQHNJK7UwKCWq+e6NpY8JvpVyu/87
b3Gb76qTJ0kuEji3nd7kcGfZxf90ya3+oZJicwp7gTcKoCQgaowZpDk1/+BwIoPMxInesA6VYCsL
VUTVM7YHB/WURJUO0NmtdmEHdxglvGeux0fuusCKFYfhioYx0ch/gg20Hz1yBefnKqDpUi8ZHgHr
zcLX65okcJPUMXqjQ9ryMRK2oU2qGwUcIupHisXgI32GB6ep+wPM/jmr3gG/K4lIUtAimNNqkA4F
TItwash6TJs7+MwqHPasM0AFTBdDmubfdTyrtC+19QFrloAzY0tSAqvIE2oyvmNhLzu1v9RwSKCh
K7D7GmF24hDFOSWOAq8xe8seuJ8dnFiXww2H0MB+48yxDmafpMxz+iMYplHiSlnuO2CGFqEhjBfM
4UBEIMinXHEBESIfEU7Ourawo43MrpNQQ6IFdaOJmPdQd1DRiCqdGWHDsFwZQcmblZVJytiongnv
1WMQVHPU85hHf7ynP+1djmCpRECfcNOQkpvnpgzhum6sKbpZHiUuCU3EfpPTbR5EorFZU8b2yMlF
CbQYtzwD2hQ2BzELuL/114IneqFhRrcUOPScgb0PM+r1vpw69wH7RYZLClDuLXTOT6mXxcTZi4JZ
D2s7Xfp9ollEC+3r8dAR9JjBK+d/y0HgQXPvxpPkb9PXk1OOoPy6RtiowDYv8LGrRRB4XTUvVsSa
m0IA8XwTPi081SgWyBqFWBKdkScAkBtfB5y5jU8/QI+3REB4ILxNAyK4kVq7az4MX4RIY6ZP8evv
665QbECC9Wh6dQbn1ILjPiU0zZsaAdeIky6bzv6CQvIkkBNteRfzT7UdKcw3QtaffmmD0aitB6T+
S6YvMIPMK6cgqSWwbVdmh+gtZJJA5o0OdL4ThEH5eW3CzjQB7lDCgbjP1+HuIi5VMqEiSUOu51zZ
y8FgOU3dqMbDTmeWNnUWcMRmfxoXRxOrmsVD/AQ0OD95hGpYBbjPVmKwpF3sVTG95l+Ed2f3HEcu
tvuHB2BBSqGGvdZoA3OJuwTsRY6I/ox6TFkJTXosXmUTmC4JOKtyJv2u8IwUQmbWEdBcT31KZDhH
6n7aN2y2Lh2/fiFRE6kq2RGPeQpI2GxZgyz+EaEbowOEySr3nu3TC8LZelQQ6rtDTmfaz8TS8oKH
ur9cUfxM7csZDnHF+cTNx2NWyV6B8jZo66CzYq8c1+qO6z0gXGHMthx3qaAk3aqrvx6pfesxpKtQ
bVp4Ez1OxF8VNFj+kPBOy/SbhEDFilrkcOb7s1Vyv0Q/Va8wiBi+ofJlOxTnknRlb22dcgrFR2tI
Swwogn6vsy/vpQcDz5P+hNu5MC11NPho6IQZ639P5PFEk5MWqtXil6bBLY/ei3nSL2L/g8LTh7LY
AB4LPBEx0vzVyhKho7jk+Umg6j/gHCfFo9LGU+A39r8UmDqLtyoERiJ87buyxidr7EMM0XzpubEg
FuQiYGyyYXu6bAzey8hGgXNRlMCnhwS2aGWVtKD7mqENByZQcq4zOfR0aaiBx51hvdLNGRXIu82u
46VVVmikdcbOqDWUsZDsrg04xSvRQsojv0KRYkR5CJBPiN9NwpJ5uJi3KObf1ldybnpkYxNF9nVI
pT4aDFzM3ewyfGHMeMUUpjBAKTOFXdfYnrUuEx/TUsAYiBMFB6BFT7U3+8z5zZx1aY6m2bI0XSK7
4MGWWaVCHsVgXmHooBe5Uv4fAVirmffE4J+OJPsLhjVrGD4UnzklFl4AIxKTYAzelAyvAJS/k4MD
EuQh0C9jj5aCAFpQbzyrh5/FKa4BUMEuz83Q7S8/1lt8jsSc1l03JIY4YochkHGjJCdHoT4CND/t
BlZzXdrb1jSysAvabNmuS2pXwC1o7GCOMypj56ogjb/+2VEEEFdXLVqkmdFGjFe6YOLfxNl25CL1
ypYOgW+vU6SsuykvQ+A4HRT85+qW3WTLvbRFLaTyyo3AoFxB44kFTx+lXu4v4NOvzubr1mv3aY9I
9r+UUYMJHcDlWw1iIro27iqvek/RL0CteULxMp5DivdilGoJTqs5goW8u+FCzOo+07Pvo5w/9Rnb
bRRnWCdlxCdJl3inlhSYPygCT16zVFCWum7f+Ufc7zdxVEgRDeBYTerNjfOmBzX8J5KsXGwfgNk0
YbvWB159PwX2mmwpwIxzIi3kzqwjZuJU1xttpzCfMFFC1eeiWhlcsTBRLl0e/iZesy14894fVFQa
9Eyk53fBiCOsGnMTH+bKEt+UODdfvKPeSAIv3/8VodToA1FStCvFLPP0MwUoEbz2C8CI2qhGkclz
te8Kp+lLX+marz7/03S+jlJpIARVSjHzm+i6UfFds5wfEzazRMU2ei0S/IXLQNhTDHpuXI0cdrTV
3nJiwW+rwXJVI962xvPakos51/O/seNE1zW3dAYegXikKs8ibihitR0Qq4F/sgIqEUEcWzSJcZCv
p+oKRpE7TM2AybAR34TakOS1OII/F4XwzJh/bYpGHIV05qJIteDMLCVu3+adqX7dmJZzN+OyBM2W
qFc7aYumTSRtBJTkCbl6qp10ghbGfjhTtpHlgqFzClV5gmlbuYSszMX2cXu3mGhNUp/OJ3oCDxZ3
hCoasHFEOVSryFOxqSNRuzzJGNBkivlnIQ8PFMS2Khwy4UwAsrpot8wnZMfuoGKgHS/RTe16VuvT
6RQk19+2HG1WyhHojzDRqC9gihi82pu9QJzekWedBTjvKx3+CF1t4+q7tDkSfFsIrTsWHCM66xla
6rB96wXPhyI+0nm6OP/61oGE3QEK+VQs3xDycecGNwZQbTJ+TU+ADfWXh1vluGoihPaO/9Z3qeyI
JcV/rv57GimWAMx3cDUIOoaLcVBzHLv2PuKjCmoxKagYNG0OiIbvxyWIsGz1SxnUMwskGNggrLBN
/P3Wx2og9yyODSwQ6yw7/m7y/j850yvVuElBQI9tI5UKXXl3MzuYDQghOc+ME/ls6LQdniuAGteT
YuQrHTIGiCja8baimY2u8yuuQwKwURtRhbFHK5SWqhZdSzJxFcJ58PO9D9EM2QRK5YexVmiZwvS2
1962FkLtxp4GiAdTU76okXBN0auVr8nt62uIxf7ji6SvI9fzVn/UBs4yZJgaYTKmxpfoJuP+Ku3c
zUpd0x8npWnUeKb+214V/cG3iqMlUAlA+Q7HB1VAoT5QjMAXpMbB3h6M0rSKsic8vUK7/nCsBCTp
tlj5i63T+eS1/VXB9n0X7BNTL3SCysYMzqsJyE4mt+1EF5dGm6ZSR2fj8tdudc6pWmbwD9MXipr4
tzgBZmZqdpHl/Sgh0ipADKzboRrozWLMOde4rWoBNmDiLAhJSW9n+eQYrY5fIie5F89XLPwxnRDj
Z71559tocpFd7QntIgVVXeSbYLz4vufPhTdnlwlYVE4+SzD+GAJB6jy+72xHWWlgBiZ7QcGYUJmb
UGH46an9V01w8q79kVJALp8zr7IK1H4bCYT3AksN2eky6TjIQ3ZayYQHJrwSTe76bVkdDO/eAS4V
oNRQIn65SYUjKUWfYKI6ae+FtSBWEgNoaPH8BWjmeje8mDk0/bPVoPZug9SHOzWGPXdvzECDK5Tg
uhUexpjwPwyihlI3F/eB0W+tS5TXnhPTr6RgFwwStL9WJY3KamaMsic9sG/xPcJvlkVfjKWwzOvG
RWYuYp+Lu6fDgqMGZ7A8bhXCeuSXqp7Y35Z4F1HIGW8aVbRyb/+XRbV4Ld5eCv3D49C89+y1O7Nx
n8IYBxuyHzzV/kiSz+Ln3e1ANxzTme9GXeZfQLKmABqt2rAntyC9fO8z0/F1zx5amtn00+z+zj3a
5qxboJLNp1RigCH3xXaI8DD8v4dRtBEksZzyw6OZVb3K0MWKtCG6zXrLwgwUnuQT9UXqgdEL6uC1
QGqtkhuJiY1swSRzeyN2Ob+rxBbGvh5BsOVVwo7ZLpJbkq5J2livpdbImkQkHNZB2I5ydIyoVWMK
9sPo0ryAUdctkTDewK6mPo+HQCVyTpf3DVqNI5wP5aHwaMLskyyGnNQ2KIOZNidx5Wk+4tgBTFot
fxcUMV4ElO+OckBEYKMIyVbTlfk/rlGJchh0E/lI5Nk3G+6xJerlV6pAOdRtmh0ZqvG6j8fw2OoU
GWbZ1xL6LIXCU39R1a56axxNLIxpKh1Q1Op1oUAF4zTCPZT7Y9emF7zIVmZExe8cw6On5Ef4MRLH
4IwnLtUXl9uXAHRLYSt0AOvJhdm2/RNTImHAaHXbNEpZbLcXFnEjNBIetLkJyLXrzn/P8rq5xYEY
GHLMVenMcNS10vPiMmiDxmtt+wc0BBUkeG5IAzkvr/XvCmMvi3KQ6ISXoolZCl18DDfMnnNDiDCq
77srZOnT+53jtunThFE10rfMHOB44jp+8Z3uLWuLmpfJyS7/o0H9LhwJE9EDAJZs0PlmWYAPrBqB
Qclcasf7WgO0RM671J3QWRMOoNggz4MDrdXwJgWFo6h174tmNLAr006R7UEClMdlargkOWF37tXG
rMPOTt2WgRrU6e73cv2aQjR4IOBiagtdyGCO6i2F1vtofdbtaiaqKjtR3L/CAFBgRHLa9gsA73Hd
SinnawZIRAVoYH/od5uOaZJIINHPDwk7nunaJZtvLDGfZIUAwN77BYr+1zZqZzsm5VK8QfqkNR8f
SEw6XaZ4fCmuafimhSzXZfP8/aCdjHf5vcJEbVWTMK29CoBYCAcczvYIBiKRjUfBnDVGQEFAURqN
CE6UESeRpYLNRDOXAettqLy63NdOYsIv0Ws+Zcrcp9HeHqI1p0ubgX1DZ1fV7j37B56dUXXa5K0z
3BT/VKM/TPC/Pyz/4UQbKVMW7+iyn8WZRI2FHX7bn0WnnQe1cZLY/Yi1or03Z/hdMcXBHjK6NWJT
THAWYjPorFAWUpye5n9n4gAGmycVl01nRy/2XYVAAaMegwBCXk7BmbWz2A+/JJGoFAQFIqCbCK4M
+q4SVqUMFMhyqJbGQGadkOOWJNpmBa/MfsRcC1xOTr8IK2pteBbLsPlU0iUVf5y5DiaaTbz8PoDR
jjYmBbY2nF0Ehv4Mg9YoTwP/vYhgKaGJWGwZ4b4XRGAEBkVQAxRu9oQ54oWn/b6KjJeNGuQ643oM
9hnre5mVwDCS5x0LapQu+CVCDEPS4scy4QMm0+NPvlzFyTjM36X4yAGrsGxDzT2r0ZHzK6EbXzqe
Evz+5+ozXYIL7EC1y/3MhU17n5XlM7z/Ta0HrHwPYR86PUBR8EwAqvl7aPmnKm7ybgXNvkBALcmf
7JjueLptuJCD6AVaEiN/f72K9C2i8X8IRPEVWZ2dvvO76/N0wc+y5bFWdFEnaYDZL7PUzhLfSu/O
TeeLyBhJ9JK+fmyapFoFqccdDXBocEMuoaFr8KwZq2aT3ueNHQsu0dw+/R8uJ0xvCJEu36raSl9H
amoI40EtNVe9l4jMJ8Hx4hzFDHyKfPAzCvguqzm3OdT1BXHmGHhek+vpkREr8sLz8KTWwbNKDjpL
npYsz3wsk8l/XT9JlF4IyfAoZsmlrs0RS87scHDSVSWVTC9nFzhwD3982GpyQxfVSawB44A0DjJw
aBk6GkkAK+fOGCmI3O6coKZ71Q/A0n1WVPhORiEJ0fPmebC4YLVvt25AclEUVUmji4vt24kPZwcA
9WyLtxHn34Cr+28HMYNje3UxCrU/GISILGuCQ3dqsWcgLpChuHuv19DyEsXltc6/NHW6Ltbwcxdl
uwIzDXt8eR7K05xFTYGYl8ow3it04FN6AcHu//fxCL1o7YmXs4jwaeWPU26Yt8uRuDKLdG+HFv5y
D+revb8snW3p5d2t+KQnL5nN4JE8CcpDmbJ1dtaeiMkSzqNY0CDW0heZ5ZRQP+My28m7tHH3XWKC
SQn7lVMOL11XfgnuQAPyOPHbXrY6EGMB1SVdks19HNw8Gu2U8CiL/MW56utdawriSk3pNpBUW65G
uYfQbp48nmBkSb36z4T+FRCWDYWjshnJ9x+gPbwsR8Rb6UAy7RTi777nApyw8VfpUWClODcdtxZH
ZwHO/TM0KTkGKUHmY5+ielkRoT5RmJgaRadJkOQrVhoVIwonBtRFihvFnbL5bbcoovVWwyGqQA8Q
0TXNZdFq0120ZNsNhohu66afQuzxMSLNgtiCWHbhQqWvPKiESRJt5Yoo4cD3V1azPkAhYULQwBLY
G9rMCDwAnU9soyHN7yaXm1EiyK2tvg56srn6c/I9y9Al+F22McFqZSYFWB8Vm47axpLsk0qilowW
+8jufse7wn0LYYQmk1KuZh0TnOfC6K10Ni8RskejrnLuPDOoy8WvaVhHScI7Cd/5BO6v8xvO5DY4
A6RXTP8y8UtkmqsDNnqEkH3UL5ukW9eClkwyKg76t7k3C9Ezz8yxXpcos0muR935iLYWFJs2W2Gr
82lefUMyERZIww2yDBZ1N/0btR4UYV/4MsaiOJd2/4agV5kRmKtkvmlhFmH0daCSTvRGJuewK+2k
JM1rDQ1ve//IurMe2IQIdZZzPQ4EooVZO9GvsLK/vaROfF/MR2C/n05lRitiDg7yDS7UKEtihbMB
TtvbYzmMf9jYKX+k6s6qIl7sAuS1RlbXSs4Ug3zzq4+wCyCNT/10eD1T9SvXmA6XLaP3vhmhAFsw
0z+BMJhezwDjkDj5GDmKEol6tTqyavFaGWlKTv8nsXWreEJ618c5/Q4rNH/IlE0GiQ/hs5SQxcGP
ooOeiXKgxyR76VyUYYqxS7ojGQJjMAT7RfNLIenD/wUfPc5awSADpQ85P+z5Ma4/Fa2xKafOxBRg
FpJUQgQFK6eQoiLyqsTmy6iy76nyU4U+pyT9mSmxps1zRfG94p63kC1WTJh3aCdVOua2h1fyCtup
ZxjztoOBHCr3eprV3OeRNC4Wq2Fnt9O/8IbYY1oYZRDPAoQxZH34pZ6akaNtmBVo/yDeJ+c3F0CV
K0zEAYAbul70E5k7sQMfZ/JaR8P9RB6eg3ewWVZbmastjye+xIhYZzpQh0F5E3ZFzcGbUcit97gZ
uFbSwBYTDy1LJ6upKumD8oEOAEb0OfDJwtYS6cDXXPfvrebC/L3VYvEkXLq8eeU8MO9F5kRciqw+
6EJVSCjOusjgPIrVxRiyZDvsnDa5r4QQcKoYOmCxjy04mwQlacbm1fwN0tjPCOjSqlMmGKTmcyYs
ftxDV1w0lfVaLrgzBHpEiTVq2gSAygFvfzfBK2H1/PNE9ShdoB06E8UYGNY3lYi/iktP7N+tI6bj
NIRc2CU3temUtMq4MxJuSFH1LizAD6LxE7zBADYAaIh/+jMclBHjhLVb5/rdzqEnjGfZhyJiVlXF
xctCcL0+qQVeblPS0vb+FvW9hVEJR694NyT7AH1ogxcms0uGr6lAuUtyC8ToEJTw2mijMgNXoiSc
GPhtUC2RalweUsWN1EXo+WHI1UlRh/FA1tCzpyVKXwhOVcxZmRVzkVtvhEOHQekr2lRq4cXfU0dv
VBny7R0rEvi9Qq1DBa4uovRea+MkXnKJGzaI4n85WYfa+bAPkKxC4cmO+Pogr29Kc4h33mPpxqrv
c8ujMS2J/cD6uFfTW61vZKktypYrIkiApqYO0Qd14dp79k4WqdZo7p5+KqblU8Z15z2yjXlwXOUh
M6IDzhW5/2pK26IobBQrEX2FZlRDmqwfpEbtrn5bZQLzhPujdr5783IX15tQCTzZcayv4z7+/K80
zhud4SdZB8ky3aXRk5stRgLz0pt1c9YndhI61tVx7WYq17QxU50VmaRQVy2d6BomAFudo8501ARc
6buSoYrEOjBKMoE1ekLDk6Q+WQXnQsY5auRtSXzFqSG8Q6qQWMv/lKil61J4wpUm+KtnzTCADqL3
jTJfUDNN1GvUCyhrWx/Vt6BsbyFm1WF452T2F8ZQcwcx9I0f3FayzTHrIbyJFEsiBXSqrvxWog07
BCnj2jC3m5DNSAHGTnmFDECR0kwH8i+opbyiOZVJDCyBYQkfgpSecvXff+ZN8vUcDb62HIYTRBBp
EkOYhm91DaleUvHbyg57dPXEAWUsmQVSZtQc5QipDfTBoYQyD28AqsKjTQJNbSsFqouzWtri+0Fy
VNel6S8MnGAu0hncsHtClgkcMJ3r5ILEr4Dj84w5/0MMktkiV97cl8NeGBf+pwS34NRN7Qd5Z2kI
Q0jXDrssWh5KudIWBp8TmX8xQrIJtC+XPpqqgqPP5i27Zj9xOLaWBSBcIQQ8sNAJdMLKx7qB51Jm
/peAmrpARZwefwGwxKnjw+kF3JiszE/SSi+/RhvuuM3YYe9g/KkC4TbSYqmnh8JlBpHxD8qtX5Rr
oqzxwz07IOu8VymiZz/FY5FUhSExmrfpybrur6IpGF/Ny7hZO2r3e15orwibXDpWWa80KM3fO+9v
ZO9KFxD31c029X6ENYmhY6EK6aR+iTo+e1nXR+FfLyuf5AyB+sRZccLD3vVpetnHxMti+LaoFr9r
rwhEcOnDa50mSH3Pmdk3yuFG9aaQqbv9VyEowo+VOm1RbkoKSphHy1w5wmS1nivYzngl4m+WRcWl
Hs7s/zx1Pa5FFtRsPH2/a7iDMPZ3Vkv9yWZM9A+Uo+ueFTs4t6S+tSpAFfMCHkh9thg745au1ICL
3gwkR0isq6sOeLQov8YIdCZtcfgCVRwmquGoY1vO+IIiZnx1vLeQZNbMB4/K08z/bajdErPXiJba
U/BsF5ci+UxjstNzTP6TTjYpjA+CAFhLthAi0/s8JmmMDbUbrQ+O+wNPU+8IPeda/DqROzAasnuE
xeMTPSsncava77WOfy6gz5qs6dR38IqBgAdjOaJ9ttNFvv5Ve0pO6rZp/ukKXRMnztbh7yfYB2VA
dZotnvZtWCOOr4NkTP2hz2H6pVPiSLyAp8kynntXKRgY3VghGPSqe8seuR2HCoK4onYVF8QXSD3V
Ibkba95DMTr1by7XjRJrcIAQzcnKG3dYTslEVur2zbfJpHHqVPDi1JTTwK5cdGq9okymNEvbr2jE
XrZ/MR3ppZbgFlmhIYjd3vlFasNNRkYmM9b/mwgwk3o0zygHF+KV9wq/B/hpGSbnOyrAC92JcUn2
nCyI5LLZIPXYtxPysYEmPYcHcRJ155y+PpRa603ZMDDVtZ4ySPdtbgbD2AugB/kiN2eA/I0dsSla
w+DbH60sGUSnMK2KzWdcrnMTV10Mt9tJm0kS6XSanBds188zZi1fP9WlqMDLztU5/FuL0wwCHcz8
QbdtQm9UxysY8ialq4OdnpsESD2NXdN+cf1zIblgS1gvKgr/oDcq5bObKF/Kd0yOYPw+kjWJt9ql
QINUtT3uT9UZKo6CK8DEj3K0f0klPD8mjgRWDpM1xzcz/jYveSJ5C8KVAOyvCIp/X2+hIhLd+c+O
bVWZ4vrAkrC+uoEMO3c8nBKFhsjnQa5UzpKVuSBxM24hbTz+r/PyckbMwlLd7j/AkjIyNIIhHCmC
p3o/ast1FRqaghOuiJEXO05qKxgMZyRdR7lWYXJ+tCc96H4mkZf+rJ6l4ll2rW/3pexZAH4cy6KN
9nltAyQFk5rM6aPoQMl56ri8ojm5ozEp1V618apEzFaH1EmJ9d9Pr7G9b/eohpRsiAbJDdL5q8zC
nNhXsDln/Rvr2WYsEXUe5pl0G+2RAK7zYmDsYQwJHodiv7KFc6QvufN2Zi1uwVI1ZIvT7v7RwKJ/
UoRSLpC/n/A0PExoMzFcpYsen92epM+usZLWGPm4S2DDqHHmVeWQNO3YG8w1KahYSDhnnAU6adCN
hqMAzls433yY4icHhgkXKP0X+NYdd1Bv03ZnhNB/WzAIpDhsQ0grDE1V00BAylN4tZ2+Huqgi7cs
WKQSlbSjsM7SZcgR9qFUIj3AsjI9rIawxQrhGMP+bCt/O/Dd+W7FayEW1KknAXfhLrpRhCTev3+4
nmCYtU30N8YX7guo4gFM8uAFl++/Z4l7j1ugIZPmyMmSWOAoprKvRk+m3E4joI1BKRS3xJQnWOs2
oyMaEKK9+e+fAiHs4iL1E7Ybt4LVvpKEXIuWadAeJPqDES2JFgZdVNZe8WnBBZIx7AMDkn8In5x5
Ye76zE6i+XcQFUrJvMGMObD4eDujUOOsW/ohi9e2uEqb1byLSE8hRbv9+ZaCTBLSMRTJIK6Uaiuv
wAitwCrruQ5mgLjAIE+2yI867EMXsySCfkYmPiUqDb/0HdZOfKCOBDTNTa5LBco39w0CBjnSR9tX
g6GrHMAQ8FnIfLnWwLXc9q8X3gAzkjRUYO4fzbSnLErPzH9G1AFQcd3H132M/Bv5PtakNX8STZzT
WhI7flliSgCnH+HeH+9d/lit2EbB7jxqX8fHYcF1JhwgRe6hFbr7wwkwq4Xq3D8VGFE8xRFTpf4K
JeKWcjiStMY9weRiAmnHjVaBr6r+jcJVf0WqIlLcVTsID0+1A4y3cmE9YZ+40H7HAybOK3KahMLP
aEMIMElTYQn/qWaLPMECu9g65EiDBDcqiUJzRmFx5OOeZGCtjdWuvF6KNqWdxfaXK9D9V3aP2suX
7yZqJ3Ah6IHCZOD+/hjoAi83F1WTuvGsbTcVov0/gZEb4L9tZxRVzHYCMk0wod4tcFte5Wu+twMZ
Go7uYJI/VHipJCJ2fZnsPq1bAoTVmMlCJ5WUlWATNnP9Ooxw8B2mZmDIm3ua7uJWFBISL++qqk5x
TJxKjxICWe/ti05cQdFgPhCQjonAFontlrt2XQQgPHAI54XOIhXLbLuwtvkc0V5WdTUM0REqIR0V
+7S6mMqOJJHCv81CEiX8caBXf1d/lizgQhRLOkeVYZm3TuXymX7WCZ/IeQs9J1Hx1dQIj5cGwkHl
Qmw/Ded4EU83qDz+D3xzoIJsay9fbr6AqLxUN+WfcCFXeFD4u0ipCFjxH3XKwwQI+VVSAw0Krejv
IuO5h586UUc8lps0u7KgfEqjUocUcGn+Cz9KvxdSGzv1VtlVQd/Z2Oye6GqA6XEjGqcYisf+kUG0
f1THEtaQuT7GZ7cDUVh5zWpSoNVT5lDg3w/13mPHYZTnGW84qDh7IfiS99wXaYcHHi+kxLfKzaZK
9d5shtzDflOcEl576nASgrlICKEaau6I9kUaPGSF4AxhG0zqonfmJMDZFnztrUEaFoujw53FWckb
BGE3Kq86o2HMj8rLSMHTNgHE/n6Db8Wo8wQ69ddCKsBqummrznqESnUEF9QtQMaDjYFeElG4ackM
kxL0We9fldQvC5+gf/aw162CGpvrnFnmX8vT7nA+Wc+xD3l0Vh5TPLxu6qFTW2CxkAScxCxPhCo5
sIGGEVGFakdkaThYyR92StOI495k1eSgTFwgq2XXUE8Fy8EjUL60vj8+YaBRaADS+iKO72QjpPJQ
G6NEYBaZCY/WFFqeUzLuNHnEun/7HeDx0WDuEArojjRLj7wr8ezPw3q8+w39KcNHXFoI3DPl2QsO
ZaNSxPhNxkw25Rm7kWndO/Xk2OGp8tQ5RtVNM+Bo8k1s89fbEBFMA98m0hk+jMtLMw1C6Rq2QfOb
VS/7JATfaeAqnajq5ilwjNNz4aCXQS8Q2J45C27eiSGX9KIgW3YuBBqibbAQOVVw+HIfS/wrmVNV
v8Mtbx+4nFhmWfaNjmXfmAKagAxNfmqM0xjdj4z3qgRNyA00OLp0gaJEp8lqXKbHjeNtdCHcP76T
esIaFwg/xg35r87G9v5XrUhQ+jao8JTrTWsifwIPBxMR4tkGGTBW4x3fvEueU3I4W7tOt830B6eU
d0osj2Ni6wMzQn3mgAjxDBGfmeWyz8OURdVnA7gBa3zEmuSk7x9kbL8dZcylTHcoYzVaG3OXG6hV
6Anp1VWaW8zdM39NoFAAAX3DMoAcn/4Ms7RLy4MgNbnxqvfbXLByhmVhRQfbHJY5dI0x1lUS3s1c
Q9kh41nAfr/bqjrDbl3VvUugLVXedzfXLR2nYrFbEY4EmWbostzZOb9s3PoqMQost9DDa7oz/cbE
lNX4YMrpq9QGc/p8+dG0hhhZctVhwgOk0uh8q4sRals38VzmCl9DA4w00VxczPyFeMgydBFeblTA
4CA54K9wsvk6fmss+2SNdhmwiupfKXR21uV0jopYXXVN7KnD9Dtp2ZZMbY4PhTR6eFtsp02sc2dC
1nVTw59kf0GLIVEIBw9o6qGC+fQov0iQWdGuvKzAradebpJt+SN6mHAYqPIUvaw8m8R393vZ30BH
4/e+qoqCYlAMYSyw9bYKaPTot7WNFtIcSU7pP4fYU/MtCZthogNJ5OZX4NUHSnGn81c2Zej4bPF4
Fcsw338oQoMNVjR/Q81HYXQgS2iz6QHeGUlneM57qAGUEJJ2PjjnCUty+5bj8PU5hGteXpqAy6q2
zCxpMwNcngCWepMi/8NwMFUf1AWhaWOJyqdKVNImJANyuaUojY8KQ89CP7/vQgIztz182UmACtpK
kaJFxGvoHW5xVbOD2P2CSuQpI21z9YL4bzLzrtpk777MMZ4/MFTXAD7+4nJT/2i5MOgXH9VPzLcz
azvVgAg3T6N06vE4XQLlTSsN3Cefcm1h0REeCg9EauQaqtMghKgNWNePrsq25+JUmu0APTLkKAw/
3qKS/KvySDDJiQ1gpp13LWEodtoqxBOcTG/PXAyGRN6uP6y4H/284ONZcWs8Zn3rXlwfJds+Nj3G
VWZzDLZyEQE947w/pBhx+1sGpQ6vp1bAXtoojLzKIdUAhYLPCe8JZDs8gWTD/WIiWHNA8RCZyGv2
FdgKPfdjBjhaihesscxrb/qxQTXjqn0IKDng59lyB/aUjvaWp8YGWu7lInybcqn9RH58TKjx9i9r
jtgaG3qhvnBAfqKZ5k7OW01ahPeCFDvOyV8Hg8sBpxDOj1u3UThDUrMZiVQdfs5/9G8dqaMD0GZY
GSMAHNmXNwpur51Nrf3CHIz7lsE7qoJzB/CkYXbd/9wRuHgzUKwJS3kcpab7PTwrPJzaRRlReBU/
nJrOAeH/sYrMYE6hM44kkONVG3oY/sKC1k/2nkGgUUo1JfBCJGZySBk1l2ASAJxqELdCo8rY5aQz
ceDSNHfqTC1LlMcuQomrqpAJKIO7Vmrx1sJDcSRPSgRc/aXoWlD1P+cX4K8GoiRu5lRQM7deCOSX
LzOmfPAnQ5qoIBX7XFAAVMSGwLlvPYuBRBJNoM2CDtx2vRFQ+g0uYeXE2AD0xY3KCv45JtvsxSyf
zJZN/B/ep2zcrBJrQF0UO388qq+URplW4kV4X57rdjaYcFZPQsgJT0j1w4E02DXVSPJmL9j8SEBd
d7sa7pWPFKvKCphfYzueDmFbxMd1TUwqlDxRShnzuJciNv6IYZBSdDemEl1fr7u6Muy/hO1xqAWF
HnKfIjqq41woUSFAw2qPqKFOlX84dfZPenNjJl7AOJdwH+SDQX7KzbmJx+fUWoaqOV42xd1iW0an
zfBV1nb/R0XtaLRBKSd/e67kyAZv3LMR+Cu3fi2N9MEllbWDBDp06tn2rY9mSwof4Va8z5+vspt+
fXWR95C23F4BLufK9RCFBlP1dTUmfg4lkegWAh8xIkXlArrkgRt5Z0L+LcspOazgbLOnYjv/OTiW
kJGk1DyroTyh0Yea9HH56vmxPLpfIXU6NTujje4MJmRypcbnt8kJvHo2LdwOyQjqoS23bfoDZfdY
r1kAmHy4AKdZozfi8r4sv6gip5yivwXNkgRKU6Z9WcKaxkXQu+UkHO9INPqCxeY6auf+jxtc9vvU
f4ln1z2kgzQbVtXYi1O6jq2Jo9gg9nndsaJTkhhJsY7wOBlfz3iMc6L89dTpF1oMRfEr0U/XaSOe
cuUH5QWtkdd3jl5039uSt/jU5JWfk9EPBJvTtiw8RKPJsS6OBZl7qaTXTVYKQY3wx2+oVsMHnLpq
RvW5xsPqFpI7DdRJcqImqcNbe7AzFIu4hxxjsNhJAUsFroxHtKRngGbv/ZAsy/ulSG7jUyOSjVU+
61UEDXmxVmmHqKOYiQz4uYZVlIMqT61j7OlxvWYHyCE8WWeHQwE+yRZEhWFjAFk1sqZ/oXKI4g3V
p5YmEIo0kuOf648QZQ/1w09ibyvlL0KcK994HuIW5TfAIIHICIFSx/BRhb/lBiIzcN4L4td9khhG
JCuoBf6orpEI7PvZLJWkTa4iL+pxovA4uAdeUkt1aToMq5QxLrd7hj3dSoZnPRBAclTZibI93un4
WeMTEA1TxLtzhqbgyL9kmWdm+wBdvhLB7eDDJBUHbrWd9U9+EvliAZhxd7KAJF8T7PFN/fjwT4RO
cPQk64Whdx5ldDCOzTLrXjO3z5GihvMtb5J9lDYMaBImG+OnTuEumgXz/KkpT5pdv8b4notlCv3M
FcEDySaeGUqp4HfPrGOx0rcyrBdbasHZTUm6zGK8EGKuuQAZzeUlughIret8qSFNO2EWZ7qKGSbP
ipDPPGo+aAPL6pi7JRIIibzIkkLtBldaYcuvLz1oKmAqZr7LXQllZ1g/WRkpzzq9IX3wn0iwxvVX
9TZyP6Zub3p4Qb8FY6VOQKEilpb4NIWdjaseKNlC/recNxkKfn0En4xe35UNFtqej8HA9P0+2K2z
EgK7FhHCmBHGJBnLP92/QL0+znfD70TQuuX22rb+zd58wAYFUInun8Ps/3eI+mLYkQ4D30tyP0v3
jf8ux/YfUiojIliTdTQYn0JDe42N4n1SZ+WoZo20gXeNKfbKrGnftjav2+yWHRxdezMHeX8Aaa2A
8GI/s03O88myCpfWa7JxGeNc+mUTBDuMZHenZPsX0vQnfox2EfZtKTEmdU8RGrWwCLHHpSZDzKkH
XsQcwUPLaaxADsYBRmfBbx3ak45UAyuPnh8edYrr/6UJSkUr73B9CnDXgFbYa6nO72+vAHKfCAc5
eGDX9h7DqBxMsv5Plddwp6WWdoNGJilyjygdKyqS4LNJxHcxbgJ9WUxko/LAAVatCzfr4yiVy/+C
7kndSbtpnhXnOA83vfw+ePB9WZFe9PY7FUhsIKimQ/vpOgm8Upb66EpWjJQptGRe9iU91VmL93hG
+O3GfOGqIjHxD0x11pZOd0g9tK/HvRAN+emYN9ATMSm3JErjWYlnoVEi6HGk4UvkO+98z6V628Cc
L1r0OVCb8rP0P3XXhSxtwx2CteQx9GHspn6EQYByfPd+2M7r/rI76E92651zXVYCDtVUAHxTxlEu
sUE/aMlsZXoTQcvl+IeCUbGzsKL6834whnrimGe9rthP4GtNGWEvsrgPdCtTE2ecT/DdN4yR7LPs
zs+q+eyX2IS97SqdmAKgt1ZwZzTHVn11EgbNL/2N4B3o4pYgn2JkWy3gDlWFe8Ja/jcWG82tXCi6
BfgExGV8T6qpEQeIus1s9GO69asYdb9E+Rl8nrmvZ6PJwV5Ruf44WDePxN/LuiPs+bjox8UmXMPw
1luUu/lHqd9F7CESJ8nVk7PQ7H/dg4r7+vFuGNUPwA+sf/RT515gqYnTsGMASjXERMa758ukeoBf
yRMP3KZ8M/RrRDORqfRrk2jG1UVLWEBBBnq0NE9c1yv9yHSvSGzhPvXyvRBeyCaZVB9UqcC21wip
ozL/NdxP7NjGOj36amnA+0XnpouIPDQEWFTTQxmUJ93FX+ns+fvNekjCy/msJ59fV/WsC9eipYDW
13d/r72XR1YWtxGUItydGxP3utfjfqEYGCMcH5GyHeUbOWMIWSHx28PFXhxMA6UD4tapuZV0U4LU
37VIsoMLIf9N931BG3+tb1HJhVIej9YDr90Jj1yEazIDERgmJ1Caqh6CQIRGIMhdKazcyqFwIdmB
N9eK9y8TzJtLGnFm/6kdUO1licKZQUd3gQ0DurLkRRUBpzt1ZVDibMO8AiukCDVvXouknChTr624
yTD6hNwf/5jxLJxX1elRBM3l2PfWkcjIcZz7lotEbDaIMKvQbwYoxsuBrzO6CPx5sN94GEQ3olmD
Y29sRB72CZ57XeZuNKEcvqzrEypqXOOx9Vu5d9FCj3I2DD5ieXhTz3DS0fMP6E5Q9iA6IXwDW73o
3yQSUdvbcmuhSfcKQO0FuLta+tKa/h/m8Qkt1dpR3J9rMBBhFN9oGbzALgm+RuiRKtRciAo4HZrP
AsWXnwDst1EDxxWRHhsxXFuWUuz/BAXuEfa6QCH6l3tCrYE/L4OC1FmUFdxemBNPIKCuH6MY07f6
4yrFx7hxFNtARfXH6vQDVhHt5R5lHf3I+4AceQItG6TAVTexqU5naa1rFh15WLh4XINcLT/g5A07
OmfwjMivJOp2un3+jd3gIBZ2Sszl66ASScSckH4urgRZT7qS3vcWC/AClEBQqU0wsSuF3Glko4Lw
Sh0EsRi1it4fUsMxXMvikTEDoem0xjZnbXbCvOQnH7MjLZOoC0tWHD5aY2BEGJSoKjKvVNHBnDSz
JY4+8dKPTuaq2UyqL+2p2i2MUb0nBivpAUz6ocNBbXVBguTqae1JYRByAbJ4CQcXi7L4Fmu4wIh2
tQZZ2JB+WQkDMktIMkoq9LrGWpiz/03Axu7wytW/nX+TN5U0UN+iObtKppaiT1h9zTHYsKqXtWKd
ISmZC9QdvXM+LtAB3cj2TUKS+yp0y60EGe1ilqEybQ/wSG5z947qFslBhAfa3aJdfi0zdL+AN5nR
/eVsC/1rNd+FYKUQJ5qFQlUSBGRpahccii8BQCnJAJPMP9FxRkfcr6MXYEhJxSP3ECmUcewoZLpk
GYd7MUZlxC4PMOKMzuWNluiX3Y6IVBRmDdiK87xix8W5Y9rCHqZ4MIinrkCcmCG4S5onQ/7aZ3q9
MGhJAbxV9I1AJ7eWqoquwAOQB8PYyxxZh82TeAPtcU4K2LuOGAvl5tqcdmTU/GB8bybFmApXRmVM
Ud8jx0vHKHKzL9nDOMsZtLrx/uH54uJMCSVMgOgQ1+Z8ZfN+F0jTUItKSEo4Wxv5jDKo56xYAJi1
75lUUiO/hA5+MTJyWhDRC0+nsP5/M32U1wjLQOTo/Ei7K/I7DyjLnwZv1txYRt9yIJziA3KdIW4p
eH83Pi1FW1pBgURxAfWqRm10wJFznRWbVsUQQM1UXtSp8Mq8vAlKTmt/x+QTmeCkPfM3wGmvLqJt
dmDMjCw1fodlyREx4h8PlNCxvygyBROeDMK3PIrswh6CDOzFUzjBPhViYRFh+qopxcG00cABdx9d
PhGoV98K6haLPJnDGXowiluw0jnI0uzg1Z9+S/q00Rxg0WqIHWPPJ/tZkedO0o3uYS43nnATUXRF
/wVZdyL79ivRPHsB+mp5zWLQ2yAS2Pz4OFf42NLIm8oZD8EArbMyyjN/BRO37DxbiDjlpvQU0NpO
Q7tneloQz7YFe7dW2t4RUqy0KT51JpatA23aw6V2Wgq3J9CFIlhrta1HazffxwJZ0GpgY3mCHZIz
WHcOAqg+sDEP9WxyK5ew0DjwkRJb9aaqztm10ETZ/c8/cK7xg/SBQ8GsL676dxKXDQFu6vfCkIe4
bCtJeMwChG9G89CgE4KJwBt040ZdqbvRMQ6pStYP6Wvxgqw2eIVI55Tt28H8qqbErb8YNfOJt0ol
s2lZNfCG0NHcv0XvyMGatcGRV/iblTd4JyzPBQQ0DLOmLmsOlB048yuxFm1yqAsM9Cir6h/oSQoP
uq2fHjFTPGXGCKAngnHWAax4ZUwpXOHk0Q5gX5zwhKCyCU/3y07ebTZWx8N3BC6QOF+jQJfPq7jH
aZd8VaYJdhS0B91qcAIBpXgBtssyMOsLR2l/MI6OEARkWv1Uw/LaybhfadJ6mIGgiBw9x1sm7VsG
FZwmkxS5FduoncFF0lcJ8pY3t64PZAO+YxopqRhdu4SHo0dtFmumywuxyQTRIvcas5zpuUDyUu3p
FH62hDgSh5YTebX503jpUjdNe0R51E/7Clv6DkVH4e0BdQoNACdQTjGnoM77zU+p9tABNRy6SkqR
zjOzT1imB3FN8d6KBHhC6lLGeAjUdwxdHcRYgvWDbL35tobb3MhbR5OHvVSOmGIScuCHaWfLJFdk
viutMwc1937eb5WwNy1gJvMyBqufpbS5N3NmerqClDW+K3oS+fY9kSeV1k3xBef16NA8lHse3JUw
vDPk7sG2bp3MMEnUHFbQ7cNuXv/OAEImJSpFJi+G0A03CPdy6klX1PPxAyHkxSk5OeB9mbwP9Z/K
v3DsiZVraFOfIsH+S7KQm2nwId09nBFOLH6DxtMTLQ/hv8Ub6uppUN9evEAHEwxareloRd3ebSHM
s5Jmm5F0FM0PQsAxBKahkxQ9vis2NSiI09pk/ohRKslKQZ6QFku/e7Cm9hmxRUHITNR97x6YVYH5
vqdF4ALd7n9VQ547c1QBY1Tuc4f6uxVwz0LMqNOl3igrj0leboByh6uUamdrMjqQRbOe5MueeCMY
MbYp6wNYIVmAAQPoIYHvD3dZ1jVPXl4cGbaKGfwzPhLN93ZjfGl7lEvLpShqhNbWT6KIK8ivcaJv
IXQcuB2ci/twYnSNIa1VUgbRj4jDwkYjbaTVJNk+J6BQ1qWAcQ3ZWYcZ4A8B6IM2fqBxCD5o11hr
wA/PDp5CfB+SJUtTbac2QKbqLihw3chsSl3DwLpeS3/Y05ZFEDhlfLd3ymQ8FGzMf6XxAXNzHt8V
1ipudlaCJ92EvzEpNv2yOfZDMEmoE36GNT7c/4gWuwyy5QbQ9gSghVehU5B5BGQmuglEhxcer45G
Hi1WQtZKB3G5sMpn1KHnCfTS6WvO8ipqV6rRamljse5+Zl9GMT0790zCgOfhcoRAQdG6zoJlSZKB
jPWdw6/ZZM40BKudKRKvEohH3WjaxDkWM3pwkE/rf2bo82nbVmZL0RUIUgRrYa+bxe1Gzx6CUnVE
wi7bBDdvKJ82/1B9GQn4EDXMVoYoDbv6oGrg+pHAJl0qlCEiVELYnhctCMGsExwbaTqyg7ZKhlEX
S7DwkP5WNLvZfX5meJa/y1fhNl6bbKsRoAtIBklpHqb9OnRCTEbkbvy8tFd3L5NoO0Lp9W0BJfwn
zokeAoUoIeBbb8mcs8+1uZGV+ZtjuSMv9wMvMJ1AiJ3jvIq6PpewZKhB1PYDVjq0BL0isl1Jefuy
NHwWrwbxbZH+Jar+0BWZTEvoJknx/58ctaTwB6o6d51CHoXSMV82NG0L8NhXxKgq63yDSItq1kWt
RGRCwRKgVcLMk0MDsTZK/67btpnh8kF2rfMXi6Gb+L3L/L8HpDO45n2IsAf9dguUfNoUjfSbxFrf
aSM5UkS2Q2QkavB/Y/YB1OgpDij4o7W0eoSz9XmqZE1qySv4iqLAuAY3aQU0ePJvKuApPh9+/Qt1
RqQeYFkRThtsjyYUSYi/jm9j3PGMEU6n/Rds78FEhcWhcOW5MAPirBT3Fv69JTjPjLUjPAx6MUoi
x4kKH7i+VY1ubHGQYzsXV1Ga8pPuNY8ykzxwFzbxOS+nG3e8RxzzV2I50OYrW+t6W2P6mVHm3BgD
/RikgDrP/iq7orZWN5fLQ3pLt3eiF8sl+XpwYFnykrtYHfBmuc6e2j4e6GcR2EvDNHNkVyQfK8kJ
GWrQoXCeCkQKI2m+5lCC8tQ7ntojVAXAWYwouMm4zq7FEXp+GolmM5Fa2zNp+NFE3SPbUn6dUtBR
FrRKh8jHnix4HLEcJIRdP+YXtNNcFtr4V6vmORde3tXjOatAJTPtq2K9ro0OnUAwZX1qmIjjh0LO
QhPyN1eil7Y9ps8ZjwwbROoI2u7/oGqBGrfpBR7bJffks5EkKLbsC9XCcs7jUdfQwxlusY5pfbug
47pFCTwnCjTzXP43BDEloUeDk2w6LLTSkPP66ujnQqRwxm3YN4X2JOL4ekaYib/ALodjuxepco7s
aC6JGWrP4JNHXy7ztNbyGbTRLVTHOIE49CVgRUcuf9gK9NCwKMVUyRhAjoBOvd54oKuEQUMWEn+6
vD16m1XlWb6/mRMAocfG1xYe4mBsnLaUygCsv4awcEsSt91zBlzXTNQHfDBT6sJQOwbn2jRvBDii
K6SGbIg0TOaVgqCYsF7VfkMvRS1ImMu80annhVlFr7GeifVQ+cW1/1x3nKXbtdmoO5uQWnkw+Lmn
rTsY0moIQ2jNoMmfHXgGyaRxqshGuDCcbimD1ApZXnAjPPYB6qvWkSQXaaBPxCMDY+l+ALQyM+GJ
1YE37Qn78ZmiD/m4NHo5wbITtFHprvNOQeWHGoaj7gVKtwqaJWZ5Iow8gYetG0uiiDwT2g+xRYX0
sq2U8IOH4RSkp7l6W2bzhFnyeKncRdZRaLe8FnEGTmbhWd2rLlj+d3OrFqXC9whmoER6g2LFDsur
H4X4+qezlmvFYon1ccd2p1YePwQIf2+4Xrbh4na3gVjmnLvhPiHM30SMC4ha71RzuE2c5Jw+svzj
OUtbnkztgbc3JASQOeP8BZxVc44rYkia0pR+3NyHtkVUjZFaYFEO5cX1H/9XC/FdtlN8KVMJ8oxI
A3K1+N9lSHTEOpBCOgl789jwIc1ZGAoh4z3BW8KNUNHIALEh35tGDShbJuMEpyiTNw8m+QBa2n1z
ML5LwAyxseMxZstsQwmjPN6yN4QujUV8E/gQASkpsIF+lpLlgRepTDLTrlbMgWbWjWsX6U6x96OL
Lmhw2mY2iyLH3wSjh9BSXf5UEz1sTW2eKVX9yrLuC2PWGvcHVEhjfNGYoitfHmambz5D+FnsjeAV
AzZeCIk4QUO04k1D+JLLKGLfPLh7uXqrykCfsTPJdrKRWpES1+uT+LnzIOI5l4joG1CsbYN5WUEF
iMplk0XM2BSLyYIoXO3WjLH9D+xxDV2IRTT1a0ObGHdHd71U6WtTbLxh2TCbMbFkP6It/CQya6ml
QLlzv4JhZNI/42TPlp1cYj2oiXwT/WHcYGbSa/NRY9zhwgqNExR8ajGJd6iLw51lz0ZPoYKwLf/3
jCxPMPPG0Hn6S1ka5qYOwx8T8BYAIDtf0MMR49VR5LQbrpKSPVNU5DO8lSXT+E2KnlDMfA9nRE+6
YDLqV1alHbYRVUajCMoOjfCX5am+G5PPqk+Ew4tbt5/9OqgHnLgjWo5ZmrX30UesgYMiJ2/BP8t9
84HMn0RNTqVbYjeUQycKZxBfkOftGi5dwJ1+64WmWuUoQJlKUwSK7DiGXn7sK9DUSxqs7JiHVpia
ZnKesF3jfm34XJezeNoz1Qy+VkdD15Ut0pzZFULIYjSpxVhMKa7M4whrs9EjbA5aGR1J+AcTqAaG
Vl5+fvVDE5ArXc9/MrjnyiPl0N/P42/noUkoynQasWIHnK+mcpPwrPNMyUxOSnjM7yz35c+dwxAE
9qdaxGALeCCKusGm7ftGJjQ1UCthoXcOIFSPLWQN+pbpBjBi4ON+O6jgqnAGWcGmRcxPrgaNgVm7
tFfciBEH5qwgJ0AGtHXL4Cg0GCybnscS41miajEn/GC1YcMSlhTCO2s4RyA5AYHeinraWM0zySAO
XQVdeJZ9GWDRRuro55y9hvfah/4z+9LK4JFQr3jMdoG0APkxkmS5R5uypYXecMh6AjSGqDISV66O
1llKnDZJN10MkPlA8STat1ZH9A0PG7LdM5jh9AHgD3uUKrHSDnZFHyMId4tYApHlTOj5bLpE+QaW
v39467zcG8cK1ejEbo/G9QkmHDTqe2mG0vXlgjPp7WDxvmyl4e9NfC5L2CW/cjHBykEEk5PxYdoN
b2W08pRd0l4Eb/J8N/hC5sVqZmciC0omQHEcOPBI/tBIImZOhyWiIc7XysWvbYylLVNR0DnYx8pv
yMkac4Tp7THTL7jGiMG8nefZh/fuD22iteemkDQLSgyUl3czGsYBSD+RjD/IeLQCGYIZ5N1ALuGu
bhwpmDLNORWdmr67KG7kF9a3oNZLE4KluqAUpDJ6X8H7vmStechrydGh61+JhWfRc+E73nhZMSWK
no+qKH1sKQp0gJmymb5klfDwRUxEmp1Lwgqa5G8SWBysJwBS8LznPgd8zka2gjN8MKovsp5YIQei
qVDqCnQjZiueGL42d4rTV3dOyhUWKSDOUQ0uAcMzXR3CFlGmSMe96dOevGN4IenQtOiCmUr6pfzd
11s+8sNPq6ikhV8wL8+gKVEw5fOMKaHDdd6M/jtWlbYx+04b4I5BCxBGm5DHIckCKOBiEldyaJyJ
Ua8+M8kjWtRQrDIRXzi3hlxtRrJkfffMTNg8IlcPxqnJ54Pzn2EHy4I1ZY4JEOJUg0Pca5Af7nUy
41/jFhjv5t/vgSO58fFJ9kkHus5LkLtknbxZmM+72i+w3h8mhNPWRPYedFEq23Y4VxrD3WQ1G12O
AuStgwlswEGlOL0ac1hfqIGpJJtAnxstEi8zOnEfQexeXnGY0W6MS4LitrJCC3cALSHR3hNPsovu
fBzWMcNSMaXG5tbWeZ3xrlHgEfHcEWQw+4tK+VTHezeWnVvMEaeOq0XNBNGlN9P2/2I5meApoCVQ
Ygf6HbqeQMpzQOyAV5/fclLN3calm0YgerX6LFd9K114FQ/z4ix7LVTM997QqlUF+QPM+6neVVBO
Hfbotq0h5r5v/FRi7e3r3lsD93qzHOL/7M5edZjTnZBlG3eBc+JL8clSviSnFPL1N47/n/S1jO+b
rB/7RtHSM/G9ZKEWfQjjRxihhyk0lVq6d+IV/hWPeHepkNlRf2CZfkTK4z6aypXg6psBpNjjoa6W
pVnjYAnhAsDhhO9tcak5NBUmjL49UXXVEjtVJN1iyY0XtGrSYV+mOSUuciW8dfzdlUrt6Epa8jJB
aDdjZtAl9vanhqWyTtFhcx1FrfcVGefvp2ui5E7eTcH1OCe0fnMGKAx9OGsZGk3snk0VpaVelO7b
ZDVVocjYCSuMyUp1EOs97tIqB+OcD7kqJiVP42RxVjgwIUbX+eS/ZEjsnYhNu8oAXa6QFosxLUBy
XFpODfa5yc7nfx6n7CHBdHugMGk30pqVLH9Fw4CF8ucUDIMkg8Zq7+6IYZqph8/3zh0bmMObm8/W
784PXQc0BCILMud9F9vL2wb/II6nctfUS9POYYusM+Sm51FEMYuoVSivt3qK5jEuowDOTaGsb+vJ
C0xOyi4KQkGTaiMM/jK/SqHo7C3S97jPreEgaAA6ezlN+nnDAvnlSRgwMuPryOzZDBeJftjPRRM7
C2ouVe/NCmA/F59mlWk2zmzfknx4xlE06GRcF/DWL0hFWcVMOS+HWt8TyQAmDUFyQim9Z7pLZn/d
Iaw6zRaRN600+/hcFjWJm5hSjplfnvaICrKY0ZAmaBljV3basW24raWoGPszPaep+p+vwAQfCxXe
EHwJ16fOgCN5eFvKeHoH3cpnNJmNkQqUXJqplJItIn1P6e66Y70/bE+XsAHjLzjKneg3sN/ul60y
tSXWaY1L64dkFJK6jrNyXIUidCNNq2bnq0MFy0oK62l47aulwFKeL45qO6NEWgYID+aBC1BI1igM
UMdw1MAkD4KAnfOuQYw5InNniyjD8yS9xDAAV+/Sf9+U86Izo2/u9BX1eRna/OmdawVuuSdGZn1n
sONKNUeBdhOki61+rvTAo2Yq94UkALR+3ABLBjxiwL/htg8fWf3JlHqD7LestoToaQK6FYj86UF/
LoF8QfzLrW1d5I2RM7QICobkm/5jh2IPFxgDer9FMHiiqaTURegZEzve19ODJva5NSxbH6zcGK+A
0LB94yFr84QZIoLsMPQ+h5AkdYVcDutBGf9F9dsDff5NY8w5mZr5CMZ4uTHhLoCayjfxs3OvDHaS
YZjVlWe98qpRcLALHIesVfjm9SDIxdzR2WOzdKzg7OvzL1PnjDzXMRnEhNIzJWCcLikXQr363QPA
dViQc5MLA8zr5brln2V/t0YXUm6FuW4CPngKo66bnNwlW80VrYDZPwulWz5RznMTG8QeCZRgXj4Y
09Npo+S5Jzr8RALIdiNu1qqIiQfhZXKHOO1tXO6f9WIeR4r/NmsxSlhO4n5IdANphQW1PuW7qlbX
XcG+2/xcOU0Rk7ss9Lenj0jB7/LsnWyWq0IkkVsY1HfUNGkOuUpAefRtCF1pJjXRU07vNho0aJyg
gxUa0aQnEWGWfWp3u0f2tuAx85NTHY1XZzNSouWzDw/ejWsNhvCGja2BDy2RQiVyhzXozCG8vtmL
qHC7VLYQM6AWfwsfJALc9wyyQamjPUreWnq0JoUSuv7ZnJHuUEUZFw3MWiLJCiUf4C/ZNuiimrLV
cIAFan/md2mlFzuVYs1WO6gh9F79RoGE5TjcW8jnXSEvusRToIx3GX1/pxR4tvfHKgm9RXlFuz8H
8QzZMVSxwz64+0Hx2aYvGugtZVrTGXzjyJ2hDbB6OdjRZpvVCYWYi6V6E7rwq8u6SN7QQVR6R81u
hZpoBuql6S6+x7I/JHXs2burvnlsdTbDgQHPWyXTbI7ltPwdVIXsCgzi2YCZ3j/hriT6Lcae6K2h
Geo/db4QtW+6YfKDFTdeCja6yfCTt50Q1BXChr62CXQ0zmGEtYgLBc9XqZU++ZdvWCqgHqrIIswv
wRxYYLNslB0nfY8DyBvU6A5wRUDXqKZJfd3UqiVOW8Sm2x8RappzagBNHFFtWkYAFvlFKTX3hcr4
5PCqdTGHSg6QEvGm5wCm/ELMDCv2Ig04wmPXXzCw6J2ehz2/BLkVbH7s+hp+ffFIzyoUoc/L82ey
/2ffpgGaLsNB5e3NOgpNMM0dmIRGVHw1d6J1LDz2SlFaX0SevTYSGrsUHGdrMZPe9Te+h4MNBbNM
B4grsoIalvqmaoBKskBuVJbAB+LyKuqx1vWSf/skiuVS7SXeGquw3c1JhEOpAYRD2wmdhspEqw2n
dDRfI5c88JiDWuDs8TZCbk5g0WuG74TzbROHe8BGsLRUr9KvLecO/wioEo+xDYVxr2EXNblFVMgc
ngDerMSJsBCY+tUfTJNGeaZNCCVD+vyqH1DEF4fNxaWlEIs00WJbPMXMJvGK1PtEWQoOQariDrqh
DGeUAoDfDy6btV4oVRbLBj56QtdgH+o2JJ5GQ+PONvsK6wDSxQ3II7WHsao0eUDFzz3UltIKY+Rj
r9K3EFY9zG576LXRFasEAtAaLmrW/MehbeX4dsskHSBYxEws1GZjhnRILTyWoW8LBGOmq4tcpeqh
NNLSg5L0c21HdpkLWOpUuErey0Q7uYDBWN/K9zRqBgoUIe+g0uVCVhTIxQ7mX8sgYUZk+D82uxP7
sz/nfPAHK9wiFVOPQ60QDOeScP/pNyQt8O7O7RmPB74XawYImb8A6A3YqaqJidATRfBlfE60XYVv
bGu7j4FrVBWSUjZS7Uh2LC5mDKUP9csDHTjtPwz0+PygRwAkWvOe4ZtS5bKPC1oJURn8qZJin8tr
mgvQ/jNDiJUEDU0yB13OHov2XHmd9yC8NWY2Sm9CsmznoiI/KGc4WdbwtB8z2gR+VQN4ga+Np4qa
B117iowneTR+FnQDyy3RXVkTI3El2Bru1wvXR8SRQxXcmKLvyfnlw4GvxdigyMyiYGW5MCyfObk4
p136lTE3m8eiQsuHuEUxGo+R7irztmDWWNlH8+qaK1kNUdsHwCHJKIkh41mIG3UWxgsjq3wbSeIa
FkJkthmA5YPSiXWSY0MKyvojfNwPBrFdbMLGJ3HfdW03jpht92qMofS7MH7SiYYdDCQjoyZdo3/2
xoxAXXcuVJ8I/JhLkK/oRTW+dqcA0gUcT9AI5uQSTscEb087U3SzhvoQdR7BIZvuaudIPeQl9Enw
4gr8rPc+3I/knIrrj8UyxnPWUqlSZGTouYvthy/8hTxoY5GkpPpZ126wCBh2ZLFz/XHgraoT1Ce2
Y5rUm8WdUPlIK8OAiERkmShwzyDzhB2BZCLvCJhcxaJFGdTG9WIKQDHHoyfLZBLb7CSnaBXzO4V/
m+sWP/UMvaPdvSyuHFU8GhDD+siB4eoLJraiqjAUWSQ1berxQM8joBmrIeq5T7r8PUJs7J5xeSjx
b1MiCKMu0s8qc2hkaSOUe8bR6/1AJLB/5H53CYSKk53F45qJ914sn7QZn04/SrM8QyK8j3dxM5FY
4QgdrQr0jspAHSLWwDa3We81dUWh331hMPYXTHHYnFOK9xU45Lf65y7ZWRV5P9nvbjFQrOOuJtdk
Sg/LjWWQ/rsy0jDHEtTraRJuutO7j8JVg9J0KdJzRW96D2NnkHqrAbt7o63g3u1DSa3UbBQUyBvW
Y2NPHm/8GOLvv1z3NS0G2dRRORqUyg3rlWdRjIv2KAeZVNj6JItMjKEGmD8zBwuw96SoQw438skp
VEuU26AWjn0qopi4F/+HhAseerA1nYUyIvZ6HUGWCtAVkUx02zCxI5Ib04iG8Zg6ChJXDcV8PdC9
Dbn3ZK14dTMBfXX3PvHmAMArFQnq1OwrGHbHoiV96stoloIi9csIfO98MwpFXAE5qoS2ir4GtOxv
iVCXE7ySLdjccBJrYad1VCmxTjlkgUcKty/ag2YHDxCrSxX5IlaJ8hnRdlJvWboKIdE5imi6KoPe
/PFUOswbCkbvkbqJ8XFuIUFFH2SAlsxiaOS57obSVPvfl8q1eQMulOVwjxt0xhn55CWgRHtiuaK0
Ts/XSxXRE6mPEf7vVZSNQWYphqDK2v3ISw75sXGW8EB81mCplf74CsefZ2pBYItBRhOgOUE58Hme
CMyPg3cWpAsxNM1O9A5bar1g2pnmT0XyueLwjcl7Z+tDlLUwZ/00r5nzch4a7BUY032grXEwE4H6
tO8QUiHO6XnqOV3A9vJO8ewLk1HmmcOX85JdrfDIiM+O/WuzYHRWCkHd/e2+BdKfWDzMmbb4PGGY
Fwq5NDriB1t8HESmhsk5ni/9IkOdfBQAYgWD7z2cWyT1VxLL1jCGgIj9+NIYG8vH4SjiP5M4vQEk
Xk60IJqJdSP3S9nAXKQXxoanhXQ65OvBVMRnNJj2E568ZVd0qT1JBZ0l1wYhY4r4spHIBOD7vT09
jd5N7YYgvlWYfT+7vlsCN1O9Y9GLn6d9tNT33sl1uomf+PjKbEDAhQAZr+076y7LL6Ne6GIrnQiy
7cZ0CC7UoLemGEE6Dx7zPX7jtsF3wpsidEGiLWmW3GPMHkV42A6P6kPtU1Q6dB19UsAkXyzEFyuN
V9IeWYFkJbNCBb4tq7+K01+7V6j4E+b5IKzpk0CmkRL9ZsA5dntZeaMr3Usb1L89MygXU1kkbvwY
Mh/rnyjCUr6/dscDwwetfwF4vCkGzGjV1aaga0Fjl5Y0FNVGs3hw/pwsCQhLOxeai9xLs9wvYgsM
BssuoFaHu9W07GiQbx9AKoIp6DSW3Isdqw3LckgYVRgm4G19sVSvHa4CE57bQS9k+vQasAtkAaXr
B+wOWN4g2p8JVjg57v6wV/OH4IkKyeqJd8+omLz3PNDqw7Yov5wqM+kDmjVdbtpeA8h8Rpor7REs
5w4eZ7PR/LVMW8bb/Hu+A9Z0w3ngXfpEv0XW8+al9vLOvG7Ey4JyMWuNk/TogJMRMs/8RlAeH3QM
81mORbQHGhZASydWiI9ReuNhc2zCZYMqW6YLy14qXaTnXwsSfbCDlDVyWYAAqWAnR4/iw19YtIsA
XYY3/JjpIye4Na+xAiV+qUWXHqA+Y9GSwDGa00VluRZFRg1uwPHqA4pKBlSOCL4fkp27AjNLKpIU
2G5HI6OpJsPwJpQQFoxSwvXHGPnL7+uM9KCRcaYIpMz2Wld8oKP6qLCbFjmdBv5Q9mkW3ninNDLF
mTx3FQat3VhS3zhAQB324WbyXY1PsR83+XFxG24dKpfuvZjwfb068mltaQG+pmhblq8clXfcOFuL
K3H5Wy88LCd7ayS3h1rEXc08x/Nzk58doHjYgb5BCbzB+DVZrUKDQEPZw1xdoe8TkVutYG88tLFK
22W33OKI72z5wRWAuUaMfaPaSzsjDKNC4tCK28mRY+O2chCe3ve/nHbZkmEBwap0hphpIXmG18aO
tXi6td1uQXpPaiTkXu0XmvBdzMt3eY73GysreyoKGRkKw+w6gzkQm63zS+WU9LIPeeIVfhu+626H
zEEONsYaoYAavDHjYamfezm9RY9VFBlRCBGU9HqM4gK68F/5/CWRBxY8YUyS7R6JadTNMxJavsWV
M8G+tTS0ao5u97rEke2No72C+i9J23GTvkJZqMqMLCaE8EJTZaxnxQ2xsTXqDkhWqhjE38La7+C4
qb/L5S0NOKMsXh3rDd8AOiPpU703aL3QaTvx6ZXwQ59K1naVOKJ9SSXoQYrJJTR6Kqll5/LRew8I
I8iXOyiTpOYHa9HlOOtFJQPxbaRAnnJR8zlSlwaP6Fb6MZkgyCo3URdC3RXuLGIVVWTfzgVbpyeq
PKwSpc9/0KgMMfccWC7k/V+Q7hlTstrTxvxGK6Q8Gi/mWSdApR/xmbdi+eP+y27YpEXNiLYDMK9P
dRoUAS/lCPDbh0WF9Ql1Jzs/0D8Utge61B+A7y7iN/M4JO2b4O44Tv8tOD4u82qBf6QB2PXwZmLZ
dD/pSm6in9qZI/Mh4R6/SNWKnyA5evy7XkVUlT5oE5HR8pGAqyabDZKdZQ0A/kDDWmxEoy9i/U7n
FUJcExTY8nIRMu7WbTpmapkBhQrocyTmbnRMZxPHbZfqFNRUr4WbJg0nv9dHS8ExpPR58/frsBDV
mdV6KropLN+Q8XqIgKTRRYanIjqulWjYEJQU/e+L0TsOurxn99AB0suViM2jZ6tuwtp/o/tu02WU
MnuQ0D62FNk2WNRtz5OYHG0NSV9AYE3okyPK0n8id282GmuVZ7gB9kbtjxjEa59yB1TaUgTSHgXe
9s9ePngqmFWx5365yC3WvAJ01zCwK4vDKQvVHFLKMpjrj2MdzuOf5SsKdwP9BG/XibdJviafz3Gi
tN1tjwNSjwuEp7q13Jwcd5CZjqmr5J1sJ3aTtSwyuGlA+zE3Ch5wYIoppt9oWqhdPdfqjxZGZ8Oi
IUgErgEbD3L610LCj6T5hHQCOOE+yo1ncgF1eQu8uOsxtgEy5hY/zxOdyzrSQyhI3Z4j4uJslwF7
mMEtFemDTZ4Z4GSvGQofE0VdSML6pk0x19Vb1t2cUxMAqDSvos47XUqdiRZF4tFyD6vUQNQqCX+c
iRz/7DpZLqXXzFL4eZW3L6Xtn0IdT3rznpj3/HmbrT6ScXLqK9ebGhDXOufc+ovblaD0pqlHOOlb
MFKOC9VuWaOCOgyq71vokigbk3EMGorL22VFDKpdgw2Ntp6SuWreCQr+oKCffbvKdKmzBfpz8ZIE
C/GtdBgqglnTGr0SznM/h3UjSTqGLS0plJHiabQ/f4FW6na8sdJgBsJDEzMMaZmlVcV/OUfw7XRU
rd3dj0ScRSb/cAP2E6K1mNWdbILiXJdGD8d6W3sCLVypD1vpFlWAs2jU5MthR5/4Sgdz5rSoJs5G
Mxy+EChn9pEd8IBbMc9y7H3TDdNtzPxMR4WfatHHKvX9XxOdK+HnEXIZC76Rf1N9tbydjUOz4+RL
+d7Yc7KslPoEUWbCXftRSrLAI6WAe7V1nIa9IW4aD6YvcqYsFM1EB3PCU+S1HltHwLOzd2nqb/gf
L8atVM3k4SskmUxCEeXzX4zfclAoCwrX+LH87sonwfiIt9sbF6GzBLn8KiDsVrwq2X3uPBYgZjFf
22G0jWlQPMQKoFQIz3BPBAQEcvnDcxlmv7KzirevKQ7KRUHTqL/MmY+BbWG5OBLk1UsFrWF7qbAI
aSyxg6uFcx5uW7QogtJJeJ5WWizeOo5eY9u5Dwhbtm04LyHDZFWHE14ATvrlY40aN4LkW8NHsTuo
+wAeZxV+Fg2qOuLrXaWiXvFDWD6yxYqm8A1kcUQiX+lJ1scVRr/RDr74KHwmaXzO9v5H4RGDPqN5
M0rTDc1NWcshFZlo0j27QGvOcHIAqqyw7AvklSDJIDZ9GmG1dVtuBHYqTJT46S7qrJ3jfpcYfBaV
ZZN4R1ntKtKe1rT3ouvgQTbbr4LrJudUf761MP1FTi2q5WUviSkEteaA3ZCs6HMxx00NhNge9zUZ
3fD8otCUD4fxmbh49NOu0hEEsmLs9lMmj7LxME/PueeFg/AfCG65edhzo8Czie4cfZFV9sn32jwR
N9cJaffkneC9oCJJ0FoVHYp21d75ETyp00Mj8Nvr7ZWIumqGxIqBPKGXhhvhGPOV+rBAOR2egwvD
SqAP/11H0XXsw8NicFQRKIVmy9BusAHXGnejflc3fwwq6C2Izjlg89jHR3GqapyBKIgkgOqQ5wB0
3oc6e3kTpddhpYHsEISAcMjcNEN0fOjSfxVWOp4VnwCCdfK4bLIhWg5E3OmXbhsC13X1NO/CZ4rM
3mCbpj/wuWXZ3Gjidw4JVo6euUyRT4P1+b731HJXve9iQzXMpcEdIzMBxn0EdTmdz6hLeqarL+jO
cYEW/j5URHVs4Rcy4LVRi7YDQcZmdnPO+2rHnptavdOqzFDCB0LRLZOrQG3KtYVAj6Pt139q47iq
I2gW+4N0AufRnGYiukbvdminVx7tNDb/ah3O4kftPGbhUo+lH5R6uR0xkuZB/0yNQRAfhXLejJ09
c+qFpBYuBoc//NF8AatauPWcPVOf6CoEhTcbd0Qq/Rw302EwRa/Vi6OFWl6Vg+Otd9P2XoYuaOgR
TPPByptPMN9OVVlAW7eS70e2+jwzyOSgepRikzXtX/8hb3jAoq+rbyTGpEIva8I5CGkDOhtlxNIC
ie97TqGw6NxkvvmYpLPt6x3W/zuRquukoy7ozBwhpjFPuQUK41Y16l7YMlXfuRnNbREpHRf9U1sC
mNMOTFX3m5yn8yUb76yiIYzaaFNJAUXFCxyqA7jleRFolYdJpNZX8xdbs4jQL0T9/nzx8795iGDy
tduwbptVU++BR/1llOQfxYlN1MF7/U9Dlj6oTQ8AYmAgkTMXZqsN2khawygO3fklEZBflBGamibH
1enMVJxNO1JCAVqU2VvOCQOwOKSutj2qkHMC6CD3oeuzAptqv+TzGFK5yGEiXi0ig/U2aXhuli2e
v0tbZZ9WtZPiy0YmPJC8zFe2GLz8rLG6oAQzsREQGYioZynFMZCLF57IbLk3LM7VftpBJcVXq1Hf
jRFrTI8SfAFX0apa1GnfwToP824Gf5sKZvf0GhGjWeM+w+vSQOFlONg0J0wYA8GpNA7TNbleUoOk
40s6T8TBXHJKEyVvAd2WC71q1p5G2zNLSCLESPIvFlNZuFCp6b6VBScXM6hf4wZfkxYTMjx37nyH
YL9qKfb/5lwmqNXD7AzuPDTcbLutQy3AP3fz1LbyguiYaaw6jwfiZdSw+zFSG+epqdwkhrh0zoaE
sZEUdKvjXzaeWfCecTyIF3xkGsYzRqJo3VAYaoDVYmAjsBDsEodOUVYx+/Djf0ji+8MulnmqWoIr
h0kqwLeBGZEUReQx7mMU5Cx2JB6j1G7n9AYO4KPdPxItPyttaDyo15A2CFkaeVLzfnfsQHmzIjtv
ow0xu6W4GKH/SmhxNpNr6vFrbZsmX0OPCMCW/uc/RXhzQ6hkTcCusqoCP40/byr99dS6NR0ctXBt
tAbxaHqNrBrD1iKsIn7kbXCJoAIH1XSihdh4Q9uIIeREJvXrn8Cree95o0/Zh9RdqOOTQOv7AkRc
LJ51N4HCGMA0wON1LspYx1M5MbQJ5QTRej3URNLuWOe6D8Z0xglf/R+PAXa5hQhbnLtgRZ/IAb4D
qI2EywLQGlrOuGkM4p+iT1FMpt441VbaVyt62cJjNi4nEWluBs8xSsG1DX1m8lBAvJozCNc4ZqfE
IFQYE5IkKvqUxg3hz+Ssv4mMW9oKhfw26/QF5ifmzR3dfZbl8u0GCLOSwrXtodP054YMQDXUIC0/
WEIcaujKlTJWVriAKYxmMlAdeNhQcRGKbNfDbqacabR6fCc0b3ZDbTvqWucJQzTRy6BlY2u0hqpe
qK1JExmJogHAaOFz2iTsojGE+mv8aopJjf/XTSZmKmhyIlgEqAIwSYYrKIzUtwOMQvpHGsdtanDl
LkANIQxUBbnFrAyUbEKp2yJcjuS5l/aYkFD4EAX9d/IcQzZXdl4qG4XY1oWVJYxmPiqERfOx6VoX
cfB3Uu5LYFH+YtkcPncmS7gHBn7ze8Cq4vjvboy6zb2WPWnD2VY3MH/pMXBYHVXBbWGalPTz0GVi
UQrJ7zGPrnE9JeLiI2v9cuTk5PbN+gMIQcVfLVPpeWr2Wo9jfrfFdgo8E+c/B0bhyuz0tFFRZKYa
mQvtmKh6zW6kDslPifY06SuGfhZXoyT1HXBJp12lTJezkLhLp3wAvS9iiTME1++JX2qQYSID30Xq
9yMeHRQr5UQ/YgCP3LWvgoklIV34fwd5LGXtE1lhShJWwfI+ljN0vTm5mM0rhhAA+wqq9vMUPgIo
ZkRxdWcv2+q067EsjZe2ng1dzwxO/fytFny+qiK24znEzkAHffIxc2kUzH7oRTOSQ9LcTLpnoTBt
aKbKw/1IXnt9Qa9i4UHY4Zd2XcpkfLy38BHPkzqcf9NoZTQvqtTyGVnnFD+j1SeO6U2JioiYesj1
YoZhgTq1X376bXTGllA7Sf/JuIAo57oDb1Ysdv2S96YAzIL79fjgZsxqD4sH9tAlYWk8WwZ6/lou
mBnQtNwT0tMwdItGYA3VGzwzG6mGLiD+JYPDNPhp5thOODA9X1GYXr+B94lQNWsaoBCASvR0EU2U
QeQkVr8eEIWYC2li4SkwrRWlWQn3lc/xbH30LWL+r5GIsJp+/IFxUa3NwIO9BGok0mlEqOKitpgR
/oWflmXsDERRUfzMQBOTXq6LCh3xtBaf22xMhoARS3VVA2kcGuT2EegFMJCglBsHdbgjg7IL8l+r
uiw94bwg8Amjv9IV97x9AQhEhyoG1e9qZnDEsy6kS06EFIbsE/1Vyj5WTa3cXjqH7QozHt6gw3Lx
PQ2K8r02h82IzQETNxTy25ok9eKn6vTbbXseQbYdueoDlJLVl2nxHjvdKCgDjfG5nxXEXuyZ2xyO
IQEoRxtZPRAUhyQCIJoePvFGhvI023gXo/geTZ8d3Axsxhz3t/Of95kZzapMDgZid09ZsflwOd0A
FYG4y5LLtWasDi4Kl5hcPM6fRZKt78WHLR5G+Qu2wEe28GWcVLAmB3Ur1cqZFvrv5IesIxnr7yzk
PjnAnoHX5mfsb8TyzUg7JU/uF94I4U5m1uUNTkNtgw94XuijP99O2pg4kJ3lDfGYAWfZYY/DKbQ6
tLVSoLfaMiXA7GNyTggkC4Ml9rQ5TROI+2pD7qKy2un/2hBwrOCSbDk3OAviJy0ceh6UCboGW/7C
qcLo3fqd471TJnlmTX3eA+rzf1u6RvMgv8WVGKjf+36oRjkDLmC+WYFYW00UaxZzmD3f7JC0rgvr
czlCUxuyX43euKabd4YDaeuOUyyeMsTu7V+dov0PCcbERJdeHdOTwweie3VUp+m6pfgVvCn7TJbb
DfwAxz6yFrqJjMW1Hpjemaai+mypPcGRJr3wRjvwUx1WDfw55akCp2c/Xk6Quls6UbEq6uvIfaFh
Tem2PFL+R+f77XI/h0lkx/cMXzmSvNTkgi5dX+3eRTlQCoxsbydTSHtg5+OEnIN4ZSBsai6lrRri
pSZjtEaeUnrst+n/fydQi+On/vaiRtns8PEa5pNUm0RkjlW/hZde1kn0DsWzUrVzjFpysiJEikby
EQOijH+FHk2DAaJqs4ztXUQLfPWmWDwMgSggAFioAnYviAqAEuLHBUH4dBOsddsk8Rzx/R74hz0O
IjJooE3e/TyXI52mLFVHtQCU7Obmjx0XxKAstjIBkPWAsR3HId5bbzQU1cs+sBt/6ofKujEy9Ahi
tsF/mqMWDCngIE475pEk2EjD4RmN7bqi1Z36hXYX30khXHU1zM5ZWaiENH7FMS8Az81/xdQCWDgg
tP2n4LwCc8lI4D2D6Pj0VpW6cScEnqIKxSdETsmYBUAO7u6hkAly41e0a+JMu6ncZg0hQcL6+Kgl
eTBv2/3hpddWYTyysVXVf8bAOF2R+s6R8EtRkgRye4ZmPgJCnZjfVyE1re/2vdVl0MuJNl43XEeC
E2bb/snXryg5uBPPE0i58pCogmj8wtuidhHFNr9E3aMl7Rim5hPBCStf5BxgbP14d9nEUecLBh0P
GN/c1OEZl8nVmgqkxeNvP8hei6vFbuvgKkxYN5IrZfvq6u7nHqzhArdyVEvGhADAMuvPMXHsM5GY
nXuCrgcXGlAz866Ri68f/QN6yIW4m67wFtd+sMjqJNsytID6o9tUWM8YkKfmz9uV5H6ISxB8aA7b
/VfR7rbdplic8CuCznqHSbGLGwQpN63hKzq1F4MZn/kEY6uWtTw2rKDWaYpzkAYXq9GLVWbhsgwH
bFFqhHISgZZVambJp41SDqZKEwndI3HOmbhQkq+1890jswfBtMmY8mV+QgmYvdBK4S1X9tVZ6/4j
ONsjE/TOMfeKOP2mKTFQRQaPEQsxJv6NhQazLR74QV+60pjL0IIdse9dxO7jLZ/Byx5v7eQKKrHA
thOn+4JYM4OfowUNILYFMLXS0NCSaMZfVhUPjnUeu0xILvMDTbfmB9znKA4YwtkqUK+JV6fcbagu
xsoGhoKZF6f1dXsywuBPVi87gGrNOWl9QNuRmSOsLk4nrrGSp4Ztj6gQxbXAi/FUxX9hJuwqTX5y
QRTPE5Lx0OEgobC/xWYZX+bOzQWh6wCPH6mrA49HvQuc+p45vGa5Ra4dgVeWezGo/DGeqY7mZWBs
Z6tYw6pWe91p7FhXCUBsoPPiC58yPV/H4z4Y/yVAutzo5NeQM5eOuEzr8Y/gUP1N7E0TAGw+BjkC
0ih6FNx5L3aAAL+B5XikufQ3MFzLA1GarYwiY3viX1nFdVMdbHMQaUHwLYTt4LOg/ZPUE0hu9JEt
gGfri5wcgxnkXjYZfHywF6oKe1ZkTMqjdxXaW62wcMx7ZV518QwFVrymzZO+eBEcIDpEcEcq5Rci
GO2SB3EVJPlEYmLtnGe93Qf4EcqOrDnU2qkoJ63FAkhisipXTIXQYBisaR9oOyxRS3w2ZbarCmqW
UbrDldOBaUxBDoKDhSUW2rqgGUoLaCb5oXEXuMn8DC2UvAVcWzaJCw+jpqfBiW2qf+tAF4c7yTVu
qcTuWOh6bE4uVapEMLSAozJTqtDjJdCYjmHjyKWBn0XvTmM7upg0l45uTblpyUjOjWtQJv/6BA2c
85f2LL4043L8l2+hwC2e98H3sdjKIyeVYbLD3KKpxAxnA5qShKxA4xIxekfNNLmeDyh3Zshc7+2c
kEFPpz3RAuC2GTcrpGDSAFje7fF6tj2g6L4OU8NBIbiixw2y7cX35aU/LxbwAywUrzz9ZCEudUXW
ocja4GUg/rNIeQloNBzehx5QevozGxb79qkROUizF/Npa8aiJkZVt0I3x1W7jy48UbnVQiorZZkc
BUFm3VR/gGKGEQE4pyFmu4U0aGHUQHgv1j73BqjsxriTzkk0SMQoCkQ6SAgDhL8xb8ntiW/6gdC0
KToRXnINSbd0DzgQf0b/HWAveXXiGPs38VKcGdYAmDea8wfUYLuDfSBuhdsoaaHPmxQ1nlvvz8Vm
KbNjoZ3b1VopIFLK0mUcjym2uCeD7CuKfL+IfhI8Z8g9wAMQHFeXbozbDJUaQ9u7mJ43qO3TREHH
AMNwo0BoDV5+femUA6oAIKQ9uD7al1ypO9EfPLrd7ECeC3mpjsju/fFlY17AemUAltRmBczlXnaL
FqR5usw2TWSCMC8bY7EEWMWYtcMkS6X9nSfWs1rrqd9iz/BBztwRwCkq+N5fVOHUV92ZL2093dj6
L9Ukx5HLm9H+5RDnlfT+Xp4OWsbYu+IHvjNV/NHD08etPPxzqIOqAuNcetQ/wkbvQcsc+ChdGDiI
6IONWHPpjEgOjyEsz6L33iiypTXt4vsiMBIjlCWl1kmXFgPmjZWiKL4+TOa6p61tDnoJTxT+XtLZ
FNzbuiKgNJYMWb1ePXp7D9Z3h2bQBFZzgd50ap3jVpYA3TySusGWkzC9wHHhWyMnBB34Ccwxe8qU
KJgLzs/PxMjAuXedocFTe151rGh4Nx5ms1C09vuW5y4ydrIKAERYDAdO4o1T+2ERPTIgUzuv+gAF
NXFW7KKfvNKabAzfugmB1fs9qI2rfJKE/PNhEMNCfbe2EloOUURTnEIvGypGuX9sppJAn4NroCfW
O/xENGLe3OtE8w4P51YViE2IYTe58rlcy2tLopD7y2xSqhOxJ2Gfg/YymUCrlooECJLY5z73nRS9
HFmJQLJFmkG34u6jsSH8LJTRSbHQiZXwJzZaWbMzFx0b6PQXcu5uwsRiJ5LT2QmI3qONMilpmSCA
58oFMdeq+6G7+owet5OmWIubpNH+Mcq7kvQEBOkqgQ2Z3NQVyJhG1ZCbLSCHJe/7kJRlVyJNfF5H
Hl0tlh0iZCNAdYXg8zM6MWrSjBHqrBHuGtcWigNSHVHyiJKq5x7027TrREq6wiUtwIR+DvvtlzMf
tY4dhCYbEB0ARnk/dWM1DZAJdEbk02S32s2S9oRH7R0GKEAN+BX9+MT5z/6pdXkQht2tTtej2Qzd
lVLFZD7fPw63OHuqPYcEREvC2aXCxO4anABs7S5OyOK32C9MiHbgGeKWjmMb6uKu1Gwrtq+auEWX
bOQU4Rggfavg3rdfDWpA24NPmpUMteDcTSklOIcngXvvoyAuXMgdruD2fy3t45v85buGwctQRqk1
5OekAwM2MkU2A9uV9hCL1ZEmGBNj0vyuA4z/Abaz8nvF1d6NAm3/9167+BL7y/a9rl23wDh/F5JV
Xwzb5NThcUpkgj4VEztfKhdbm9q2dDg0oCxU3VcOhh6GDRAKvDm8EaI/mYu5xZvNZU8lAJLPZ7xX
JMJUzpZQH/0/BUgngn2wD09r3Fy805saXrqgNT25X4YwyPvrVGwpA0SneulGaiqDDMclwJAiOPz2
EN6iFJyAdldYCT8bG/9VMCddhqLxS+w9WRBGh3RKZEmjFdOzWytRLTpVdI2HmUFgA5FOprQsYEyc
azBY/flKxLJ1aqj6EzKUmmEMZo2lNvHqTnNyDtkTarwvJXJ1x3SAwG/DeciuBY41bLhaL8VU2/Vs
p848IMF8ONrJsZJN+Fs7RKlgWmJYMVzpxEg4ITQYfBBu2ro4QDNkqGs09yVDFYQXogdJSIvet4S/
E0v7FEHWfx40ZbAWeRNbiaRLyBhIRpQrqAMRVeghG1tWKfcqBsSYWKb4u6F1Wlw+XmUKNPvHJ+v9
AFvAvoM2NcR2c6XwT/u83xuZ1LWoNxw8xHG4QNIuSoFV0g5aVbP/W7NhhoXgZCgmBgVcyZomwe0c
RjCwRBJuSw9jrzigeX4RW4THaV4wXQY3uGJhNAErkfeeaZb62ihkbmlcVEuN6uBVJnX3VNSOD2Tj
gZq5DmP5kbQOzL3wfiZWYvRtBhBH4QMW6PAbBQiTLjk7GW6MKB97vfIkozhpbtThWqMotDG6E4j2
KO1GELH/Wo6RWWqS7nYoplXQGO5MU2qjpCf5isCsF3VvSTC1SLTI+PbLyFanYaBrhPe/mkm1jbTm
jQKee0FQy0+VqSWemGxDjWpxHNFmdSLKSH4S93d9ffqFJt8vbs3LZL143k9xri8yUbIxryf/UJrl
cQFrTXmq08WOx1CWcpzeWA2CsHf28K4DHfdLoDbwHCUInCOHgs+lNEoxIQ4RtBI+q6BD5Q0NMKyP
8Y059HvX6At6iK6zN9Shwdi5Gx1OlIY8/NW4i27LW9kfUJp5QKJDtsPXqvhd48jaHSotODyL+6mK
6iqRNE6rqbTVbAdwgGnfFmzT6qHOtQ3RD5hL9kRmkonh/zAmWn8+AlqqpFfbrDS6zFqP9IbMc4T2
dmF7CuxUq5BejsBe+Vto1XD52O1g6i2TimF4MTiLG+vJTrKcetDLLB+Hujf5DUflvI2s6Gv5j4/z
4dT6K7I2MtKoH1k1lCP3GS9z2E9h4xw6EMGJSrbehoUWitIJHn1IuZc9GoNLpVFcf1sQsf25I8Ez
rA6qJfZe4b2dMvN+hWgN3jzhhZUhb8DdJxln4ihTBIvNL6v7UfeZ2oHgDPFS6Qg8NPnZigiDZO4l
2rKxJ1oU0ULgvi37XUDZa078TKoPvFBPQqS87EmeGY1zJbxF184vkA0IkxMZqlEtLkERi5nbQZpd
B783ulpXKBI2EFjVm9CAizRcnrxgqTrDF7HS3DulHt8UStQJNz17IynTcVM6dMUpcqIqujM+XtBc
pWqaxasxkNmascuJSQuOHKIqHe4XZpDvrCf34HuLJEmxNN8mHRh4GgatlVkHM0SEyvaoapmo5jzg
M6es6s7X09VQ6G5d4etr5/ZTYSnt7sJS2RwTPb2mbg0kBpHIUl61HoD730b9wIgJKetLY0uTyFWu
a5mXUCiXAUNVV1oPrxgyO/nld8nP9/BmYBUbufDE5FYNFk/+/L1HdHLv/1crxkY1SoPZndM9tbWQ
L3r7rScxhd5CJEjBgHWOA5GtKGGywBOYA6/o88HNuaDzckycuh8As7wuvnESJi1BgO2H9tLK0oPD
tA+bqDsQ771ZqjTgXiF05VDDcMJ3UX4Tot9/Ir11qIMjvrcKOe7H09OEnBKoJ0znPpR4OEvWhk8J
CdRcEOw99ZNmG1tARGuOlbpT1jyWgcM75S2qZQoPZDs+wLyqT1epXfMb5jMon7H8DnuddKgAJg+4
CRcgdhnQIUarT3PbBdAdMfFNsM1/ttsJ7dzAK1RJbL9ZnaxWD9MjO4CeZRfp8yzx4DEj4NSaZVKM
r4LJ/T9Ue2JFkPxxIha5F3LYSJwuCocjoFDQNrgEu5P+7/LzdrdoWchAAUdFI2QOMbBtCKNUeXUS
rlHPTqEuPGPuv0tUQZ9szr7VEvIB9tzdPFkzW8dufJj579UvfH2BTwjLFfyPYp8Gu3YhMoMO8PCM
GFn9c+OgLy267rqPB0yuN854LeiSxmdGa62CySexmJnMQF7TYyRD3qH9NR7+0UYneUJy+OFfT/hq
1z1bT44vnLRT9xTlOeN+01Ri06/JlU5b76pfCbuHyIzkNgRaLRq89MkgB8miXoUQhEfQU8LnUBBB
4s+386i2cTvDiPSDzXCfPhNq515OvERp99alyBD06JYTiYPjnMMVVr9EnnOmhsPSlGaG69utUR7G
Yove1DSFv/G4oeCHxNZ0ay9XRUSl9UWQhHqdPG/V/JTvKkx/mbMYj40S+hZ/s9Tk3IZLla7l18J9
3A4LZDSFk5sdYtW7u5xxruTGNU1VzsNG5WPoIoi7STRi0hgI7LZ2GgO5B6ez+PjgJ9iuP83gJV/8
pNwwqpiVzwsog/vgR6h8F3SZ1Z2Cb/3meF3sSAoMRjyCK6KRu+EUB2QoH5dRwhgvKHhdJF6IsIu5
3NMhYeKfm+MU+fiGTX9wYxIs4xnFgj8xmiDuVEyIS+HWnyy2BcCPXY7ZlcAqRwfx//wREWW5iiH5
X1vPjJO6ERlircNCqL6f6zyScnO7kY+dZ2jM56DXJFAHJws3nte+6+QU8Ch8+kxn2FYXnZ8Dzk6H
N1N5LbEy1vGrUlrMFIKdw+MGLlpsHVXCaD5Z3ioPa28gWw0qUH2P2flRIoGkxCjcHZ1Gu2QlTUPA
cJRgU1u4MLcbSFDeda86yBtSl7Ybz4E7S+w2A/fxticamIM/DaByurM9H6yzgru71ztCa2n7zg0g
j4dRcbSR8H1PiDuP2+rKDnm+FcE8aeP93eFr4qEhdZiNqMaHP1V9REHXYGgR/De402iykCfctp+E
wCMB7auCr4JSZnBfYPBpLyoKlNCQkLbtw232P8XWd5KZ7eIYSu1p0On+5lyFEIXozrvpz5LL9kEw
gV7FVwhZJILct0M4evVhIGElPCnf892PqjsRDsPIDqwWaWnFSLZQ8d9DgOcTHQsj1MT3NlIqY4Mc
2/+K7NlQFMx6Id7iwdrbKHqY6+3XvpO0EtAMQJS8LfsfYFnu42uswn/D2pt+w4CZZnfH0TX0UW1a
3shmESzcdeE6wKwZBA1JA0dsUXS2ooT3JCq0mMEcZeU2vopEzqYYDkU2KSAiVvE4+Hb/C+t8r0XE
tQYFPeYp6Du/lVqEnKsdUQTcADD+8dbBovPgpJ7MUnptq44buiuvdkPlqeuHmK4GTC01lig/3KeW
L0SLkS3F6Eh0USPu5+kGtGmd/T1ZwtdS+DSXMSurLYK8tV+mi5P7afNYusF8m7kAexfWkPYjCmEx
FA7Lku5lu4NvgH21iNMN6EosG5QPd8YOGHKfJ0HF3UAVoVWi0tX5eI3SsB0cA/quoDbEo4gKUtcN
W/ZSg3RtKgBxkaj/9aFewBiQgM5xaenHlojwCmZTFyQ1TS5sq42Q4pNPUhijRSUNmJGT9V72KJ6U
jQDr+ONgIXWmhcypu69F9rncmWFBrWKrLAepOLLDBw3I89CEIIb8JnkKTWZzn9Ii2IE+VIVba5xU
/eNO0Hxqtw+xIuTaop1x177B7dXtYnERkL829bRK3DD5qMfBnbpy9fFfCwd0DP83eELkvR4nVkJ+
2cFfBfh1cuWh45dymTf8cqQYQ6E3NMsD5W6lriw6mJjTAdsRJZpD3CVVktEdJwZ1hf8Uhkb5LMCM
oW49wJL8JFGVlUpkjEfumpCk4SvQy87v4IsrRa2BLqkpuHo98tmA8Owdt4bgM/qgzzXgp6SnlCoV
5KsllZkQWAnXt/gmeejUzHkX0gYOVMXCVBoY81vgIkmJvQK8scY3YPUOKdCIld9YPzmfPnm6WfFh
Oix4yapqaHYc8v7DsC2OP/la/HJobixaeVzHzCBexGGzKlxhRePfT4hzvks2E5AN5mSD0bozVU/b
pOXYS6u1HHtDsL8O+yxVU4L3HDh6bW3CZclgv9OxcWX1o0pr6xvI1TrR0YvpxqaV05CnRkJewlhQ
DEriodxmyfQvbY+2b1v72K70dXo4LOg0nFe5FugcX3/zse4RAUpnMRseAOcb8vbanJuhAdFHXvZ9
Ar1He5QhqX1raUjKhbIu+2bnryG1LJ73RjXZEdpc0lNuRKCjaBbrWWiq6/cNhNGkv6wjBKJqG3D5
BFBbb4vNayINCWIjfxWX6jszE9Z/47kSfjItLgfmGamfUv+uwgyVbWeVfWec6sgmD2/H4b1PBRz6
GnnjAe8o90NKXFrdA7tOSUXwLmjcc1jDGLU6LIQRijMUEMAKt7Zd+B4rMnWq9gp9qZ6jeqFFENMN
tLoRwTBZoSJpgkB3iuOSFdLtLagkV7tbj81+x+ZYW+hoOvU/zI0g8MbVFZiXptfF5hALdua60jc0
jfaBPrv6aIJFrgbveLifXfbOLxJL1V3Sp/gBoAEBlO1miz+Rfyo4Lg9h5L9xmcYtcMBpC9UKqv2n
2dKFvMEy0quNT5dTXWLvdpoHShaJtsuaSVy1zP3dweOB8EWRlVfG7kP7v6G+yDygZpqhHGEInI8x
+Xnw6/n+64AaOrhgaIaQbpkjLG2QgSmqQJtuHJ5zWsYhFATQG0+rnPB7bbACs2Pg+tTZZI3SfqaQ
Ew4tQlM336o8gwSh1sgX98OSFNhWd00WlefSS+mLPrxxI63O0PJB8nlAG9At9r9HrHvZtaEUVBxC
/R9umqpV8oNCJpPNsNrfn3PUu+rL6GCmxNo6H2zLbscty15h1au4GlLzo9HBd+OPIiBx5nNtDPhG
9M/3sYeHh7URBVPxmsHRdK6zx3zuJi4LAJ33j44XQ8HwYR2uzjrb2YHF9k2tEi1REmlQtv1AU7s7
lMk+zNenrH8AjW3Yw3+Ig2Y2BvooKcGT6G3aMhW9mGrmosxtkyhQUO3djcjRfQlVULUhsxhv8Fvt
9FcGzE3JZI6/R0EGgtisFklXAUR1ZJWpDgk8yl8ld67ejtJ+uC3ZIPZuAFjgz5hvO4T+0N2OKcbF
gaj1OcMfPPlN4v3WiUdYkcTkgWWz7A9xcefDcHvBnJ+J0B9rslcU+Wfpz5W6PxFCagGAVXeOhL/q
/LewQzJeTUQg1TKm2EhWTW2dQZQbrvNjHm5X3ghbdsqvokaF848HDHkl1w1YlOJYTPFZBgAI5co3
nWnGUzdCEV7T9A0DXAAUzvn9v8mBklrHT7rVqU53UWsfUONU+nF8Sm7KzEnyONA91//w2E71EumO
6eBeejYEXQ5N/rzyhheLwVT6BNDXzn7UIgJ3AgxRpPBIHzU0xmFfTr01lD628u+W+KF3+vezg/7j
04MH4fi4UAr6T5st55TTW0lPL6v9xQXkarcrb2LETUGDSDQOkASXN9O55kalu1DqRw+lkG6mcE+y
VtNUTW8eLbYm7BrtydMbzhDml8Hk4YSa2xGY19Uqivo0nDhpxLAihJhW2Zh2JI4hWwQvY1raW79S
I7qYpsmhsmLReUw+epfa3OLghgbyLRIhzgPBpBLTsLTXrYzPLRdJ3sOGbLTv4AVbHkxPUSxHJJ/0
9kjc/Q3G+ekh1Q9DMfLla8Aca+UtaUootPKuuP/4frEg3C2xQ0Xj078j4+zjF5txbDdenQUYdA9e
oRok5PUm97DRTjnJV7jhbFvbbZthmBGj4kkEHpkqrpeFAbwTaZRZyUUle6RtQ6Csv/aBiibxsYuQ
ImpeQ8HaMAp8z3o8D8XaMoH+pBBPDI1LfE37JiGlbon2z2GFyUr9FilVu3Z/vNWXsqXP0CCWrng0
dE2DhsI/1s68DFlK3sEBzuSwt9fzM1FlxhymuN3DJxzpYdgRvvIhAFv9VrO3AfKeEmrfVFprtYRF
4syRwcMdXpGRKO2qmm0Hn6dnuBxWzBeQLt0RHZxEAVWTU7nd4q+neoBzCe744148/blFKCGOxQrt
7Zk2D9jvDyDnSLX21gQ07UAcZiuN+V+viLlRj7daot8lZYbRFPPVwCOZghWoZmQ9A1OMG7vzQ7K4
GAkr5c6s/vqlVzKj7GeBfPdVTA+S3pzkwU3qidQeIzfFg44nzEZ6wlMEuSmLbX3mziHhI/gWdIDW
Xbd0UnSkYTKcmmfFCI57/37x4RTMp2VPGNkfx7xU99fCeNl/VwRdx0rz/O3p1TPJ3wj+Cmd/HSRm
eRGaloxgSQ9P8F3qXqAq1lXGYSo/93XI34XAOSJZ/v3S+wPA18M2rUJ7XxB3YKbWJv2sWqUm6Us4
x66GoLVB0K1FJPqEsGKkLCZ2zUVX+rciiMhFYAY2UgVLJyPUutuP3TZDBnUSpC0QESHCVkETVg3n
44VT5tXmDJHw/eSqolyyawkdVTKARDQHzFTrdkf4Lgej1AAcB3IO755yeQUwgMF9EA8AVGZf10KE
WAxuaQqQSJulAtsSgzFYh+XzV4J8FvCMstG/rBtB8w2G/amX+OPa80PAHJyVEBuCbrh7YWApAB5B
cBmSRh/g5mlrcNHV42c91CZ0ueOx5RG6rrpVG0tCjcLwEGyXQsq2B8VfeCIwqqEcySu9jNqJGNuM
rMjqovXmQUfH31XH/rLflq7WVXrsGPP6s9IrEtDi27nbieGCmlTD6ikTU7b5xWd7pG8Q0SOqZteB
/kUqCTmwfSxuPrWQ5WZtpQ3aFEVj3j7wcXyMtbbWKlaCyxwePPZnlw8ToA53R4RsZ/UPHoWVxvcg
FZiedpmGcMuqZl0g7UVLJP6Kk7MTdJQIA4p4MzgRtZRHKfhsNVdzk8IxMOR1wNgKoBl04DjSYsU9
xCZHjU4nNclpq+NJNQFKwSHoioVWi/v5lZQszJ5Tii26E5PSbFzU06c3lL42AzfVGZCeAZ5A7OJM
RZ0TzAMUv0cJOD+ZMRLjYR85Nxf/mmvIJBSuilcCVc3wLXMsFZYHugGXsr0hX4E8L1mr0fjsQUNQ
6sdBElG4hxzsXSGT+AywGRm0J3Tjalqgc5sz8rsBFfC2qn109V1IWefqjwGpq+RzVVrkrXMqLYSi
erXrvtHARRL1gYjFbJLIabTjGDOGGvXbLZkwa+3866/pioY69RjeK+yQy5EZLN5VUhYGW4I29TDa
8oqjGHwRC8r36ywRfwFOsLcRIJCo0H4uxiaK/mm8saG7jfWrS8yVTShGw8J4CIIc0NSlJ0g2IG23
yE16AHZR8e+68+l0tftV6M6atPtv0DovtpAcAHn/6zXy1XiZutyeTiB6MtMXPAkKzM0KA/ZKueJj
zMN8NUHdBZ6QPONdYeuIJNO0hXwnXyeqy2QiBkQgswgmESMYZn0v1S6IsPpcplNWz77aSMZQvAbe
cb+qQLXpdcA5PCl3Zg1zMBwacjUnEGZcFi42hySesn5cE9tEmbQHB5iCLEhb/zSBz0M6JdEgxK3m
yOebIoF28CjtMghVICFRhwLNhV6cYXtWQJFcrfLDNTV+ciZvLErS3pF4cDSfxWIfpkByZj8iRXkU
L6nPPp/6aFZx2s0DqdPdk2kPU2lXAAPo/gW/QM48eFpQ0q/YjMMzXA8gYNV0aSzPRY7TcnT/ARaL
KQxrbVjpowTTDIiRWJBRoE4LowpFhtf/AuXBNTqpPTGrNt+UfoXRa1Q35FvkOLRJzIGJfBY41j2q
zOkRnptXcCcZvkL7A+Wk8DHl5x5hNTGkLxeSS8aBWY4jaG7HXjoTiHBvllrBA6idT2hS4+BaoEbt
r+T7AEtZlduYNkR7oD+cKD5eKolmwPZ70yrzib5hXja/Xds4e57RmoMN+KgBbPez2TjONjkdWGf3
HqDarrUc30Ewv+OS5GF5rU4Ux7/4U0RUu5akRuSR/LNiIBpL65IiiPNERcZ+t4+iqylEVIN+9EKn
PZDQ/5lhCabwzm8UTF9SCkrCBLsxaQzVbL7I30gr4HSzHkNb/lDG8eduMpzUj1XbdKeDYOLas77E
yowkMfZEKZR0JG8v82v9pifFrHr2r9L01jJoFqtrclSko0Nyk8jbW4WOGGTptUr8xgNSvrTaHvY6
P0cddSXVeuQ/gdNotIYEJUSxqk9Tshrz8v5G3jwEdruxQLu8Jh7/L3ivZ0TcNSrWZioqwzZ1OQ0H
MkW3Reo1H/lcl/JP/u88AB5nxfVwWb0OMdNZQVRD7G4K2IdRTqZIwlpMy4KIpcWYEEivEaH3KuXg
YhxAAL6Y7fe/ux2TZKVfT4E5fpEQIt2VZWI16qhB9xWBwmYtPHlXTFAp6FvU+gwAsQH2eEit/d25
5OVrtVMoetssTzqaHNI1XhQFTXsq640SuDC1yTukD+4KEQlHVaDRsxx9j0UgWc1sIA7MUHtgERVJ
W8L7ySL2/M8nZ0dI4Q1aruhCeldhCHFKg5nV+LTOQ6GDZCJ+3JucDhMETNJnk1gOydKjAyikTOXu
+uh+T+uTu7QLe3dkv7EZtnJOws68Jcu5u+KCsWR/HKaL8UJ1Ad4QPCWhUaXKsN/d1Rj69RfpgE1F
Yz2Zu2aDScwgU7U6pKffALQv/c+u85UvK07dl803EVLdGc0mEmZvKZL7FIAEgYQ/ydOvGRFsJlkY
CwHK9j4Z46mQQtCrNKvFVlSzNiYwrsrFL9692rUJm2C7ZoxkqGgophRHAU/z+zAQJ2ukU1FV16ts
ln27TW2gRK3syHNhP1ChaALYlqsn3VqLCpwZrLWslcQSe/4jAliB/eH/IEfyOHZsVeavYbJ8o3gP
DhmPVSthhmsV3LEEeY+UEx6sOiJ1wk+MFu9MdXg/LJF1a/OuN1xKxOAzWlDUk40DsseohbuVLPZt
xb0FaXwhCgDgEmqDsT/gYxBcDMw42IlbEttOhHOXY0RlFPf3IQ/TAQHGP4DnaWyyUaxiIv+Vc9+C
Qin8kqSpN8P46zBOESFn7YsGs9ngABo+s+TknU0QhYjnN8pvRbOMhikiZSIS5x4jiJ9iBcR9ZUTD
AJiZ6mMFvdRamSaOMjXeXAPaoxNtqXuc5nMkJSYmjor7HgDTPUcM4+8ShDr2FPl3WcJ4GIBQYJXD
m2ln0OHHRtzFXoImfWwyxI8Pxf8gCPDkHOLFzegVDB32mkiAnf/LUlNIkhsFdYLVQLn0WjmDIyMs
z4OVqxX/e9bgTv3JI8qEmDhRgT0ZlxSGaVJMCKCu8/DWRbMAeWtvzE1ZorigDN0daOfb7CtSXzr2
nTNuLQLQEJGFcQLTyLmSPDSM2uTp6uX5GMGXgmHcwc0itI2r4Gv5d0rfednw6kh0IUEVEo0nFiic
FzGEvpw9kOocsgrodBaRExntkq3ZqY3lWkfOE/RwuAv+v9ojWCZj6I8+0p2BE2vZ763gVb1a6OIR
+Hdstl+ExRwi0WhXkPkPuYEXMmONuKQOZXEqsDPXuisaaW7c3T4aiunZItIv7MU4X1L+S5zaFKVH
8ZcyVmqaMOBazDKMHQ4iL+z3uMIp68H/GC/nyOmXrdc09RWGOUASvZkq+WGZl+Tl+25Pelu9FBux
oPSHIzCjJ7POJynG25zBfSyjFBHA7r7oHtTwSabIHya9oq7GQa37pCPbhe7fEAbAgGpMZ3BXs68L
6STt8lVTTkO/KzA5KU0i7rOlBdNbJdVLLq9mUlD4Z6NR0FvDyBQdZBrFZIi7MkuQdWb133UID7Au
CAfTx+EXQv2U+Dl9ImkLQ4qevx8WRGxNXTbd0Ke/hM2ZQeXFOQmK79vBnnqR5jOP/6lV4gdNtwDH
yiCWZoLie01GrGHSgqVvm6Vo6SkEV5/4suACZ/9QPbmECwgS7JTm4pQ+EzrMEek9G5TibNrcKG/J
IWugpLL2wdujFDPu6pLfJW33eG60/uSJAYj4gxMpCtz8hUEsFvVN3M6MMoVEg2tWSqlIkMqaUJgT
nYfoGbAJx9CgRD7APCIc4ZKPG/miETgFDzFHbERg7NlKI17oIvhzMtmLnefqKTkI30u9ONFVyee7
tVs2u5lxyGt3iMSDzJcpSrrervtFDYdcNlWQM6Hc5/CK0YsLv5sYbvg9LUKIDIH8WDM+brjMnFfd
/JoBt5MFoYw1ex3bp1IA8rYDA348CukarIwOaoS93tkP+PvzO/Q1XLzA2tgM6hZBv3qBSW4wGPDy
d2axUE/zqd8BQESDhGsytg8bCT1tAMkDPn+mnoVFqcakrRwAABWb98yUm91V+eETpPeeIK1ZIck3
snJWJRW22O9aHHZUuNVNTrPq0+/fwdzvxHNdRe8kvj7/UWsLZhSgaOAqrbnxWvMPFPWYNCoCgCqR
oF3VvfDflbjWhnUjCsvybn4Dh1X18KGiPR7MtWbeJzOVUV5y6a/faIO+SmfUoC/3QDKyWg/9sBDa
c57/vFHKsRPTksd4Bg8FVgi3MPBmdwEv/MtmbRIanZEQJoGMHlofQQ+qI5v4MvjqC3SJabRrwRen
R6HwR4NYHtsxbczdux3pfO3UHrh6J919G5J8p3BwcIiBAxPlNOyAGe9bGfYYXyFBoHqgaBLCnKLn
f4/XstPKh50udRM6GZ/N3Obc+O7lxO8aJb5gQ9jLgUGmfN0V+E6UwVBqss6eJD1FPq6V+mdSlBSB
ANLir0Tw6nZJOh5L4cg2grWWpLexjPjTLyR91fN/yAA2AGNPWEmdEw71CyRDkfxP9KnvdxhhSSLZ
cS28MGfS1EI0nNZp0vvo3wt2rJ6vqXCo0wGdTgRCMfz1WtQLI/kmdE80w/+gaNj79DbeDOSjlqru
/hyjj4n6p639Olvxm9oicyMLX1CFAyrQvwrxAU/V0Qrqynx/xwCw3zH1DBRX29FBirdS7JAGKpoV
zMiBP25+R8xkLeAZMgFvA+4FNGGOHPSvEJm6O8yPZh6Lu31ooW3EDQFX2NCigYpMP9sQYdpNKVr0
wXOu2mA+drBxkmh0eROQi8HG+pnrTuPo1eaih62CWV6pMHqZzPzkOsHjONiqGBo3n72nXQHEokmO
O7cWDQwHYBYpTLdbIGeZc2cSNK0vnL1W3IplEhDLjndNWhdFox5e9BwrRi9Xk1FVdH75Nbl1Jb+x
aS3hARv1Cmaq6hRXjfBHr22UNZkVYqOeCDfVhA5SjJIodHoYGlg2LhdeGVnT1SpJ697GAao8ksJU
9faFaQHzLvCuQ2zNAj6MNqq5TNyuqXwWfvxCWoC5S1SxWWtcXt6qJ05dKalw/Rav3gBeaqj/7NkZ
TVLXWXC+3fu4zMb9+V4p2LmSqBo1zUZbLZH/XTrnM8xU7lSaH8YEO+oj2Kfz7EkkGT7y8GmoUFMK
Pw7i+WfelNv1Z5uIky82t7KdAvcn+tmbPTHBEB8N4CEYWseO2r4KqHHr9GgBFpgS6vQUA7lknUfd
rV8byUWJo1c4xKPCEEqRg88b8JoqHeiwWpXByASnbPrPEZ5l8/cSgw7ZGVXBF81slQh4RWXRd3DG
bnrHCkE2jRCoTE5gCpNPzo45iZbbZWon1a1+2kexvwb3Rg0x5wmMdw3ZQYYZZsRDT1WL8ITLXDGe
hbU52OBw0EKd6LiRnLl7iL8HVWFd5uUG6bix6qsc7Ok9SgtZ0Z3nnfyU21BwYx3Vs/PX3+QnWdP3
u4OAlnrYOWy/PwzLIAEMv1OeI20rV2MPulVey3U7ADv9Bu6qcNHGKpHuXe7CGTy3UC5nWclZHcK5
6FZdhxY8ReY63X50bA+iS0xMeDt7PeosjxbzgpP/OCihxc9T0DCruy9kIioLE3omfoOTHdEszivu
ejonDoaJnGpebKi6UGsIBIvTjT0JzGPTC7QyXxiXjz2cHwnHNPmDNujY/lWTQYNcs+VI3c5YQpCB
/aukGcUx1nI9Y9UmEploPGM5dT538HhwCDE/bnttsvfEwDt18hlxMJndj+9vU5sI7H2Fz0glDfKb
6vgGC8e6wM4Ume7hRslbFsuKExAcn0W/v6VgydkYsTIxgpH6h8+PwAF7e5mtS1RSCTLNEd6Okinb
u1931ZGQtRNSJ1XUioFeHDb73v88EUj9vMtcesi3wXm1RSKB2+eOb8uVcTujh/bEnTmq8zrXZGoF
/ayQawb9d8QHiJuexlTyHMhR4gV8045gwCRqIz6wNvPvWTANAB4ej2TrKlKsNr+i2/uRiCeU4OHg
aI6/WimpJwGIfdcd/uG7h16oxGwIDfkJpyjYTqppsGznFmw66N0zhxvWrSLo1uHLKc420ks1WcYF
thoFvG4MbJV5rlSFlRNtT4HmVRdT7PCH7ocaTssvz9m8fsf6MVPDznwf0lmITKmVj7MbYyWGebDF
yWSik6XVazSO09VJ2X0hModXXZLq6e6dkTCULWgP8K6LYjl+7BnVReUnlH1fQowiIKL5aO1CX/oz
fqzcqOuzS3+eySO/Kto+hlEYDGIgl2d5nDjA0BI+aVjKo+TiEOz4nrV+HjHsSKKOJ1FZS+fRSEJ2
kKaucMIn54m2MzayX25qtcEc4ARLupak8AwyQraRTXohotoiFPhoIqcE5uk69m+k68V+nIasTeMv
rR3AfmXSSfEI0xMXn6/v77GKKVtzhhvpUdpffRSvbDV2YsooiPXv9hg37pbDjFWIWRpSdUA/uLQQ
iGjlEx0us7xN2ZVjmevaF99KsBegtF3eRmMlJi73iHtni2xD/3B2Cdo9bsB8nJ9Nr7wrU2DEjQP1
LGk6NBawLxSemFKWf9S+v/THUF80342Ql8132PHM60sXerzEMO7pfVqGHVvYlJ4lXzraibk4EyhF
14ScY4V9Z7ky+2fKTYaFXj7mdyO2u4BvZ3atAOO8gsDbXuASAR+qIbXppPvOXVyPzD/J0na2/5P9
RLI5SMy9cJQXM37255e/XzDsPOoo/K+MKz5xqUk7X5dWSbvSRII/y8PU3QWe+E61zvDtT0jF+avY
uFQJxJXGNQeksTTF0ng1ZO9XZhK0a9ShNGSa8b6SGKDG/rt23yQzpc4SFGN43NiStEw40CcqkCrO
lPh01Mmj6IQiA7vZPp3vrccsy8Z2Tnco9ZkvU0QzTZiluCXWY7HmK+TI/Cw5vscVSkmYBdz6loE5
Vrz6AahOrZg/AZHUYguNk6XaPdqrfZwLim5ixqDPlvQ7btQD7kJQB77p63Poe1oR0tRYELI1kjVM
IIj+02JCPM6XNBFQQGT7V2HaA4PQr0uoDX32Gl9w6EEy25Sfv54r46nsytBBHRp9iXlNKm3+Wx0+
J8oPBfYGXFTWtuRJ0sL76ZW67C8SG+hqfA9r4EXypxFYGo9lMNR4ZhudzJdnPUm5VXpbUksFgbYS
V5InHESMFT9Zy2rl7C67Cjt/OdtomRqxsekmBz0PKR0TwjEIlNoiyf87LHO1A6XUnRbieREGMc/X
+BkFVC7dGYCa0cROtzcY/hPIjH1TnlmLjpXZGZqA1g6A6IoFgmxZw0mNBG+o5wUZVpY7180tBF8X
rplKOdViLon+bYsjHC9wOamgCb7G3GP1ILklQUQTy7QJrVZO+iswYAgbb9t66BxHERq2/fXT2saq
RV5+0BoS9YF5oE3Ji/TTDqfStkYew9awVf1uTTl5GBT6gHiy8RWuNV9LDrlA1cB8cGb6aGDBZ0qw
GlfhCJRZtdKrqkTbRDOCr7nmjrClptYSQEUvwu76W4XOHC1eeyS7hOFKO//FLKdxJqrsaBLQQDUt
J6F18MvuHuj5aDwgSrefmtaUb+02YYOfBSCRkaToYAD1mSvEuBuMtNWp6p8qmhrL7gMsjBWnip/s
oNG6gdYuWk0fpm7K50/vA55EYjH/wcWZJq4pSYV7V4lTS2vL1iFOQ4Wzggtm8J5BUMt6pQYlHxDV
nNuQNlOAh3EAaM1Sks/KKX2yCffih1774SVzv55Ad28VaDfDgqWUy/5ePZlPl8qQlkmJJUxJI4zL
Uy6jMcOSlaSph4E/bYb+NOb2nEnu9qkM7EvPP7nbmE851vlpQOKgRM0nJpQiNhi7pFyehMQ6nR6e
Fkam94NVodNG47J/dDbpSj7hDS7eX3JyXhmPDZaRQkKINsyJ87Kx63rxgM/E3T/gHj5Kt47P2NCe
QnxqtGGm3F1+UUIsd3JrrwJXJO5QuU/DxUPtGzcazNQK851mH0LPSi5vI7ZnlctTcLhfBjxAZFeC
fuHh7X/u+T6SgmYXsgTdJUrx56Fx/L7TbnTG4QtV6k5JbYp799wAsrvbzuxz96kjKpFhYzM826Tx
9BEo/Ea+X9UB7ceWcmSqIT7f4iA7ysZmZZM3vd6UcuyeY3Odt42UuIr/mG2uuSbyhS4xiGmCaxXS
eX+iRpwCE4XjFGhElbIcIdzQnTSgqF34TcXj5xcg15A+dOSL3xKRNYJ7PSBUJneIfr1ij9pVd8AG
ewaK/MhGLSzWfC7fi2ZNGpiqr1GFwQ8783PXcJ8cBr4hK+UZlGIpR3tRQcUrQo0DggPBjeMl95B+
YndNsGCfQVSDNuLCylDwsJ3bHDKjCkBsv1CaZVXPOXMekGk7Q40DwPQhWNMFAnVK8Vs7jWcP1bj6
R6JHN6WD3eQFuP+JLeBpl3b6ipLNNgY3TgVTzRUYcE3CgC4bE+qoLAZEnRn5deIhylSmSSnRRkW1
zcsStfhebGQyeSBUVJtOPeL3wJ51qnM/xEt3/R9OjfzXRbeVcDd849O0dMUsJx8YanV4Cmrkg30g
C62j3P1R1phsfX7a3spQEIlp/8ldxY8WQR7Q9KOnfKVD/JMVwMZX76uxJd+loB6TxgEFwAm5l9HI
ZUDMzUG6ymHOEQ3N0fVu7Dth1SuSKte3HFbmGAhlkVD1h//ijxkus3RRbiRlEPEAiKEZz0ofpjtN
DmyWhpNDz5zM7TvhkIzxHHwGD5hxknS5V3Ds4w/nmmRaflr5tbUkZJmVb4cCGhgSGnaHJ0MiV2DA
oYOCS0P7v0QQfBHKViEPJvulG8DCFVXVwkzDRQSASnWUtUDmAKfRUDvmbpHmJ+8X/iVgWcIjrY/0
pqnK9NsDWYNoKDq5d2kpjA9r7e2XvZKboek4CPKdof2BbddMkxyYPpMOPxb2YXTQFM9GByj+v7bx
5P6xnJ74WIrDm9yRfUb625sZCFGV/i94/aCjfEz/AbaJDU5QQH0XDfQLkUz0hy4KeMPEjT4AUyt5
3qRDe3bwcu/0HPVUMyO/csYCwaxMVN0ph6+K1ugLoDm44BuvlJB+VhKti+rYS9AB7bnyYTcaE8uF
YjWctzDv0RITyqzfOqNv+/v6bFDgGdRwHUs4Qb7pZ/Fajuw++OYeqjVlt7w0nExKNxA64e4nVuc7
CtZ5dFOdjOrnaB+x0vFtrkk0YH3MwZMimoSeFqDqpWpAGYHhDaHyEAAvWsVAj2kzWjQBJOVpDORQ
vOruKBkrxEz3U632tbxhM7NfIFZwqcaW0rJlb/hWRYLzsS7cuxMtTLtRGDGkUBlJpiVRog1I6uDZ
JtcIPMCbRQu/i078ng7svdwJKBZHufTEIZDQ7z79f0zAixy63qYmXNOvqdg1zQ0Xb5sqpXY2mE3+
yLq2c1zbDkPbzPy+fl38M3zxdvX5AGA3Iaq+IJ/Rx8qArRbyTkD1bWtkLfwFr0Ge781FN0wW082B
PeTMOZkf3GHcLk7qPEhcu0Wg5/JMwXCheYwSxAm0ZoKDvQVyb7AblJSh5u9ZXCZ5LuQnOxJ3LWB1
e3Hs31oUV/G4gmobrO5bGJF1V57csmupTCiNac/L/cg7uL8TahTGgSarevCKtVDwxrpB5gvcfgFL
fTICGO9HTlsU/s3Hx8vO88VwnUB2xqE06vtW7nAQTb44k7tJnu79Ne37i11JprxEA4uIi8wX+RLE
aTaRvgtDfhrAGugZr3aZTl8ehB17NFV9RowWmcE5Fef92j0h4IVKmF1YGaIXl0CKLMI8/UV/O7gL
QPb6bMgKJDRtjzuIMGavFrTHeHKXcbY+qgJVXM6cn7bz3SW3DTcSOofv0gXuuNc9EuJMcl3YIDhH
fVzurpohqkUZslfx4iU8kkv4IEah/S86jNqzUUPpmCj4KAeJQlou14YkQak+hLryiuoISwvOJVQB
HJLMS7xn/att96Py2Ze1StbtP3fG24GZ1lCsyKeTXYwEkQ7OG7VLInEuhR7ufG0fZjtp4lSJv7Ch
hGxjop8JdFFxBk3vW83gxg56xBHgBar12hV0KSf/XEtJhNRjn+8ZP4GNscxdvNqQWkVF0B6exTXG
r4QNIw74cUBbSWyJSSUgQdklYQ7LRVzF4KYw4XaZsXlSYIWyX7V0VqTewoWnEO3UxLYgcbm4jcYS
Gqg7i0dgrXYTeekRwPwyPSyHP6KLtgbpZzf5UWfNrSSxoiLHaOemu64kdsypiQutlZIQQ1toQ3N6
9vQfhZBv340eqVAIP8Kcdl3iR2jv7Pb9Tv6MdRH6PnySX7dKC0uIsqbB13mhRaO55RbAuDW6N7bG
GSQvvLSsTkXHeILAQlPdGk9Mwf5eEFaIMZb7Uc68yXbb2a5jzkH+4nl4mh8R99dKMqZ+W4Uqh7XU
jqWzXlE61ZzzzKylB8dCiwgCX6KEItyk0NOK7CfuerU5WzS+9fwPRBWG3/0CMx8ozIKeA7hoaNnu
EU3+GWVl/bJq6I85xe20GBngXmA7j22VUYSUI2JUSOGyVTOMcXHv27fVG1cE2508QSEFb7BPvy9Z
h5hwxM5AIIWHTl39c2MhRnl8HKYKRAUvAUqprrvzfIp2AqBrgOIceZqnYlX0oU5E+F20TPcBsBUC
tkgnkwNst8PZSEmIAGahar2yAhnU4/2ws2LOF1kidjyHVIY7KU69h6Dd+wwBk2qttT4Jg9UKUXYQ
qMq7mPqBXJyHNejUg4YvV2lc3mkadOAfAj2urjhmeFYmkqqg+l5wF9IpE2H/47HBIMXAlSjXyFtI
ZlB9u5heaNxa00Nns6IuElfhU547cf7SmKSO9k3p3ReBkvwj+lxn5U2ViU9RFlLkLxjdLTCFj+ch
t+Z26DmcIqDwJIVYvXF8uO5xh9yTrN2dDcbiV3kS+P8iVwuBU9SOWMnaytaEdLMBdb+XYo58mVfK
GPmucxW8hKZrXOwNHQ4ORit52uzCN1D1kbCrOoXtYA10mA2o1naVfsu/pnXoCrKmdwv44I/lAWFr
vBnBWddABPWLnZOK1Qd9dpPlgcLc92aXlnnHaHINSMJuW1ERDFeX8ECrcqeL1UQibWzDYjN3Ypei
bxsz72Lb7HHEM5okVslbZh8OgjOFiexVPNhc940v6ssMRiYdwwoSDodFbFG7XIZHZgHqPd5zURU4
OPXJih0xV4BttMFO2tsT5mKTHh1nfZJXv11HJLmCxvfDJgGV7MGZALOB3LAwSKEwyDie8cBocTk4
e3+HylzZtO8P6fzp8c3PD8RGc2FxRrQs/JqhzBLui1xVe5tscGGnFlN3s6QLUi+RptkbylkfJi71
z9WtRfn47hedhHuyQmWPRWnZ1RDMHPycKIY6djay9Q22dvv+b1LLJevhUZ4URTDxpJn+SHr+068m
Qq92muqOGcN6woKpRThSm/rWR6vy4Z65uaJpp9Zjz878CQjZNF7Mst0nXNEEKmbHfYbwi6c6Kbfw
FybhqIxgaaPTBI1f6IPPgi2WnmxAGBzO+P5m90jMD+sBHlOKkPutj2sAUq9bUEPL4C9U5MOv1mB4
fFhKA8Btylk/8xxQNZZTfnzAq9xF1byWqkUUxwuvV7stnmdeGn8+9vzM1rMzxTz8C7mi2Goa5DYE
lKwikucRjV1+nczZRPf77AlR88SDAcin7FrFegnj4vLYCmOapj32QgIt1jfMJlSS+oy4RLkPdylY
MtOhp5KYQniKdJIrUpurPSuuyrfdukgrt0SMqnPfJ/STvcd8MQTqWLkTZN5sbX8mIe5+ynDmVRmG
N8VJewoxS5Z5ZsSmOof5VaVbpdhG4lSW3Tr/DePiUOFTRn37/fZs7dr5sVF0zXXS2KvTdCwjuXIj
0duA3elraaVEeqcxXjBal4YmTweg7RTP85+Bk0Npnc+syJZ8DR0LxGkig6KEUJJmEY5nsoCCKf/y
M+wqZRDX3fRzMLCn1Xf1Ma5ETCMv/AWs1JYgZA73a/RGSnZmeB5c/TORC76Rbfx+sxJCDU/wkzCB
tFYTqu1N9RZEeV7Y4bCxcAxqMQjIP0bwZPQE/k3wJ5cBCTGVDjUC6wI81MdmqlX7RcB7Ao7ukFPy
zPu/9391SOz6R6OT3SnFaMPEOUwy9qI6W8QqyDRGxHqAyJT9t3zzeGwmyaaGrKPr87yx3f7mw19D
aUFm4vW6MiPa8iJ9wKcLoib2wn6x0GsjpSVeo+bAMGIE5TYDA8ZJd+jxLBGHiv/ZVinqp4MNYRG8
6oltKCIHSBaKPjL8fdkWRysZqgpSpdtzmH8hoXnEfAm2JCOBWzXXR/O7Ba/22ixNDzHrlZfDUt92
QnOtxRflRiSci8/rarNZIcAf/zreizlnSizwQ0NhNK3IAly7VUNoHTiZgoQU46ZFmafuZlxsEPqF
5ztcqdVyChvFQH+oiOu42WwJt4ZyYqvIvRDYWbygNHvwcd6aR6kqrr4XyLsUe/3Tw1zVxsD3MJJO
izt3mu0MhU9TUxtHPElHmTWq+HlqFMk0FV1ATiwnRap0H2MFnSQaH/R9tYgToLbODOve1lRhN+6H
AulrnellpKH50QUQODfnuj5cFAzKWUxNeSV0vWH8+iD+wP2VCEygf0qAQxnq/KoPYYLY1DblYbmB
t7TaKJoVvSV+64ib0JntyYla3U9WkARFlRhMBL/V+S0iAp5szzW8lg803yIMboUYmh5rcExsfS80
8oevZE9/b0KTTspZvy1vAfpT1I9PgAqps1iJhcis7LUGOcln50RV3Uq6Wqj3VW0bnfqTWnoP9Z2l
+CiOtwoHd0is9jvdmG/KJX3yFVWg+myiftRZu70s8Z32v5ZscvhNytcpHXucUYLhJA+Q4/e3RNBM
JC+lZOcyjkRwz5kNOrfg28FTjX736Is+X3NsB4e6kjoBcf57mQNXvAPZLtLLzpv/DPbb3I3K1pxs
zhbejIDqmi9Nh2sGfKqAV4B+oasoxwJcsb73ZHbExstkJed035D1CxvhXFm6I9J3rhaAmTaxWJR0
cLhH1jar6gAyAnCK5Giq6FoxV44tGInxwCJgRLBRzIL7I2PCjowFL82KnhXYnGFU9vYvLJmIYc1k
+Etobv1gnBJ0c1qiNZQuKeJ5OKvSLDxBYpdi0Qw5DrKjTwtKrozHHLKrk+5ZczhjPguaIUvwNPUY
NsWHwYky8IfamAZ6kNXNBukbv0fKWdB5ZIGyXqNDGqXMSTCPoV4GHL71Rp7GqDyQSiShQfKgR393
y2RmbW95Na+2P5r3UztMks8+w4qXMAfepQ3gjU2aRXQxYVgaaOEzZ74fKFXgIDkO4xkzKpCd+bu/
23dMPr6TdgDqrL8W27dP+YX7+7Kb3aQ9bkI0TiKzj1mAYrYwgwk/xGyuqTr5HWP/h1kcGOVw6Iqw
/iA3ZX3vOD6/qNGfJlYOY+jJjqoHQSrHabhGATHL6f0Bj+XiGywqlj7+SkwMXElhcu7m4Y4V7z9+
VKF+pM0K/co7gMoIydH1DaeLL7yaEcEcnLupXh04KEmwRheJ8RwYw2Px5IpiZHc0fJXCNA6vj2wW
6K6bZrg4F95VpsMioqhjVBH0FPOJtYx8Ns9Epm3Ao3e89lLsLZ/EUiLhwjCR+P4SKG4pPJE8pMqk
gP1d0KAoUCZgOBpUd6lZ4sfbKCidT21//aiotGMMlUlUKXuzKZ3iefB1nxtvfCEgRYXZcQSoQFiM
96+mgB8vCjZJBEXajzcpX2+ult+hHmHPYrfM6/o11aGPLajiO04MdrybGSbT0CvnJl4FpjdTSbry
0Wpa/g7MR0oAxr5ykkV1lFzMzsJTnBSZpMdDufC73oQB7NZVoHdWXNOOc3SJ3pfaNm4e5vAeLTl7
4AEj0osWq47umojjNLM+XMG7BDIRcr1RRTjiDAZHo5HWAqyU34FPokgCFFEcrAYpY0O/9qLjvEEm
3kL4dSDDYGR7lcXWWsCxb/77CZPgtmT/9CixJZkT5QlpLOpSobNCxJjqYnsieh8BudmnMRg/eURL
0X0hrGqMuOeMP6Dxtf2VGoLk2fAi+ryM5R0LVT0BgBP7ntnrRMExdNK56Oz8CoJJxWAx8vFFbHZz
DtEBradDegoUC/vc+T1+Jxuf4k9BwqaPfoG5eakW2ul8brb5er+Sq/0kMxXaiRL/MQ4QXE9nrJlv
PPYeKf4HNtdccFMXuA3rmNXXaqbC7L293zuTto/rzXhqkubvPZ+7mlhzGqr/l7GkUKkllJYyni5i
h5CbWskIXCtIbjfRZHY56/OTtmMkQuh1PhOyTZZnu+CCV9zt8LKLWkfPdeVALeY8wQsgm5tFp3ZL
UW9cnw5EruTIhZQ9JG/g4CsRe8+MeP8KGIG3F6dV2CIX6l/RVAUlk8nAcDHYmUFpX+Pw7XtGrSxo
LbcYMmTqKxSFFlv+Cf+t7Sp9idoy1Z6IwzeG7xhcCXQh5RGmAgn6ZH4EVRElRYm9DMxlYXvw8md6
1V9nMcYN7qIZ2MabilN+RUFxSPthOoQYbGtdOcoj+bO9m01g5E4j1vHDkcfJ6ymyh7/J2QZmMVTI
q3BbWvsbAQ6vR3wy8e5l2PtdNXTIrT6+2H+k/VHYcVEkaVcX8oJKD8X0bIq1Xa3vHdEnTyZhVXeI
ekyYJkHyLitiIz9wHZT/TLm+z17Zyl85gIEqTvor3nEEzXbZftWXB8wcRtfP9DGp0n24hwFPKZyF
YLrO+lBwg/vl7acbQifJvjZbp0rMDsxFmrCXR5lI0o6rfsatpvrZxNAuTnWossbFRRz8qvXYbo+s
LGLxHLzYQhBxFSQFS793z6D+9fPJW9DTyDme+vk4e1zNqyN+nXVgwm1PJbVTtsaCrNRMXRrrb4Bz
7fU6MVA4n9tlOwncKH0DQ3xGSfSwEqVJ/cG63kPhdHL21882PG3HaSUKizJecwORQpZDZx/rXpKz
8JbiC1kk9i7gOh3sj1Y48YCaqvb5TQ7TSvqghei8hBejxQQLY0RwZtQFXGd7XY4aVx4mG6DQ9b1i
Nv9tHJVI1JqYkPUqy8dnUnZ0yOFm8+yDU9rHWWwzpEVK1+SNGE6+nrMov/0z4WMuslFNfq3XPOE2
h2tdt70m6gaiIhGmBQDKmp28NGGwv9bhQpLDIpcDfCuamkAUk0YNauEe6Qo5wLe2BtX09KeNPL0F
Vjk5r/+fnK61qVu5ipn131LeM3weQc8ujaS181UIpag+yVpOw/v+9HGY+dVfJhpCaW0jUuwUIwPd
hvFjqQWFT/jMx9g8A5ypuOi1I53qAy1D/nSjT6fzEzXCS6+/Jx/j6qtbRxb7KkAp6Hs4eJ9rpgNK
L/3SNiot1Dm1invOm+1kuxN7BPR9szUoDUmdvU9qPYpQvxDXOmElDAlhiCbRApCUX8FqezSBPkBn
QsqddP/oyeYEDsGA960HzYbIhm0R9xbdp4aVVfTGBi4j0VNO0ZTtkcSHsdzhxKaHHCgDEqXPdqXv
EsgEmPcrgJHrxaTFwkVOcqzvUBxyUEaj63SakpN3lQuaRNqcjdrKTIPzruqNJ2ZsPZT4lMQzgM4Y
XhZnk1gSYZIEBYYYu96Zs9jSy/GmfsypwUOaDzoMxsNdOfBt56j4zpNZSovZf3D/5oTUufkbz9ri
CxcHn9LCQs+8I9ISLpjvhrDsO+PxjGVdQlhlmINHA3r90cpLBGdrbjCr+5Of+qQSPsThKspoJB/r
91gvLCaGLKCGq6SKHL5mw7M8nvcXAPys2oAudZX+AwXR0fEikHGlM4b1j0E1zVG0uBuLtu048ged
/9F/WNRLcnKzjdxEoAr4fwg+sW41/UisNTSYRvoO+rNU4M0hJOoK/mMnGEUvhhr7ZUQIyxQrU9Fc
YK1ptuFUjAbgKozEQLbsO0KF3l+A2zIdn6d67+DKFviKJsfg7rC1jMdk4TWzxRkoImcyUuqPMyGc
E9JMpx+Lxcf+5IHmN2NWTHDVc0Plxj+nUZ344xmCs5gXL+tY72wday1cMi28EhzsGGRRXTR1u4cA
0IMiEk1HjtNqDz04zaJPhvj+Kp4WWlhVPwpGVsxjob1BHP4hqtEktX/Rig5ktpvWPZWR3IPKRR3b
07KkCg+zAAzPPjcMRYIw+ZXeySglITF/JrEd0MsiyC55diEnjVAWMMcjTMM7CcD+j7zvwcJ3tTlA
ZC+qgkzFEVBcCDod1Npme5Psuc1bXuPV9MK4CUd1I129RPtB2mpvxpJgu7o5qX24X7/NuZWTsokb
ZCuLIfaVsa2I8HoqVSek2TCGieBFmZqFAiMT23OWQlKtdrx51vrgfn9kiXsFkj29kBcYI4T0G6AJ
0DfOZ698fKVuZFAIVaej+BKO7abSBpT+YTDGUd6PHMzhnucmqj3G4AUQzjaTXdQAhwkA/WynSmEr
p2/Oz9r1pww05yL/QCBlQCEXapQZWuIDz9jW5dmJs7I7E8m+8a0sHUZncagv+zrN71L3JJDdwh+b
+VgKgS0rSKMEACaMAl+R9WN6Xl5vRk8FPmIj5hQzJEk+wYU0cyqL+E4YmDUGpcCqTmeITg07Rrk9
UHNfBu4KriU+2wDdLKw9hbYCw7VKVO3Hjtnl/BBbWUufBAnk/Z1mlzxaYcLd+j2bhY5lg3aXZhS6
TbQj1d8MjOLw/vuAnMSjhqkdWP7EJsARFOLTXJf0bCAtSva4t3aRHk9ElQ2aKLEuA2TtMKS82fGv
FhFOow62D2wVj+wpcRiU0N1eve+azpSDMCOKpq75AnF82GBZY8SeiCCEb1NOALJ8fd0Gm7NrOkRT
p9xAZyzmBiKwqBoFWJ5YxkFsuKVFd0OgnBp/qaR/pebkSJOM/T0Qt6bp+efrK8IoiZPEdCihmexb
fhh27vTBWoAL4bhN8WjxisccAQzvbxQqohc+S5coTNcJYT5/OepK7B6yWL9GYELDTaVgkLToZdzm
1j2JhPYmuR9goAfCGzVcoMpA2ZCKdWC8/lr3RmeeQDOy+8gLpHvBEwffG10nCL6hhmZiqZIfhihV
JZS0e9z0AU+49Fro8Mnl6XjrL/syCpTTAmhbOOW+sqtSN1uyJDJ0mr3LIwde2HyoIXqvXMrKohfq
na6vSQxBQKjrPWm15zeqLcB0cXLIOv0Q7lZS16JKYRreOjzDTU2zsNaPiTPtXagdLrIeSZ5FwvZJ
MdjS6WK/mW1SoW8dEpv/Q/x8Sj3iNw3kfZ8+26DwhGmaLQTscwQF41P89nGmAkqVFBlSnonLF3qO
rwMEKqHR8Q9HpGQDN4X2a/Dmflv/cepNEm52uj9YqxishlQleh5hUBK4V7NudhM7UFrMY/MpatcS
bHPTzdgICwpfeihLWp5C7DNtW34DVcITpbygDM/w02vCpwXu0fJFM6gnFUh9Vi7sWBumugS8WU5T
epow2KE7YY/TzmTNUKdkfh6dEvRIss/FtpMXWkHLKmX/yS6jppVbsMgZ5w67bVj/NUHa4Bpdk/5I
60eP4NS+GDsnQSEZDsPfRZNlbZUqJPE6QbrSuFbfcxjvjpFP07bac+JiqyOoz9YtnIkp8heGeu1C
M2XpjoWHMSRKXl5iz1viVO+8015kVhsKJhbqdQN7EOx+Ypu2xQE17qUsyvo2aeD+OivqEN5buStr
gG7qxVdLt7juFQL2zO629PNOMlpODGKOVM2ndhcYtTloc+f5UEIUiORXGtd7qwkfQm/JPxSIOlFm
0w/RpBnXBba2NcjvgUFP0FiUooFD4y150oakRLMYTWkDnc9kw53gVwSs+xUPOs4ZZ/axDVeBA0d7
LjUufFI0diuHtykccJ4UVT5uErStKwlpsTOA1IpcXT6AozPFfutDK1apk6/sFg5kjFdIbtDokbeY
NDKF9N3NDRMW8YNqdCQBsBbRpHmPDjHTSayOo/3ucGhbZJ3skiasv9VOo9L2Tg+ydRdslWaqyNkB
Sn3kbZYnyQ7V788BdeypvnZDhSRwWVVqUKIX1ZQUKcHDIgJhCK9jN/fW7h/4OSAUHwqvw/TGY/zz
3ncJDru1JdPpPSZd9c3mDSh9MdLMdr462HU+hBeBZH/KUkGo0S7ug8wFfEK2pWHoqUUjEoXDwtHM
6O2D2HqkmV4DZXcL4FhL083vSTOr2j6m7OfbexhvPidBm+z5SyvWGRYQigHlGJRr4L1JT35e3CML
lqef+XK6i0933ZVp6BY+6r6SezLTmjuV2F2crtZhDe00fiGRShdapGFaR25ZTfpsM4Wh08Ih4vhW
3QJt15/zsE/M8tEgfKPZFlK8ZUrtwfP/TxsPSkuEpSyoP+Vu72jUegdYKebgZiwoa9Cs8iWMlwvZ
Hxe2/tgb3cPOUWT/NiHlf6lDQ34zNAnqLza2Pj7RBpqpyoEpa9nSqHlWtU75XXWuQttaBIBThddW
nQErgzoL5beL2ofx8MXE3fWDayyjf+sTQJpZhYQABXLe4X6nynICcrvewhfMXQRNTbGCUR3Sa6mb
YSfK+1kKqHf7vfPesM+LL3uYJRH4r3air2oTAI2KQKggRPiKisQqFb5xWs7NbSkVMmAfwE5ViLDn
cbT9k63fvILx69d2GqJL55+HXxWbWbQOvVE4m8FUBnw6g5mNScn3P5dYYmcPssJkasiW8LxV6t//
0Xdaf+DRN8opfrBjEA0LhFY+vnj6RBvlSNTTRMaZ7RM4/UpAi2ppkkUg0/gHanbDRcYcirUAxYZ3
dnFJbEeWsem0/55lD7s37LTv2g93bQmju5nmL4fU3FEcqfHCx5QEwf2Cwn5tXntKfVprSsYiBrvh
1LSxU7lMlNdeHfE+tJD7Szwaa/FtnyIp/iVE5H4W/sqSYancpsr9cBOe7FvpW0741UPMyyCBQdt1
ldO6+qorVP7+73NiU83q+WDN4wr9I9acXALU5UFooPOgktT9SFv672Ufl8W87ct8JHwciLA9PXJY
sYvjEpQZWB8CJRTUkrvkYk7W7O3KuOoGlpAjTCdQyjYa48UsF/gYt+CtdoZ4UgykaiA3K4sCwSUM
uhxLqMJbWUJEFEnogV64cZN3rnA0pESZ7ZnX+SaErR6I0AKF3nZ+41YZhinIQpwazjXSV+NlN61p
P1SENZhIZUPyq56ZHDwfgQUvRvbV/KgUsWYk9QO/bt0PvPNlVXPtJXLHAYvVTvSPYNKJDqt7+CdG
wSmEf6GxYf3XFVX6cgYVHilZmYi7uT0ixKWxUfCwoTLIOJaGYwlZcye3cdHLFmfDSsNmYGnBRnUh
x66m5GV/OcIlQ16tkk+wrFEMZ7KFRZqztKc7UUM4qjahdrE+c2K2oy5PPczvKn5NN5le9PsD3zZM
r9TKUn7L9ISpefM/hQ5PIdyXzpdKa2Dk4XgQy6CzS+coXvizy5zr/ZQ1zMul6PzoazN+FaD3ypdY
/mphBW0n5FvfCdgjh60PQwxrzSx4W0QXEjAftpmQwZvxTJTVM0R+I7hwOzubMHd729841vAiylh1
DdTuYZ8qvurR68lhihBNHBImyXNg9s4Es93fZ5/FXIv4G68xpcEye1KcbTrMuxWyQs+dfd6hzBzq
lOrQmfgWNZsQ4N9ot5DcV8yN9n2BvRIotEPWqHBfedUYFsFRT9cyChdS9PA/p1yr87Mzw8KpFdn2
dR4p9hk+nBHXx+irnp7pmGh52b5zt6YmDQ63AKb1xuJ8BERS6hSx7/2FsWxPhZj+/XJKDyux1VKl
XGkXCsCv9HfvkXsKu30ntyNE1rX5g/6xiyRyInTvPdn2/0nfhQGtJXHwA2TeXg3vn+WhcJERGZSK
fZX3GhIpLV1MqFlKJ42Vfi0lueXA4/D+Trv3RbAfYac9JaG6rjzRNnXcu6s5pGlEqdoHmMrnNKVF
9W5NQa9+Mvj9yDvazkr1RBP8R5RFOkLb4N9ZQPMzSo8AXWOhkn+DJLuiROITI1tGoVeOxVqXFsrg
O+u0yALkRbEGhMXIUdErNmKSL4C9orkInu/1R7OX4CHl/HkYvoSEuzPQ6IXTG1Ogjzs4DHfyd1Vb
WXBnBsb/CXlGg6sDABBz3C/RbCJILGzi3jPgl9SZz8/q1VecLiMle7uszTqfHjgXjdE2XOPrFSeO
SC7AM6tGEg6yLlCBDVAL30H92RCQkhkST5Hj41ziAsVZWa75764n20VrvOqidKhLiLzf6R+Frzth
xTatzqmDWyT/ZwFIFqB+lA6NeKkv2iPIsnPtZuIefnIHyOdzQzIh/sPB1jbsGtFodasKtkIQjao+
y9hGBrvrmpY7KCp0y+znTYcRgjOma0B9jafq5jgi7Y/rrONM/sLSDkBM9GeV/PK4/fjluL3TOnNh
XxD11b8KXlZs9l7aNbv+zvkriPO81G9ssZMtTeFrbJqH8VcQGaI8ET+Oj9Cf835Ms09RCSyGx90+
TPEUtxFzUJ3iJcThWKVR8MCKe7VAzrWi3edmeFWskG93Xvw4HEBlZG6Q0SZsEVVrbGUtZKQOOhRd
Zj8ggZn3EjQIPKcoW/5S50/+Qhp1sItjger/HxcoSoPVa7CO3hWqdoXqgMGQW0+aDL4TlzNtcd6w
M6ceg920wtWi4PYPVI/SfdOAhLNF2b0uBYOLkzeLf2bTQVWp5CdVBlShLDsRXdLYPwBA3IsyUJ3M
HZsyUNNIi0RZ+yasHH6g/DvtmcZPJL9hMZJlmpNY2HVMyEpR+bdMn3WePE2N0/8OSs/OjqBJTCew
fwDlUlJ2BJD8S/1A2JEKjw7oeZYgYWUAAaEWH2A+mrteGkwEjGltrNILUVaHT92O6r2T9Mle0c7i
NpLtJ4gKoJz2Ykvw7yVYdxX4pBr7lg84slfxCaGUurBYRMz1DXYdxgo3qsY/ESNE19ZtkV6YszVP
AJwFO2aP9K0dLh+KgnoCXzCgEd7nidsuOgKRzbLYHVy3o/bTsoC2M9rDg0WBxH4rosVEGJ2JyxI1
zWTn+IZFQfq7LA+3Nv8cu2zV1/vfRYMKlfGf65tDkYEc0iADkjAaiABE+GWNT3gbLk9oibx98U90
ktLF160ii2My9/OOj654rKJCBH2ykN9UtN2bOo5b1UEJUty+2Wxn34Y+V9kRe0XYgDIMCVEo6qVh
wHiK9NKBvcFJ+xwEd/GeIqrWtwl2b5grw6T2pa9bFGVda+V1LutuhmdZlo6oDT0sfKERqtNap6Xx
ESy4Z28an904RNEBH77sHrv9aafqlsvfGBXMpBym3P5aPRDmwgjBPW2o1qfYrhHXW2/or7F4DYi+
KF1c1Y4roOrgK4Y+bICUerGGJi42HuFw6TsUOymL63Tat4ztWv6guj4RW01F+46vwD/aVONq4n1K
4qISxZiVPh+X6mRLDeWxMV+8dhDqXM3zreNE4RLoROcs0WEqIXHLYcfXIFwYZXPaVpsCRsPsCVxs
ByyCii+n3ABq6DOCA6j5+u4d4eO489G9U+EPMQqLtjU7d6dw6rRALoCGzuLBdkypPGPqApMIFcqv
7nsN0aKAYTLnZOzyWevjOeK/xcr1j/nRVS3LE9q0IsKYB0R4f5/ibyiPKqsPe1N//FZR772uc+sd
pk+R6unfcjprB8iasw4JSqkpIaTlk0sDEdd+tb9EAH3LWnCek3xqac8CwBgZvnwVvqAzRY4gSMuq
aTHc1pZ4o9VNEtw5ZBXkyay7ahEden3Yqt8edSGMup6Sc2F4vWmHOylfKgdta3wy7t1GrZWtt863
kCF4RLV8hTn0MePs4SGWbqz5KUcM5XT3EbrR8SHaZ0CXRYSTVmPZLj/IoUned5R9ztYNmU1k37z7
jsjiQ4fgxsnuAaa++uOUvb6RP+3tnfAAZtu5ALT0pfKte97L0pDUMsycXMluCNHeZxQ8twsJ4+gT
qTIxvZZK6SDB6fZWIcTtm3ISCcKm8b4y4AfSA9njJr2KQlD2tdk93InWuG0u1aKqV3ZWmnBtcXgK
hCC3WzskwHQ8wZfQT3mpYionld9AWX+2ZUSzebGKxcLQ87fjFN/6oG6Av6mTb6HgR9P77sLG/jIA
UaMVRl00fplyxsR1ei1OzOWY2Y6KLbX13pgh3FBUcOJFohm2T0JEoX9L+CPrsZ+AntJ/cmGbtDHn
5pb6GAp0aQwL2unfezkNH0F/cq/+TNn2HplDdwQrBek3iek5DqUqVWS30f/uiAy3vFYkLXiZAx0x
NO7BthrIZCDq21kZJIuvT8uqMMrsGDb6iANZxf9xgIayA57xyWzKxhohXDzvRuI4y1f6wg1Ycyj7
ehWztIXXDtKowhw1bjchgcsJWqYHeoPTbBeQ0SJyFFVzeKzKIWmpwdCYzjrtcnCjL0xP094IWU9a
D2XvB8fLa5Lr4S06SXukPrtBY93JHFc72NMb8dBqWsG4TKZx1rToMyYG1qr6jS5xUZzMoo3+qcEz
V4ZueExRSwFPLwilwkeShVuOOX9jMx9Qdv0/teKdZkYQXthjHfQXBMoaf1rTjlx0Hf7ymGtx3/3G
Io+WclQ0ARBKW2ggFM89j2P63pX2H9Wh+TucIgsirhuKhYfFM4g/wJrcuhj1tfKDxnXtJI30nTSz
PTEF6AeMFocx0NiQBdNX30RcHvHAt8Y+qF0ZA5ZQ2M+rTdueWuJ6sd5/GjwRp/4LdThlqkPitLzH
mBbhsPIIgHyTPLkTuNNUHregUuoWjgcpG0P5I5v4FQXwQKeiLCOijBaARi93tX39i5zciy4/ecV4
tjUE0UtOScC7xJheef36p90jb/bhHxrBg82FiUW2VK40H2HrRoRe9m7BziaDl5MkdvwlV099PMIo
Qiu6jXuo2+6d9NQhE0Y4joi/N9b0wXgUJP9Pf23v+kCIozk6Dm3NRQYaByBvlcVlAKgr2rkbncuk
eaQbyL+bPxU+I1uCxVZy91j58kzXZd6jDgOTIHM8OdjYRfCoem3RPYK5fMrKrr2+oAaN8S3XP6Ze
mOoc89UJbOZ9T3RfUa/o2yvqCtxcJX4jN30EvLP28uPHd/kMg9817p2QlQSttiiXsMSfBNmCakWw
QDBvUL52oEl2bMuk/uVhG3VUZIZuw+X6gNDE1RZuePggHCRoy4Mp3rhBq2dZb+SlUmJIQDUm+XCr
PI89XqbwZciYkoTMj/YYKeR8lQO+4YoQumhY9hKczBpYfl2rSBkGnC4GjmKovvm7B+R/1clcOYc8
drPKaBpMqN0fW+MTnqYdeobdIS459dDumbVLgxzicQ9GUDr/uaTa5IvV2jQBTT8W6Utdeb0pOxtN
Dn4sSxpVkNOav77LrIPhbXFS49tjZ3Hv+6DAOlfe71d6apOzCmJNPRlioSsoMYEAT0uVN0xaOjPE
rCrZ/sdSdbXCTx2MqENOIbdZIpcMy4JD0c2iY+qFcY6QOpbGqQ1Q0vhB+01TN/Iim3snqK3nAQum
moKms5fsO+HTExs3pxqQO6ldFT2cNyJxGrxk/0ge0IrjNmlCIJKgE5Ukw6s2s/usTr7Xd87AuoSV
H3kM0hL7JYX5mPg28/fuN4kj3zyVnJpH/nBzuW1q1hoSn8n6/Ty/ZowDtL/4rshHK6pNv1y/7jJF
TFqXRK196sx32Ov5LV7noUmMdC1XwQDOTbebo7XpfDHcLODDa2F8DiRQj9ETHDEhgChqgOZyWYb4
zVsSmF4KshAkjY2z+VkAWuSq55B9zrmQ4h09hyZBw9OOn4Stdj0RzEH+EaLRev8TQfiQJc1TKcIl
/prFaiBeXayGxh3BVMwcbrjORRm70F7N0tX9pUAGPZMUBWvZZcZ63uvCTgLwKBYri0psr5MLfPY8
EJ9BBnQI2r7u/3iwthBYLmqPi4LD9yfcnfLd/ciwn4IAobFa7CHf20/Nh+xKOOwQStvmqgue8SrV
hNXvEODd+uB1y4ftYr7/szuICJFj5DYysPOQ85CyA+HbAkJ6Ian3/5oaHeRFI2Wqr30IwdPvdh/H
V5QKthtqPjcQriOU53Tqgbj0LxtlY7ZLIPuPtV2t7nltnA0Meu0+ROSYs9catcYz5lvmNJqTfpdb
EpH4YkpBKEKPmhfRIo0pAp0Mkvjx/K3jzfa/WHWZ5qqPwOQhbDZWSm3kOoLf/Ezm5PjSbjzDbmY8
xp5PqwQmiHjP3+nhitLTjWgKidXXHnGMg9VZyyi7QxyM59AxsUvqin9jyxZCs6zund/mRNxC95ee
88kJ8MjFaAmfB6LWc9dNLXbFOpTaTX3UXWE95N3bGJj22bcxTWrrwgVI2ub6Eo99Rx9rqdcjGSZ4
UoJd5cfEDRKYg2cA9nLDUCERbhZFnbCI4u+7NZ95bTb57pQRoe4Da7qj9Dd9eaVroTaNZutoTTwb
fvP79BDd/sc8w3PwJFzNTcQMST0UlcWIJrjheUrvAvkd0xCgl/DSAEmPJFrIBrRAJ5jpe1V4agw2
bY50dO6PA9TIJ7IMg5JvzTw68fArue6Ass230kb6HsgzJnZaK5Mj5un9U5ENl+MitY47tfqTGqyO
Xt6cmrbH+fTDUTDLziF7MWcNxTqfD8FiH2YQSbjikbBapDFXBFiMn02jx7YiQwueKnSK6fsm63tm
UtQgb32ddHC6VQmy3PYkh8JYLYht84EU2zxXV9TqDlokKHyGDjNDz8FyoaEupoxh2q4i0z+xkHmX
yMA+MLtf+3ME31SP5TKLaJ/kMj0RblYLyGEJTWnCHIvd8iGsb+iJeLcjE6F5OXrq8go9kNrfjKAX
SzMdhIONgC8u1BSTEUVzd7TxwMFvXtqnajA3AvoWzJzoYm854bpyz9eQO+BH9CFrUHDsZi7kjqJn
kYwM/jtNzwapm2ZdoDRFYUyNlDj+nglB8FI28rDsQgPyQCRlge9h6YrASNMO6qoqEqjFM+Zz3mPr
+6BF0nTKkvrRQxURLF4qZJ9YWW/rmf/ZToJpTSA5NFEHuVLZr1ILTYc6VgwgnMqabPd5R32F5aEp
A/XcAFGqRj6Hozoe5ZtHaIH2Gh4WK4frFu6s/FNdTSd/xxRpc6SJnUMwLXIVO/mJtzLBNgG3ykPe
/++5zAf/HXOd6O7jhXKNu68j/CVsYKTCHL/+ZstTIE68XqU27qDud4jZHWkxoFr3HxDeMX2n7wEl
P8p+XM97TfWV9eJ4eNq+RhYTqwnWFYLrpMu+Qh2+i5YfSC/TeN+4ywAHGzw3wE/Bny2NXj7uJhae
3B7IEzZeJnvSZNnMFIABOnSJXLAzRk3mx6OzD69HQ6x9sWL2PdjVWSd/ETtr+G3ommS3geGSv4E5
rtCfUrAs3ZH4klRHoFG9SotfYIzPtLzQLnv3Ub91PYK4KKZ9mf0fojOcj/uKm5lXhF73/S1HBTQm
IUSEI8im/TDEQDNOZXASYprwDBvext9xgzRq5bvG18rZG9Hjd7tF90U82N1pqgHDEXBafpmSHfRZ
92IOcQQZLfXddArcH5mQYuI8yAknpRXr/CdX+IrswlijoDdN1Hyou4eP4Um0YvudwttPWGcBGnH7
mFC6CduSH02kIsIIBR+lkjyXjiswETHLwI9GRUHB2qM/lq0FA3mEBwfK3ltvLvWX9Ga3cY5hYVAQ
WDJubmnCyUG0SeahNBZU7WYga6gW/prowdYYBkIo3QasSDe4ZJC0qERlGkIaHNZxkJyzZGRkhLRF
PBzTuB1nefcO+q0q7LX9K5/+ATThdGxhPdBfubSSVfplaLCOFArOQbscAN+DGrwxnSSRjT0tkgok
01WZFsGyIk0rbgjICjOdCqGAl1HcGvNou5oGi7uTJQoU8iJYj1DGhwmIm0iVZ9KfHN/DknXfSItr
5feP7T5x+JNpl9FdyS5wmod1p9jRXLCljWRKPmQSrd2iX3kGC4+WkK3V/8yDd8E0SFJgbWaN+fDj
g7xURzrug1WrB7xoxhZPZ/iNAUlSvt6/g2cZ86kjDx8uqkSoNHUcF1w4KsBf/iR63sVWj0JhWCKe
L9jYx/VOccsejtfRc1au/dpkOecVriHXYzj48rfXy76BYcBzZUyF40uTMCaLz3AUu46rDIi/8Cmw
i44PNtgCPb6447RPF3Hzbk4kk7znH3hMasG2u+UjwlMRf3bFQtKBTIkc0gxviB0pI3+JWSLzUF7o
Jhw9bP7xlkZzoKSQr//5lcJjnKlZN5NiGTJGHAmNVZcSOPhZ1T4WjTj0cjV5c7Idvyzg0EPqElcF
J384mZLxMDoGuUzOb0nlbNU9jfMT+Aw30oyz0I2YvkR0T+aea+cIHQENMant3kSBgb1m6hvWBlus
smkYwQLcxbBX8mBF/LxtE7i83n6Z6TDO7Xn4n/Gsh+TdGY5CxHjLlo85c1N3J4n74QUXZ6SENdyr
VY39yvXUJs6rY/zgM0EV+Asiqm2JRhkmc5r4soPDnxoybp63MbokjBSP80zGdmg5W+KmnxtiT7XX
biUYajDn3tAReHQc70Zx+zwqgSZI8XaPnysvmVxi9/wtYYx6jEmJtSMKPA2gJMwwnc/2cny2RQfz
lrase61c/OISUQS8VCBwfDYh7Twkv3vLJrYJ7cJtiXKl3XJLakWAhDgZA/OWH79kteXcnx8H8myo
wJXgJq/taeyj5pH7dV/MvAkmyfAAcPx55su43ZtXPEtdziEt9Bur8RPkoc7bKSich94pm1AitEf3
bCcKZrd5jWXM+MFmqo/RQbJJWK/y9Y7s8uAZgXP8AQiRe+Fl9yhe4lywUWgWjIEma7I8W8o/hU1A
CEZ/EI7KzqDpRxlZKVyvpiiMlmlNu0F0MYbwL+/iPiNvlJlE/0nq/z3uneQ8u6kYdGn+p3KHjErp
Yh42AFkS/YtBqADlqTgJisd9+AXjzfjW4CJXkGNADYLASc9JJIO5jd9VoAf5RcMomYLT6hBOh7zZ
6pstkAUQVzc+X8omC+PfJn3IvcqqBHZayuVQJLlAPAV3zA2AShJa4/nkVMBlnenhGL0/KW0q9haP
5TqtRE4gLmPkR0JT1nJPmQk6FfW/CMlScnAprGJv/TMpdAHjtM08VLKUWIB5AgnllwTLClmttKBo
h4DwRpkEbJaoJZTsTKEwzOMJPh/fgAyxUimVuCOFjqXxapLSyZSN1/zj4IaVRgE/nNCEsLvni8jB
d7RwiUPcd+L+z3/vosopzdGD0nOcRA7RAIWRVjhpJthU5xlzRwm5r30ZeAa6sMAtgFcAQLKEZ6Zv
F7f14q+GvzxiDNziosMcbCYseSr+pXG3R6fjb9AjiXOz5gfXvddVXtiCuiyP9NJwIQY5I0p46hYR
+o73VE8YKVHkMmaAAdQwekjsJqgPJ4h86PHuLJCKHa3y7u2ny0Mwhc0aV/m+reySRnp7D+pc5Mg4
pNc7WRnPyux3Hw25E/D3cGWf0o9ygoECLPcP0ZUzBiyIwWR9dOqchKRft8t4jvrJsHVLv202Osgm
pt+0TANKZUpj7ClNtDDhQQa4EwgGKw4hNtMgaJv/JiTDW8nw09ZuuciVwCL3wE5YgWBpuJ+A5nZn
mC6hA6l7omtdqTMWzQ9eHUmB0CQTmUfXr300yJtIo0MaLJ7Uks69k5poLhrBVPDX50/nf8/wVw2Z
dmkpYs9RRAzWSKP9YHbE2+RyZyw+CRN7RS+HZtjS1aaZQCm3z0zZ1fX1hUKougir17+MG35HpU79
YA6OeeZ+7niTP4EJehD0PgdT20mvDtqycr7qkdphpKRS6p19Rlk0ZAODK4iA6G8MGTIh7tNipFUT
dwCBtAwhr72IyW3AhDKjH9I0zJTiLhTjZf1rYNUJUbq6sLXOKYspAKjmlI4s5dU218fkdE3SSuBG
nfZgGvmPwoO8gFHi1UPE6mKOetPXA07Ku6AY8mhSu9kW2963vy7eImDAQQEpVJesIR4ExOGLDySM
Rh2VPyFCsn5zOJTe000G74yLhJOr1k1iXJIsZg0sfksNpArJHUKo7WCAAaqQPrdxv36JIDnt2vCp
B4qHGR1w12iw7agVSfF6bGIausYxSEQ4A196QIdVHN6A5QtId9TlJLdZseAIgUVEAVr3kcrJGQIq
xbQe4eZmrniF7DqasHlpX0h4L6Rwml1O1EgNRuZsgaEFUTm+gELXuK1A7hUE44BSoMDtErhkELTS
4BSsL4dOtXWZVnXsqzKdG6CNsI7fwlofy7/QDJESleVQBjTF1jrQXCQZo44ZwZpkEpx/iRKAlqup
nu3IWaBT7CVOfpFkW+fTAsw4MqtRMMsfqmek50deAp+4QDRKx/iDYPP2lN84RweszsSTfDKQymIQ
I6dH86W+YCkwD4Tbh7noaRC4HtPUoAoQHlPI2RtbQF2XqbLPDQlQadUv6jFW6XlDX3cdSNyS5hap
F2+ZSIl8ZodVW+5DUXFKIZjXS1gdubUxdmPziApm1mDBggUVu5p+4feZX0pDzdJr2TB31MwrWjh5
Fub0BenH1h43GGd7yGS/fklxUPMYesGwqqFJ2fQjXXDCOCW95QoArvLVnCmBv+BaUAdt4d+duITX
WnTWTJgNjwneyHwXtaxypWnQSA6upoQ17mj1RjWaLnhI2wGdfK+uh0j68c+LpX2v7BPaX47rQB6X
8ukROnGZvQDIMTWdSKmdTSjRmXWmBDXrIjH2iUuO0glsFxZaV0DX7RE5ag1GpUFZMqBaYlNTPVvC
hN0bylEWhSLauRbs7Cq/iHgGEbfJQ4ta5l/5qrqpIFonefIhwWa+okVQVQcmTczx70OK33M4IZru
EK8u8kyOXGZzC+gcyuq4E0TUwzM6GfW6hrmCEaHJO91R3e+JGSsvL4U5iyGD4lIoaOFb/vJkqjGS
yCmUXN2trJvbLyJ47yCPQ7tpxlyjvs5GctB1jPtux9yjlPkz97uXMdwct6mlJ0aB4QtU4BUv2YTj
lYDCt124W4B8KlBu5PwK/5sc3kS5UFCCvtemTYoF2rkki8eaV+yhfIPRWLwRkW5LRqSHraY/A7U+
IMGvGmT9I0O/I2gpRYLIVT3gG5o/Fadcb9a9ytq/XJcvYsDls7cUFALFsgY9vptOmSfY5F63Qjmc
Zmfwj1qAIomG5q1Cn9+e6ANqmsm9u6+Kr+h2ccJqa3giLtNcNGJCW+p8D5DhBxIaxL/X0NkIwdoF
+Hrhgrei1/ihMC9vRTR+AHIlxMHXMTOkAZY1WEoxjyFTstTmJ8wh+Ygj+/AksKgZszsKnLA93XOr
CDDsLewEJk0wlh9yCocHuHOImLqjVl8T8C++LlKKto4+vfPNJ67Ey8n4pHXxv/IE27KXx5mM0SfA
9S9qulhhAXvC3n7D2Q7k6pYSAOzhmWZgXXA7MDyeq+b6M73vvwo4vS5sE6gAcR4iO2PfqyKcUb2R
8oQcZMIjXdV+KiT0OFuwJHhtXsvSIPtT2yT1nBSYy1rZKMaE+oEq1cK1y/yJFHKpmCB2MemReX6l
gKc20dRuebXOxMZ76DFbBk+DkLJ1Wg7tVrjHfhbYD+DHaBRtokMtlV/MP94WyszTAQDwcKFln325
UtYHPPJ6add636vUfJtWeli4QfZiOHLPGSqbtEwTtqt6nCV2lzl3s8DTn3O/PXmmMxvHSV8f87IA
BrWDVDWZYjwfowLLhqNr21oPOdNL2YHi/udChRiiEoBgMpB7vgxP9kEzQIRbGdnXmECvkBuZzzwi
v2fj4vN4gjaohL0YSLS7r+FEUqSDQXC6Y58lBgKeWmCYdh/ziAWC/uLq1m5aoguHGiCjIQrVmARc
OyRDAE1y38osLj0YkAohkbeW2whk2Hkr4cwVxV9kOEHf70ca8H/STYOgfgOT/hYJrNTHd4VtK36M
5BDr5YEiRKMeFb7sNv1GhfFlVSnI2dj7iOXXiFG0jYUkJl8m2unyB/PBXROZ98xtLc97JPgJjThD
8JNFimVgQENo9XYkGy2IR/zxpcKaYyfIBYRkxySxP4Wq0QMsGAi2p8PXcCO5q89rygfDRMqymaCR
l0tZe3/63Sx23zRvTaOhA8uxpQsS0UD8Bmz1DJK9RMYn62WGIJb5eusnr9k1CKJA0OOAjM96VeGZ
46Ql/L0iMtTYSJBR4ONgTShiE093zZZ7opFQyEY7Wprqlh5BzkkLBAMLIOgxh0UVFWFG+KHCxDn8
4sEAcJrxD+H20diKFXOORDbGcIDlQxuGdEnuTqx5ifJrXJdSwkFy9FM+dGqcIK4DX212SsR92kQO
Hpry3KB3IxJj/izFItaVPL/b5DQ/KInbTEvgmc3YAEn/FWkDJfcyNLuUs+K1OYGRnh/7UZaYmEX1
QSYY3glh/dz0Sf7J7VJktIzx4yk89z12Kw3GYkAiOEVT+Rpv30/766WScaNanyKyctW+NzRX6dbq
PFjcpOeshTt1gNFTliNZ+G8ISfjdNCST49xEoy0M645rq03Qinm2Nikw7H9ozpiPugef7szEfDQf
Lh+hHO4XvN7//j2n68pRtrbgOKj1g2ekXldF28Ot+FzP/zkcMUt5b24LNekoK9sQH1GAukbg5x90
Dn7aaK2X/WAU91FZ11WcunM3ovjqT46tSCMqDXyEqbtylPzyyhVrbVoGSUnCfBn2aiJIglRRAm9b
D5bbLnSPc4MFO2FhpW0+V8Gi+l/b8tBWtMPYHHYHBmSVUS6vAf1eyz8hMzBARZdRHiPVc2xNCBJn
wPryd8MHisY/96fohcTZEGtvLviPmWO5zapF85sqJIjB4Chlh6s/i8apx9l4ePHT0JLU03G/2kK/
X2WezHyvcGE5hmLyDMkv5uvqEVjcqe6lfTO4Rd1l78P+WBfWeHa0kUMTzPwkCny14oV8656AfYJn
hY43K49keaxdiPQRbcZL7SE9knhFPLJ1WpmVaT2zuW1JVYMXHeKgbcgkxdGDK6VPIE6Mu5kxkxpS
buRlYp5My4WOewp0HBTI8l5inDIU+4iN9nrf4dVLKj+90HPJh7KTX4vW0InFbMMznsdNn8WI+oF/
iUUjzIVyIt+glPVm+G94J47v9bH1oN/4WGSTLQBuiOfXyz21j3/4v9YQQdQMqF5mVtGokAdoPeb6
IG5jkrJnnpjikyXs1+FbPZHA0FyfOipSQIfSxw6UhkFURpiyA3TH5Fn7oI74apBPWR5XG9YRnryM
gdTKgi/LN99cS7otNvhTTjcsfo2mO6nPnhN7j64jjg5q0H0W8b8+cbY2KAavTkYVq3MWP4BAKDBP
+w87TelFmHbsoI7kSuglLeL9/TUQ4udhsjNp/3AOzl8D2CZ+1iYQpFf+7UcTngfYv468hEhOv+YQ
Gk1CQuhPDweFuRcEhe2rMmrn4sPLLC1gD+rWnPdR95QRRZ3NM2lyEVIxHv6ceRS17OccoaAWrhpC
jW5A30Hbu/a+Imofrc+qtiJeUgPMu5Unz1Wq5LXn+hpzcZmXZozskVt4HX3QwPUofnZFiVw9aC0I
jjVSnxCsFX1CgYmykF1obYhgD6AkY5jdAR/1/3gp14YwUfZP30zAohGISiH0SfwznSKmy9DOWSf6
byYY0/ReOpRViVocDSDkVQXE28JlVNhalYaX4rFuIXgUtqd19FDlvHAZTIDEw97PtO6yiOnEm65R
x70T8DqMC4yyAHp6g4K+xdLTDFEQNVr+RDeusYAAg9OJo8kxWxxjqSUAdIItMyoXthYZOxS4sIiE
69N+RkYKy8vDXvRlJAhoGKnmS9kdM87eHn5swten5V9rEItk0dIutpq4w7RVtRDI7EhV3hT3gtb7
y55XRVDAPgTW0PilyPEp04eaxtnLHGJUU2uaes2nhk3bHn3/XlnKESm+oz6HcKG/qcTyPDyl12nI
uPKuXRBF2NweTK9pXf/Eu0KLw6jfD7cEHGi4DSJ5NZhteSEs922HZFjFveggF/GvIGhzTgzzt34f
jRSdKb2CF+Kl1CFle89C7vPQVCLAAouHxQ07WU9TPq+/Pv39GiY+LBYuoKshV+7A+OTpzikxigEl
s9BK4Z8B23LQXHO39dJRHZYDH6pyYibLLBpJKEwQwpTOBIXMcteMPxagK9YtRZdqcYojezBbsip0
A8TuznEHf7xbibc6+sFuohXViP8YWa8OMK4M9ujRxhQDnxQ06/144eN8MVTSnYBj/dML8CqrU7oJ
sV9H8IHgKnYESFmlp2hIJIXnBPwDylO/UXJCSdAMqw8hMKKh9QX2W9UA3AMTACS112+Ym32yNb31
juR46O0S1BJiFdJyj0uIeMimht6EpQ3nmSKU7on1Effa37gs6RhWpxwmRQ9eCrSXe5vOv60Av5YY
lanHDKDZPwCbAiNgmFi6yh2DfRXNtxbX07AbboBytJUvXz05HFqvE/2f6pb4DZ8HXG5DnpzZ6v2Z
zNKCeK6HYVaMaRNrsWQxbPDoJn5N6TvkQicQUPydi8Mbme4RgkiFcJMare/SP7VggJOHc2ETKlUs
XiC8HveBKsWGwH/tjI0MxYAZz3W2FuFm7iIxA+bAYteEri3vyYwPzB+6qoN7uTZuPViFZMi5jiHY
cBLfKDR3suc5qSeI4yn/T+87S4eVQlzfWNjZVxaKNFCCyIdKaSpveSbPbH7BmoXC0BV8+LZpH9Nb
7yaAcLURCUewFUhjUqvXl/QOg4fHvgR1KtIY9ry4cwr0xVodM1/QvrRSac6wVaBcPLXHVDnF8QzN
cbezI2XKJmIBJgPsCIjKIZZGdtheENrn8kuQkDZctZvt3oeE/Y4skN3rmJfW34NwOfCLSuIb0fmr
aPHingLXkCXKObaZfUmAlGCz648FVxsYd6xYPdbqV9Bp8P5A2j6FDaRtold55e208ifumZWIGKKk
GpLsFYt2pt9A/YI86a+/Ld6RQg4x7UTrRhCK6RR/GWI5wvZNQes3AFecfe26IavJ6x3OdslmQ8m9
+0rrp/1G6PqJr92W0Iof1LbS1zLbZ0YUqGvi690IdeKElIbZ7vb98jmCL+e+YwF5O0bVGHhRx4ld
4eAydbLZ1Bp+aQc+N0uijISEgMxobShidoXKUYPO/UH+wYaJasbr8Y0e80yXFlFJ4xjhdmwHusG+
Qc5UFiTjM4LalnjGcqKg186H9mUNgJghjPPpFBfjXUJc2tDc7oQ267g7MC7VliiJUxvZNrp2lpdk
+ZeqFBtJUTctgz5gQw69zL4Rb2a/IQMMxy2pSoHdp5PvMRTIGoMREfOs7dHhUMr54OAPDh9hsVO+
pFBF2RDbuN4GbqH4BaGVANt8lztvqt3TKDAilAh82IAJ+cNbmNQi6Hnw5sm1YPUt4Jrvjp0kxWKG
+yPMyW89xdloMXr6OtIKK4IZdUKVbQOOYtiGVFHREePHKeLNG/Lx3GYYiEYj6+aZxGPS6gEqBldX
VraGf+3sCfS54S84af48JgZlMTecWJ7kP6GNcfaqDU8yEtUBfIFtEkMZPeRi6go52gfLfMTK1V+4
ejSUOMQeS/SWy7PR6xH/2Us1dm/lkKfwQyDvFoGthtLM/+qB/BPYShEepRPk36gDDnne8BQxy+Lp
iPduE54TcaVBjHFAPh5Nny0ySRzW8oRbnYxeumN7rSz36fczfvfLYxO/iru8W0UsiDxGxbMc2h6T
+bGQl2c+dkgDgY14p6u89ZF1r7sWboFbFP8mnUS6LL5mwYobpWg4oRGv0F8p/AiHelxE9ByVt6r+
oh8gYah69GcTphIIMPkcElmCjljm9IeuB6Xtk0kcwDoPNFl4t+j94p3U6d4ZMpl2LCh0YjMh6xJ4
dHdASR4tr7Ox4BkF/kpO+LIaS/tWm8z10YMChObPNZGwRph8SK4eYkMhMyHL2lfGCHGIG069y0ml
guA1qzwktiwc6cEr7aCO3uFroG6PJlIRNLvQCxLFC3N+Pcbtpl8Iysm5GZ3c/+GOJJ72HRwKn+/x
egfaPM6PSz6aEd9TWqGIAsSU3B1UPRKROlY7mdkD66qYWbDp+xVtU2DojVXRoGcnhlS177OO+2fQ
ajssVA3Slj/Sx7lhicJbw2tCQLCAQbhfxi4w0+vBuNjnttE6g+IaDW3YNG3VMsPdxdP6Upw/+bc8
wo//We8hxmcijHrlXqnxx9KKMKULvrJrzMggzPMhBSWFRpGNTNEHrjMxqq3dfZlJxC3U9u5dkE5z
BLzmnZoYrTT0jqj6My4g2BSV2bWRP9MalbFEHQI4UbRS/o3dQwO9Lkn29KqkWSPHYH7wYIbkJtiy
3LHHcgWAQNw+UkbcSNPfPrh3i3OgbRO6haoLewlA3Nr38jh0ufG5ZyQk83a2fkO+C3764RyWBrAy
Mz0d5VWRlLAmriV9VNIDB6uXSa4wMVSAEwhmlYnKvYdrlV9rpSeSs745gxfvFWsV3QrsTZ5BlZoD
Zvd/S6JnO6W4FCthZz+uFF+1Ysc6ADjYup2q7sQOVT15+43ctxvEvFFhRQIqt6RduAXJNNm5l6iN
IslUEWk9TscjBbOWkkShKvpDAtQetuygk3rEomUzG1IqAyFj5lYvosehWo10LiGTdRvSdC9vJSht
YSIvJs7oryxZzgByj9A5m6t6kbyrTT6SMuJU6MFxFphvkLRoE6D+UnRXe+ugvlj7xuNiXsSl1det
qnoClSQmR7qqq3xZzQEmEC1ddjZVJ3v5PM4DI9A6NYgjb+J8rnC3TKpEqT4j9NpDbauiHLNFFSoY
gV4iU6iAQp61ptLj6dNewbqWd/9P/JnTrd8GmEeS61l4zBDrL1X1Kqzl0zwNHQbpEaZ1gNdGi85s
eCDwCyfPK8g7vsTx+CoBovlpsxOlDHEdHpn41OOHbDzS7NH7Nnt6PUMpFtSsV+v0/NcztuqLsJqJ
PumjyOsZlZXWcWkPcETTXkMgy1rV9aVk86PSICEHMCF3Xm4eRAc6Ll8oHHkP6vEFcGUdZYb+aCjl
bHeefAZ7c0be3yiO/i5o9e/2nRNePgHfMGlt4SNLoBq6iNEkb82J+xTcWGveKetoUcQpWfurWC/V
LtVNf58PlKmjZf5qvgg/C1OqMg0gzONAxCL5vHNcj1qnhTR71cHGB5MMVY3SV31vgt62i+TWjmWS
mTOjbCRSeWASFSF6pjvtSDHGf0uA7W2nTp61CLCq4cmpkFO1NvOC3tjW5VwivJFbBfIsvIlw7KHi
iJBp1coTnbE4XUzw3pEi+7og96eWHb30oateyPwbiUG2Wx4EvoBiD0LZKD655CkU2Q0LE4zXYe3Y
iKCbVIdh7Y6+DB0YNyUqqa1cROwYWbJg5gvYyg1lfqrsKuNaq1qzewrbbUE2DPrXqBIo+hjkA5+c
DV9dlxspCW1Xf4pTkrg2cpYxI8MXOsKbv1Ioqli69iZAe3P3ScBubgcYW40KslzFTsQ18Lk8uCrp
eQEFtLQggj0XY/xqu1HwpjcNLLro/MpCNjcuIyJnAr9AbPHcBbAVlrM9mx7AzJ/MhvjWNmexDJfn
xFQGK2DjQW8RsTW24xp7Jy+1du7LxmKDBh6PHfYc5IbsqhoLWzyjSFO6JAqhvaSCwIRrj3MAKcFx
nlBimal6nZ3rKFYHlUyY6V78FWc4jmUh9rTANlloqSshtXtxWQ4k7yehDaptDnR79kdsb/dyUAzF
yq6mmV+/8wLbT/LL5+s1znIWobuU52IZkNaQUkDhVUcBYskIBcBle9j831PhKH2cH35scRv+2eRI
G4/JMmti0nhutWqBAz+FALZKH/G1QHPJXAH15NCZFHnmaLRGaOBMB2QzF+8cnhCFl2/z+LgzHSg3
c2JBFSkeB30kBZvNzynfa4avdrssglyr5MDGlAYjBIXfsWIunZGsNbHVFkC4oXevXM0AEXXRSfYq
eCSjD7w9DDSRuFGQ+evbRtbgJLgifLkFwYBN95D0iZfpm33EsaTggycjEI1hplBMBDv65py89stO
pet6vydt9sO1Okvw93W7RuMJHv4ypc9pr7TGZ7rWgnG5/LLSkHw4H+z1xII8fOGVK1XFju/0q0zQ
UmS/nTvcZfwZSggJg3+DCpnzZbytsFYv5VOb94hVjNP78Olgq03c4wfAJe2fRWViJAEo78oKcQ4F
CwU4svyrizzaXZsJzly0Nse/oba6Q6lYIxtP4mITZiPp42SFpB0Gn9YFPgOjPMySrc8e4+HMq9wQ
Ye/0oMnLTW7qeXU+9Z+ifvmPAhNMkhngFwyeijTkPKC5zZjpRdAcLN/FaUR9+fOI6A+dNOfBTJGh
t8aBUeLBCGv/RLjYWOOq35X36E2PrhNUSWdxe4gXjaQ9dDiXn8dCWZEIJIrJv68GMK6ojiAmFfWO
2fac+0CB/HzZpAEaI+u0qgkW5xlQFXqMW778y2bKReUlU4IH5APIFFvkZSAyHWEwOLq1vzLd9UQy
vSlVGaI3NtPfJe8n+K4oaMXEpgxhyHwljwaXxAtKnzg+kE/a80qXSkHcHUmsoHcX8Y9qxufvIZAB
qCTaOS9Sz2QmvPnzg2bi1HmMsylnq153/zAW7qqfvemHsdwvfr+oCNYyuFn3HxeRqwJdLYlTdap6
6yX0jF4kZo4VD5FMUmQQOwu6M5ZOEo+w3j04xvaskbyb/LK3NIZJ2YyoX88PIG2GEiO60tuJafyJ
auRyZCoP4Ik/CGKIE4JeaNRfMykmzVlXNJuMfwqFFqPQs5NJRtKzNC+tPf31E1wItif1TL6EjsNe
DlC6JCX04y4UHWzMIb4oupG5OK7nhqfpvZb12BRuHlrQltT2CH16v/VgzQYAXEsJpnK13khwNB9a
BQlogFx/u8X0KHDEr40U5zoNckdhVUBKECCQR8PVQ/ToguFKmBw4SjHmq43qerEzWH9uQHxrTMkq
eReT2l19NY4dZpTCOQEKwGWWW74hglrjD42OLrrA69Ny0yN/IM5ToW/Q8gjgWMgfhtCLtnAZEnua
R5UUtjLoc0DsIa0q89eYFC6hHIOZuGUFA3nSe1BTyQZXYbNQSMLfIwWDTp3sOeQ+qcBUaQJ70007
MAbNM0L164vOD8S+DCPhjqfbYppTDaMLQXn4A7nGO+H0QFZuYreyTnHfu9yGtqhJDezIigCapSVU
RifsToVE+RIwBHO+JhkkCJ2c8UVR+3/JIx8HyJXvUtSzZ9GjGcd6BFQQtr0NbJ5FVDM+aBXT792n
M26MVVQYob5a+9ygUalU0wmfDuNrJS9K4QR+uSfbtO5gjG83EMJ7V1eQ3IxqWuqQNJBGzTLieXfV
bak3cw8qXRMeOznKPme989bPFjbC2pYuAp1OXJesrIw1GrsKWqIx9ey2E5RIGE4OGicoMndXo2AM
y3tamROrPDEUCxxkGuUjCSOZTMvJExwY7bEdQa5ZAe+FDHoMIiokuS85FYriinOHxgw1pYbKxIR5
OgLpsU6yMFFxV6j8Du9m1vyoAwaHN9IxAMJtc9lPe7Zx3Bz/IHnBYKsoJfZTsRL6gOYe1aOKm6kC
0NSILXulpGA2QKPnOjlDWznTOsSUckDHrmcWMIyKWqhYj5fubsZ5F+o4WD5M/Lw1LKPglBw8p2dq
mZev7646YQXqGtJDtS0BbBr3zYotcaq7kfTgZXmceS1giP5OTkTagWr8uN1GaQWe9s+yazxCjnFx
wueBV8xgRCVFuD2wI8vswgvBB81sFbffK5C2EJ8rnNuI9airZE6UFQDL2je52EpoealUxbBbBOs3
YmdZiiJatnJ54fXrUGiGeum3KW2dfZnIins9ZE58dWgkyPg3DuAZb/1StE5Rg8bCMxDZl0d/BfLC
4RiD10vNLjACpILE5XCnScIYpOLDRs/BpW/cibzMjr0YVfbE6O8SDwQG6Cmye4Y471tNak8/gDH5
x82nTbF8V8I4Z2EtBxa8tatlH1AHYmiYnP90Sv5Gm2wA8+4S237Ii1a1YBoTklgX0VyBEP/B3ohh
++WdFlxjrxE4qIsgK4pUx5tFcWNOfrQ8sPmCP3tsczO09eh4fKsUbwstlZh/F0aFWNGtAf+Gc/C6
9ih9wlXrTrM7v1+WGBz9XRIRAM817PUILibkyu8KpEEBEMjxE2lwSPbGyGz99xTuyNRVBlo7Bav1
vFw1MezpNqjr9lqwPKU051fvfmEIqUSXIFQqJpsNiRUur+wb12nqn7UB4yykNJagKrJhHR3b8gCj
bRmwOQ31Tk6q0Czg4N9qeb44EuF2mfnG2L0kfZO7MxpFYz8ouSsmg+fVLUwtNzA7eWOUrZq7at+c
AwR6X8oajbjap3kZKcE3Tnj5lZuTNLxfnc2BmKnhScsTd4RzdFCyChb3JBI4BXSIBsbQ3Av/vXpB
ZzHYCBoQU6uwfkUCFBKr0na8u1+pTTbkogwX3gzRv2b5E33mHCsSdpVyTzmdedSfQOy6bfGmMOwo
vc+AxKIN4ajkF5CytXxxXdg1ogDmgacjKMQZR7J3iMI7IVR7M5TfALV+9Au+nfyG00PFT3GjHGCO
QFo/eMk5gh55BwYDiNGsXLmAc6fyYMEfuOWGZ0scMY5jUyC2G3lezz+pIn6pUhf0OAQn1Ld+LAl/
bJxciYoCIqU6QOO5nUM3jXDjd13QHyJ8HIUEFFevy0KTGxyo8e7hNR9gwX+3/l0ghwq6kmws2vb0
zWkXn3fZ1Uh9SiutbBHQVnuswQq5YGpFhM3YO9qVmErAUy1oHJDrscfDKM5OloRKE+znCBoKOfQ3
csEDANA34dWUHW4YysCLZQGbwvnLRW4OGKew4HB5Y2hY8f1H9Gkf5Vi5LnmB28xhWuC9lagdqCAe
dyZKagqt6KVcufY0NNHATds7EM3AJNSVWoSBx/NqbJCbKWqr7Q1vtzM9yczJlLOKEXK0806QkF04
+V4s1P9gDpT0YSLeVOcdafSmIk6a9k2RrIf3RtNh71SFmItG2yYiphAjSlALI3Ib0OolIqZeN15h
VmhDcTTdzvdCwtBEQTt9RI4cJLsHb2P8a3ysgxquR5iylp8rIhPLutMoXOsxbvr/9+npRsb5T+dF
d5iUKzbUTFCJ5DrlxDTpSJSYTBVwz7cLaSA3z3UfkKAi9Z3NOVtJ+KLCsTesqKF0jFnsdborNwyA
nnmqCLRWHgWNCV0qStDABjkHD4IgYXLuvLLv40nQzZQ0CtZ+JdSG9tMpmdEmBsBCA8pInc6ERfWP
hZ/J8++IBHZ18vaeRPAT+ziIBD9FA990Kxe6Fypul8eKFqaFKiJj4IBv/8+3JvJ5zBUMgQcuD+R4
XmspcN1n3tStVUwGUpo8xYRt1oXAIHke/lv1sJZ2gDsTirB5MAFzpMeabC9q0TPHvuXqO7fkoxri
wR4dy6TFYxx7NQNV2tC6ah3wNVbszhknnSm4tuhvm8DP/j7S2TdUL/HCkNvM5dkmqlZA8vSToclw
QX3tKdxKaj3U63ThAk+AdwP0ZQGwYaLvJbd5fCLxg3VdoLJCORObfHOiGRMfGSxije0mqKaaVQ6N
HE0u2qEnmfcUZWG3D58lHOzFC1xIaxm2bediSt5x2rAf511+RKXRiU72IqRZwETgEqo1yYpb/yUR
Nor0ySP92nM6MzOUZz/8QwwuJrwaZR8qGbCnRzLNV4fF4lVpvjNQG0tXy+R4NYDLovNSlHLCWtCH
OeHzbu9jDLZrtFKzmxmRtkuRDb84HpkKcFB4d/UCrkYpUwYwN8eh1eGa5/vM/ExD10Qo/PTosC11
dWgLrwliN5ifwJUZmd+xyDo25k9b5v6y0jtNgHigNCqxBW64SVrXKB7RZX9wHFOWl06Bd3VqEHPk
JZfB8ExhPSndlfhcQrvvpnR4vIyFOrFk1a3AH4WUNy2UpiO+WhPiCcwica7rmWlPtDbbxhjQtGfb
1JoTdkh6jrYx9AyU1luUjjUw/wft6uM8R8V6KkgyNPGTZK4iY8/MNzNFjfmqrMqx0+iEnGx9eVIa
zrzDbF6qB1v5hO1+Zu5jWLEp8lQh+GXpe/SXbPTHbVqn4uwv4qPv/AruwMbd4xyJHsEKIkJQ/iPO
D03p7icqTZszitz8AxLjnVbya4rip6Zzt6c5Xm2D/IazjXUHbJNSt90qgQxHxH7dFMsQkJT4apWx
acmyvA1uM5boeZD04kBNjjJbgqbw3I4em/8FHiI3BmljYUc36uG7jQLjZ3SJ0NsnZVNaKHOo2ZUV
UW5w47D26ccOsXvxsSB4RxlztByNfFH7pl4s+oFKkz3doXWN1+QzXcwpg77l8yxOKtSN0RPmhWJj
B5silJ/Mz5XrkpCsGNyjN9eq7b95y5cVX2lNFJbh0iEfiAoKzuq1SWGGiHCkYGodFBqW6lJrty6m
LldBuI2rfWq2Yvc7VGpONsK6cU0cqtfQsh6reKSl5eAoGqlKxmKDKh1259r40+qEutfilelwzxVp
SI9W5e1Y9CmKo2LnQBEa3g2QoFR9gxEOp4evXyklRvgKgvRVitcgXDUrFjBXVfCBDGJjwRmXQHUc
ZYFCDDngQbEmlnT0xrq89x9lFv6c30Wa5srsU+4OQlCpGrX1SoWN4I71fohmXO0t7bUUIh/5ZRm3
6w2181T2QAgzkLVVN3ycC1qWqMOzgHjQAsuSDh1GX43N+iNa9bD10m4cRJOGLaj//fsGIZDo+6cW
IHqLnytX4TPjJMU8uHYEK0PuPH4pZKXD5m4QviCVSF/LDIFvSeMWllevvv+yMDKD3N+b0N3mU3PA
Yj8ebNrce2+SW1wDS4kqivBl4lH2YT8xkJMcIvxsEyQPahyyD4xcMVmpDU6K4S7h9a6T56JTRoQr
hbu0vWUldp3ORzzPGEv7zmM8JHs+cW3SYjOYaf6UEcAlLwIeZ0NwO8CMKY5KwYSCB65yVqlindYu
wdXQstHbjEt8DHT0EXeC8WlsmgLFv+Ccr0/T8hrTNw0GzjfsowqZxIt6N78pS3oTikzsqRKW2GkG
yajOSND4jJ42I6BN3TMDMr/baJxVTZ3KntXonROUTG6kFHMAR1X6F5JB+noz1zXjo/HJeZV8TqYY
5SZg+0lFgMy5f+UAITnVRAQvEd9d7NjP6NvqqHcYjniahU4J8xKTfChcBTWS4af3utG3nq+QpiXR
MbSqgsI8zVetRal+JdU8QlNBJrtRuZZ7iZqZce2qsetwFunIaxOg8DIFKWFYj5pLiKPOzoov872g
V3TdCOdocJUoKv6EFX043lt6mQr3QLnISU0Dyoq2LnPXwzpHgU+p53WrqkKPZdrZv6qUosT8Iskk
ozmYrvgr5LDI23+K0/H5wDJ/oPcTQLFSeBsIhijER9j5w1sxdrd88QWuPi8AJ2ndgKlIaDEpcbnO
DmDt52kCKTalp7UTzAoWoDXmYciucJMcC7e1gocEgX5x2ijEttEYeLhuV2ZBq97HK5moCAiKktpU
WHJgK9u/mN5kDcwEuTPi/AlRbDiJtr74Ksf/lEXNfaYPleg++ybx2nR0MMSYUdgwCKCk7eu5hFlR
ZhAxQX31NYrsSiQe2zOVfdLOcpj5Pqxy6iRPeQuPNgB4ZD6MJrF6GMaPT327MR1o/wGiwsuhZ6KJ
aYZ9LsDOfrVvAr81Ed2cuiyiwHNenDxDCC8zyXh78PY1oFXH9pwOC2b/6Rk2gr/QWRtwwdUQmxoF
a0lq5qaTgV5wm4tCn4gN05L942vrDiR5KkqL9YEQT7x9fEGL+sYclyUO2OJfrq7GRQcWcGhhNc65
fp3ErUmssvDmdF8Nmo0VCMgL/crp1UsVnlIsO09pDNbMbq/RvAyzVnSjIhtiIIv5e0oRTKym5hkx
pK2LVesRsA7dNIkA5W/wpAVBf9jtxP6vfsf7WgeSZazem9858VS3R0Jj5WQ8fVwYHeDkwr77XYaS
ZplBhUzJ0h4x0xCEMJefxwmvOpVHOkttgc7rri39btYvbXiem2+G8z+/pWhNVjuia8qAeXyED+fU
OrlUhoOyb9DGiUZirq0SzLA3wkwSvJu8M6M7vfM5dSr4/zNlyw5rJv5gTvzLYaCCPC83kxOCp7JU
zfkXjO1ArNykXElwabsy3N2SH7jh4NE8dDNMiifi4p5v3m2GycjYqlPcXDWRFu9AJDuH/ZdHUdGi
Bj86RfLbHDrOZhH42epy8GutSlYsbShLuhIKBhnbi8jxSD/9/Mb+nUt+pPaE7InibQshnYQRWggf
Vx/ewPWR9INe7G3nR10OLXjHQBLrf7azVZYIuMRTiDzJMpIABjKvQDXhBXpFKzJh7W4zOi9+CnbX
t9B6aucr9YoG8Unw7YWqEISBB/7a5Fjodm47BUyBXTixNqrDT63Jykr12oi0SNHh7niUx2FySr2z
lqWXrgbDnWjpt172QOJakvL3pBNFJIbELOSVOz6G4G7/U8OJElPpw/Ywml8zi5L3/1Tf5Ub3gRP+
C5d234eBxVCniMUZ5VoRb5QJLqWMUMqovFKOo5EIp9aUlXfySh11m4KbJ+NvJiTdq5ay6BDgyqJM
fzdXrttBM9Js5nSNq7/aIfnlhVKsqHi3UQAlI3nm1k0SKNVVbNJY8UxYczCPmp5om6KL/XShCPdj
iB0LFjdOMARvlkYoy6pBBHgjHoJTosxZ8Uj7b+jAhMFQa1DT1vKxOpJ6+13TpQ4Op4xhew2b61Rs
qvw/TIQL2Yz8T/E38f88PrCHrqlEdc37y0oHw0EmaqqYNQYSu6kAvF/zrhqXwprc54fxY1T/AA9c
6ZOSXMwOlBVEQTDTWiNjhKQxpb2kuOhdDD6l+XK2KOj8zyrTh1eNx3yTn9deRbzMBEeg8OJ1sPsJ
2m5mderJYWeWpZ0JdD+h1/KmQi9vA3AMvnJ9CBHCwrxjA6jf30rztve21JXayPaj8EFhxZzp3jOF
G1sroioLpxu8HzFo8qv62c9tTiWDzMcrCQL4n6AMKzJhHpgksrHNFqUeMy4M1ekaptkbntJXpqWQ
J0yyEi4eSXt0Gf5pVMzwWluBDoQy+8vwy9FD97nhhjwH+piluNm0jM1JIuC2QPNv63qyEcxHLiNx
Yk3hFUilAUEgMzJMjfQxeeajPlwNvzpExQ+msNN8mBgNJJNKTf+mNW16TglJyNw6QKfO+BlK4Km6
RKeA0y5S6FScxnROxJd0/KowoVDwd6s0abCr4vIpWk1U1/fJWtJ8exd0Fxo10X8h0L61MLuwGJ/k
QsD95wHh6MU5mTCyE7bw2Hr1qKhVt34R2bTr+ammQgdsqlKTQt+FMHgVoSTffShZXWtp9obbQT/h
CkZx+lEaSiO7eFDYl1XdGwbbb5QTS53SGKInuhyVbXaxs8M3crFv7xv+LM0BjT+eZGa0M1vP/Zxo
SjtaI+mHQYJNmr3DTAw0+KA03g2JUP6P8kMmJd3tcFPJIFKUSaPMQ/udmQNMsiNEFEstpe2KAJxr
4GEF6/YfkWiSSr9fozUczMbO7t5c/YvjEHj+Lcm4Xtr9ObJYF1j9y7CgX4gqIEYUwZBNvdZYHT5l
6TdBjFViXge9URtkd88DLn1wKQ2ZEt7RjPecYU7M9klNQ2V6gbn2aM2v/Gm4fmeazfcuhYTA2OFe
TUJ7od9KtNMYKrrB/5/ctIsRwoLUKGtYcRjGJHhSNe/nKgl3JQXj75T1nwoJscq34zqhLgwB9u4J
6wMRkvMQhOhkZ3LXoi3pnoOLhnP26xKS3B4imqHhWG+aZEdjLGVZ0efThgUDdm5NUtjJKvlJDMgn
gW/OY1VBpC3SktUCZCfD6MVYClPn/FdzgzhD3FrntPdEV8jiht7WjgoyRC4+OPIM1ak1RazNIh3B
PN+qP71huiRm5IXQatyuMEhjGyYNJLSVA0IBIZupxOLVVE471LK6au7268uYLqakmHaR7198Ngn6
oOsjhn5hksTyozcgJCI9xoFBiguhFNE/DY/R3aqbdda3FD56bZ+y29okKpaOR7JOemkNETeAJfdj
l0zb6ru8GhQSO4Ss8030NBQcUF8Y7sXLcLFMHO02uMbO2LqWfed9MaUBcF0LfTvvTkfW17fCkiqD
rEhDJKPgW3K36VxdX91KOg3TV0nzwJoA9JHfOci7EleWJzJnqEQPQ1U8FyVmS6znWtukhtRuJR9Y
i4RCj9/5Q29o+pk8IVPeVaHZIMZ8ago/srqKNzHSkDL6EmE7tr3B6vn+9nqXaxxWmgnD5tkXR/3/
jA75PkMP+s5aT6NzBeBTkvVy20x4RZYJUHv+6pVIkyqF/fdNQZN5FClKIbS43gqBm+seCnE/+YlA
wu5F3lORgt3KcgyUeCW38yJvOaFSWaR7R4VDQXbo7v1MAUocPjOGZo3lEXFv91cAZ8fvtveSdO2x
t/H3qYHLNHLJdIJQZy2KYrBLkkaZjhn+y5wpDc2/+FwMhcRrEEn9wZY3kDALkulORCZblmCCNE4R
PUKtHr/nGt3LSuLg+8PZ9lXCxzBvzTHf/8TgTUqrPpFvREessH41TRBsAbVYKxEm70n8F/IKyl2q
UQoQ1xj97v17EsZjw8+GFI0DyFO6QYZTDjHMNsmD7prGg5FO7ZZdJKUYb88x4d6fRdAKeFFMmfUy
1glTCRttAkb1JO7ZeFYAa1wr7DDzjBb72XRFsOjYQJ0EgMDbaAIdeCW0Ct9vwDBIk2OYPWF/h+iC
M7BDjVAdWlX5L3nCSjCRXGQGDG1ZwCB5mBeoTxAQdYzz7MBAn5wIDkfbRoh4V5WBjXSdU2fYUH6P
JROYS/gj6kPwSXx9bfcTjtl+j4J4tVVaxVFCL3jlACdNHTkyI57AwWCTCYdXQ+NJgZ/pveHHZKIo
wzQbQoY47tq4c81nccTs/Ak+s8lLrEE6p/7GuntkFv8gA0jdc3+JHFsV9kk05cbr3cvTvuvYYcNb
Hu1chZdCHg4Kj19d1gmCQcH32DNC3pu9es6o3ipxSvNU9lRxQmP6TRbiyoHE4pl+a8xwDD2C2Eqv
KPgArKiMWkWiigOP1dg5WQDI4VVUgut9lTaxwoXNRQ79B4RSna5V9x2B8TANIGzwQ3gBJ2eT9Aes
457JjXmGGITU+JcVq5Px17Tvzu0yPLWGDqZcJ3pucJfd1ltROpt2D9Ar6QCsHuDIlXaXCgh1ca2D
DBAXt6j5pimusrV/MaiRx+zQw8rh88RyvjJQHHk0TZ4LXvwGsMu49wUcuOm5naRsp9F61/rpah+4
Zp1tN4QsCCyi7fvJ0azLNes7GJkzL6tDOD8FHsTdXqgUNhzLjvevmksRVnocCM2fvj+OTwvpFEYx
UYqzzyNDaeGioFuzsJvOSckHYR4GVb1jqsVCaRZUnOk8evdyWCpcFLxrVknblMeHJQx1h9VoNvcS
oIfEKTl8SQRRfAQPTiJdSbl5R52Z5x9+EVDnHEnGILgM9oMLZjBeFWfnwiJ7rZJvxMV+b7ltXl9U
sf9Emm2BFGcZcOmX8zzvGQLeIDu3QWWkc7/FdH/gMNaBJa3+5f1pQtZtR/+PUEynut4pBi/hbj7e
xvnyRelYHO3Agn109GkER5zaLgwEl+vAcyM22T2w2z2RbDWhwvNtLADOBgxqpkMg1Og/TEXpcF0l
BophbpTiDCQAIQKv1TiBSqF2S1WzqDtvNskjBuAksaMD9sgjG0ZcBJEBfGdwI7dOVxwSYpWQt2eY
DWv6zv0W/c2R6KxZdLGu4J9yAD0QE0495/LnlneAftNdyhF4I/Pk90KMOXzF9s0ntynRYtZz4iSO
/pM06CIhLZW22Bh8MenCMYue85u3WgJeKDc9DmOLNkulVOJRe1SGW0QDHZUJUHQm9NA29QFzaLVY
HbbTV+sgH5UO/8LkkZXRw8bsrvEIpmZ6MSa0y8aDn4zAL8K05Vx0P1EmPGbGocowdJMHDgMtWuO+
3c5eOQQR97DEWBlofiZ8s3NQksFW5l8wPjtIPkymWmjUzem6AN0R1cHJ2KLYfD7GUNM4tPA3IJOZ
wgknnzAewvXTKacl5jQuIvjM1zWNDjhTglfnmauRoukWqCLhyPeKkzRiphLc5Ek8VLP3A85kthvc
Zr/kom2+Pk/t+uwnK2ht19OSH+IyqlDtFKXBdou9ii7LGzttL/bQwNxz9cMu9lg2YBjjl2V2Ssj6
NrnZwIKd/IQuT/BjUmWHYr+LycuFC7nv7SY5W0ELwqMnTXlaYU2PXEA7LKiwviA4XXaFh7Jb4jfX
OAbxocTlaUQ05QeO6mfsGSdsn7yFPDIrDDyqmhTkxMzab8pGLszNELUKFt134QyL/O7HBvMiuK1V
OgZ0M/FluSzjRD3DS4ftRTA/Y/hDX1fWk0a6rGkC7XvERUdcny5O7WPFSLXpw+BRwBmb2RF8g86X
bs2/61z+OohU2fgqvYECOYPuWYkoxfJZi0w7myJ8Wq/z9bpve5jIeynU7KnLbgI+TbO04Fha6RIR
mT3UAJU0sSMVYR2R4Vv1YXPzbxhHNqcrvfH6CgeWGkacwVgQ9bR80tRjCYjgMbbr2KlvaqZnY6wN
k8YhpHf2yJfHQ4d1LBZxyvuoLKaV7FtphQkC41BNQeq5F+opo8ghom2qgAR6N4EikUglsgRfRGM+
1VozMqoKXlZ4zq96FV6z9z1tMVIlsijm4WRCDRmJjNT4f4xmIS9UktfVvBINQ4b+hSrD+EUcb9rz
QndhvHkaTWKJL3rHJ1aTzvDVEv4AaYDyo6qHCrCeAERlhdLlCMptGd3zmNUWGI7YU+eXCtVBjhRD
Sz1vx8JUxmowrgpi05uzSJUp5mByZnlbGV1qlsMVV0wsTnUQlzY83zrfoJ8qxJR0a7jeoqwd0J9+
ON54OIh1myOvULxTatzcM2NPQ/onDQBPB64nCPLF3pxI2oGyGQbAnjxT97W7LP+ONzKlzol/btOM
s+R0teiCQl8SGRZjG//6azdk1USYw1Weiwiqj9P5uwpg79HBkkZdcYjYkPr74FfEtzI/9KfAmaav
iWxpRRO2M7xQ1JdK28RZhh+LmJ5t+nrwiiDumhrm/vvYn7nPi1udVEuHcuoGCY88UdodR1Sgq5WT
qNDHOIb7UzPjX4vRgE6F/AQjquhUdQdEm3EQQDB352ZAGNwCcUDLwvFG/V+QH/918/YZCwUijFSc
O7HWxzdkHe/bGthzER+rmCE57MvaBCyW0m1EowNfCTylTuJDUbXus9L8MK3tveTkSD8zi83EzY7E
RLohs8uEixiMVXvOyblfR1HqkSHlz9Ts8zCMmfVcJDJqf55rkjZYDg3XdXtZqCauhLzIhM2/kp2i
A2jmV2Z+rvsB8Gr46YLznqTxv0kOV/DALvYK309jp7vrVA+CWgpUHYYvD2qtQh7S2W7mdGAR7q0K
eKxzttb3VNxSjCUjd1jb49MjMnO+gxcE6eP06bjajpCqpQKCLH2ugAcTCqMYIqQPezoLkmhRbwAa
FqXQHMFOTYayyV6xc26fgN1j0hrbEvbdvPZuHntrOZy7u6Nfua4uUiVLiXdytzZGBJCk0EQw69zF
YMVCfKv2fLTBrBRblIr2vQS+EbxAifd9LCgqt7vWVJsI85ax5EZ7CVW68ivQaxD/ITw4R0oXoF38
Rbqa7T2j+3Wqx61DrFoVjpiTX9AmKJmXF5SnIgwc3TEYTVdHYIQwqWAabxAYlSQVRxVkBJd6jtBu
Jfe9W8uFv7XAa9ZS5Q+FQI48kdHnEZUZhc5WZgAjRjJbU4fNTD2FoTNlVFmCL9r/ZlaSoSnxBpXK
GN3/NiPCicYLSBKbb3K01J5xBC7+wKflTKf6q033A8fl8oENihCfvFNea2q3Lwx9Wv5fvcJo84ae
h2PCA1aW25AHDniVz5Kq9iJG1n1tWYriJQABH+luAYACK/GZ/xDSY/6uOHp9v4sa+O/DORIjHCqT
rYm7IBsjFdexsanDer/NdWVUx4S6RIuUZqmwahlaLhkV8Lz5UB9RzFZskuCyiH4lMYb7ERQiDfcx
1K7jE+boLLcpgR87UEl3k3K87BLiI++ltWl5wHwwmqmlmSvJRavtiJiXSZWVMXlLfQDBkud7cEPF
8DNqKhZajfmATb3p3DuDXS0HWe0UQqUnZZI/eXmFD2CEuQ30a7TxrHpC11xjaO1l8SiOBcBblFAb
Wrg8CpJzJrgzaIX3oVyZy5niiPLu4bLlfQ07wXbSPoOWZe5EcRy1QRwUlyPjTTvftUqijm6/+Tql
MuEEqhP4SMrmWfBn7Tu2iNXr0ZIa6hjaQeH5EvXm3hT1xAmzjmftgEyCyvHZkB+qFlj6Y0iRgNxb
y/njNuSWSwyQbaV/1BFmd2NqF5C689oKOIHk1A+DBPqOIw7Hc4O2FrQSK6D1RDV+g4flc8YqxQkn
xJdAaMEMg8/KThoyseiC1ga7sucMmRVF7kLiQvtgdxHzS+JmFJhq7rE/QyfO8FSqBO7QnmWwTDw7
59h0ZU4B/SOr1hcf4GqD+k4U/z0i5rH5IwrlniRk852H6F6FY1rEIGipunjRg+/4PwoqY9+YITFt
lBTnNTB8SS0Dc7w94Xxfw7Qzah12UQqzpXQhGdJg5FLp/9CaxYRE98sIdjt1IJHPbUy0pAWV+/+m
tBJ9n4SIN3LvXp4sbCabrIUn+z47aY9o6ArviVBtx/OSmusLMJ1XBfZoEWb/Q0en674hFY9lUZrU
sTzSoW0cYElv9p9DmgNGgeEDUHJhaYlPjCvHdJ9urCZLa+OS2vLsU6Axv0LGA4uO8XBQbrsdCsTd
IiIZPSYfQw7XiRiWPF9oT6pH+wiwjoVlJL0NLtnvpvJg5UnMVtB7SS8gcZNHpnK3Afq5+Db97vgR
lZs7q2Y4SfnctJouunB/MqAVDUn+nOVxGIjxqT6u/9oKGmnzxwQVyBBEo4YsI9fjyucDCj9GvItm
7LmlSNja3Ga9AuDmlnkhpfHqo9rlJ7efRHdcTxwO9bzChTnciZI2IdwaihCL53LdNcU7wW4TqkgL
ZyYroX1kUQZ08AaRF61MS9o4yQWZ/m/GCvLUTD2/ySQgFRr6ZthI+LI/dT6a7FZFJ07Jr3nNSYqH
fyO7St5EsGtOfVGKTQ0o2Fcvfxqh9BgnuSkyMXpLYgrsUTmISgbxEGZjQf3Xi3WvGt2rffIX0SBZ
qIFDBcSTjFeLKby3FEp1thbtrkAyMIVE+sw0Dbk1rp75jaIzw91m19+yMdiB23nUaRwgaljwPYK3
sVYwh5DUAL9DtUba5hy8AjkT02/BYMkR17sdCY3TzMHdYNNFOg4yUAN0y+/ow5TrXmbfNVgYefz4
lt1yc174GfvuTOE5nHzUnmIUrEJrDGaZ2b3v3IUiDhinQW4djZpCMjZ6RXhPcdWlIqgmC6aXIxfQ
qEKZNF2mV6gyON4TIZ7CyUewE5FglZL5op4XpF6SX5KTUoqrVU4OlgpNKk/uWT+E3XE6JIIx1l82
Gp33EzueES3e3SNC/ekP8i1d4Soj1X1n/BkGgt9amJ36wwkvzmpGscdpx/44IYYHhfrfyeFTfeYa
CyhFpoMCHJN1Q0J3YErxq6H8tV9fu3Mrz8LH6PE8j8D52q0ku5HfPz7GiWdv15wWKZ7/SePPer6N
d/eVZARVWZ3ULIOy775Hfnu54dUdTkK+d3Tt/wM+ObB+zUpfbhfVYMpL9M7WKOgRkOupERzzMmeb
rzKBX3II/4eyOFNYLe0fLsGMd12tneJ+XKt9NXtlEhl8lzeRQiGusxA4gb7tk+DR1bpu36JrsGk5
3x0eaWlRL0eY6gVYmbW4MA1YeZy1ikuQN9CNXYYsXXoGUSw1oiI73RntvehyQynCyX5lCZzdlOki
0QGkMKhnHMCqdlbvdRKnGx9L/KfSByqai9dSaAzg1uVsov+SJhY7DzQJq25z/FR3kosYo/dd2h2+
YVyoj91+SHydXDQVo+87dN0eKaQO+iv/fv5amwpY7c1sMDIz7KSRRosj8WEFUXbEAMzkgWR688mS
qkoUlB9WzIVAK0Oqioiw6XFp1A0cb1+M8DA4LKKQ86fyWB4et35F6pRN5RkzmveEeWZmeiqpN1Lh
EsFYTNBdcbRsadYWwDq7JUgkcmIvHe1bHolLWFSiMRzKYBw/EQBPXz62GvkyaECS5YYyrgxobEix
o8UhFi57be1QIqpb/NuLtWDJ9orn7+taEHd/TOI6VUNluCLEzFnGk5bDDu9rIiDp3LNiiyCRnVop
oS/6UxC6W0/iebS4rZophylx17j6CxN+6EThOONnOh3QZAqeRKU2gcnUlqvQFsik7BtdaBnfJDxq
W3gehg234PEciiQgAzB0r0UOzWXkUY3CbdEq+pfTGxz0ZX+sHeXMTC6JtoyLcZW+cLL4LmgS7zWi
boVfZbdAonGTmXqq7RljCzvfNl5ATRAiOp2KJIhpgCR+scrZ7yVIGh1IOJrIEnkCYP/zxBse3G0z
jE3/TfFOqO/4u6rYTPovo7PVDdWiTtQ+2i/kVoAaqWRIins1hpy5akziZ1fgeHK6BZtLBH35h7qM
sKTAxnQkWW4ac9ob3WqQnh0kl5uFUjPmpxIiCXRpVmV74cVqSUPlJbakaL2NZ5NtfYgjAgZOtIgW
sG4b4xpwyHBVUgqBFWp7A6mhzAdqvo8Gh7suRzM/nGK2t5j3J1CEFC48CTt+KpmhE+3drsHpfD7G
Kbkkq7nYnu+xVNeU2cDY3w8I9O8HqujBq46j9NrZv+0NgajT3yteotSG2ii39SLjbvwFxja+whUu
nZX0fyBv067XtTcE0fxcA12joDhIqzxMiiAeKVf+MyeHB9U6/W3qGV90m74duoHIsQXlVHF38fYQ
xd7l9n3Ecfw+yMKepL8LeUpsKlb6HgdXDErGuxPsftTLLO4qkcbeN4QEqCqB628sgZCNqFBQWH7I
btTDfsGCkHzEjwYQvsuwZJtgHeiMUff4HoUhhDKTQvxo9jkO7xYwfIhqZ2k2J4M+YbaDLVVUBIuL
WSOaosnOh8x2CArh3DEFJElE8RWBlf79Ijw+C+h5QL5iXdQaIyhIjIKqbgI8Y+/eGg0CVVhNCUj5
bIhf45g+gAZl+ZpgNfwJJGDLj15BMW3bb/fb85jV0YQJxk9ANZZwPMqiCZYiUdGMdLwM2AO8YM/8
N8z9iu5dRo64J+mMqe9LRIGRKQJNVZPn0FCqP3OjOwHl5cAcQNMZmjdID7PVLwvVbMBi8w+H0KF+
UBSOea+s1uHYiVSY7rEpIIvjh0MKRWha79evaGmTXTF6drlzQBxpyfwmQWsutPRiYRf6g+TOG5lO
15RWb2UyETbxaJwxR/ENbTkqx/4kjPmuzywsQS94ICnMkTqJG14TmS1uN7ksv2K9v569qeSKbwAg
JuBnwm5/AXTcdLx4ySAnYnoEj2Vft1nyl1WSn5rMFMPTapqDw1cNDeQcnWOYYmDzhL/8TqhZna6p
45miDnj9++b/Mqdac8mP82jORFdzMOR8+R4zH/324BK12Kdz2EFtHApBiZwYaftPCFwWgGiwpKqM
GWJ1WSpC4a/Mmya8RrSRGkeMxUNyk3grw65UHsPyVA/LoOC3jQfP8ETGzr7YDMaY0UbINo+GOHmJ
E/XlqHH/c7yChtl6vit+BZ14qhX52zHteGGP63+UWEl/Ur2RKr5DRRyGmGUAWNDX6vFF+c+qvM0O
Ypiu7i8DPGa242AnAnKz1IWVw+P6IVlfNGZ+1kNHGatHsWpWiPPDdz2RAVguUaovqSZW05mgg0Px
F5WJea3nbXIuig27hElXZVso+5cgXBbdraHE+EWkipyEUBRLtjFFbRMpd+LsafzZSYhL68x0AzUO
PtSo9Q1myMJB8EUz6aqGrosxcwobuioJuvU5Dja69C6/azhW9PY3z7M1bXIxGEt9WdsvG5+6IRqI
34WhoiJPdB1bmW0zttAg6cc3biVWI5kF3wSQcMkYCHwS1pVOBl4dqWdJBkP2PFEyjNiovrua3W5b
kSikUjUfV5TIhNUapq2I4sYLpiYouLJkrhGueG61bxiJU7C0zO7Let0XSAYVdLLAyuKMJBz8mLpI
YarztSQcwEQU4j89K1StkG8BPuP6lwNdaiDVIZxkw8e5zhN07yDQul2DLfCwKWTCmyQbhvOebwrE
aqayY5MH88L1uwspvjXfOsp3qRnJF6a01ZWG3mIA3vMOsRbt+o72gCLeM8zNkPiY17u/NCyW1W7k
Wg6oLe99pp5YAr3V1qfg4l+B6xxzNfmHxI1XvdaMWm7PkpmbZi9dg1KLtPjcr0tkMa901qHdsI/a
EcolJQHVQa7gOIwQRPs5VZGR8wR/mSm+L57N0CwK7YRjz9p+gN0U+2EK2S6ula9au+vZofzcwISs
XJLrN76GzbG/KXUHuZWM8XEU25V+o9ChBTKgMxNUGXnXO3jXcEhT0MefUTegHcqkr24PJen5hI4s
3u4OjDzEap/asjDjH3w53vVPh1xOzz16HxLNGqCJ7HZ/8PV/h4EO7QcNcn7xPFWfundH1qUgCuQy
Wzut6ggez+FEN5auW5PuCRBErF7OW/X4OkWIfwc6l23bnjDUvYNjPZDgtZoUIg81xUztLXCoq+fi
jNMmUBLw0SRXEiA2QyUJmbIMswrGDOyoJhh4z1wFy5WLPDqMZ05duRwNvdPrKdtft2FoaFpokeNH
dUTiDJLcoco5uCVyq+t9MOBmueZrMsep/xz09m5TCzpzJjz5SGBPyn/Hkj4n73uU1Ah8mxuX5SE0
qMPO5LeCq74PgxIc0ggFzedqwVHOOevYUcLWVsUqBwCg1PwxpE4PMp2nW3uY1YcMUn5jcfoduYlD
Cte9ygqxtqbrS/QDiHA5hpBHWm6+kMzroF//aYi/y8COTqO8slxfynFhbuWKl2R/mvoKVzKgTIvL
nI8px+jF/Wb0Mjw+y03BNtvpojIDbi/s3BCiKVAbEdKbozXAn7X7DTxkARJyPSwMLs5oT1UhidAH
GQdYfekW4PIh6yRCK/p0UsOLLLKS13MCcH9ZEzbq5ArtwgCaY4eTD/wKdLz1zs3I22dBoV4YD3i4
xmVKrNjVOqnY8sBvDpjNLvzOfiBnGcONqdbvTWy1kgJQ39l7ZZGWQCRlEJTxzg9aQ/xd7fS2rUiM
Am0tXxkyL71ASDUWf9lS7oYrfR/JoRp5dekmjNpG7SK1biNNd+uYGfyuShstGKQ/ZUgBlwGlSuTr
sNGG44xPbU5bSvWaIvK/Dr5dN2E4IbbmZ9/kZCFKAjUTO+Y2+sKzwzqicioUzlVbcTsHfhW8YtlN
0o7yJ5sNDKU1OXHu6y3XXVVIe2lr1d8eFxBQfL2cmvi8Wcs3HeqaKO2/UVvCM2BepAQLt93eg0yY
J1uMT3SZc1ImzDBHWe1CVz3D5ro3/UMXXpMcjYt7CDQi5JprH+Wf+YEg8E+V+T9jSEn5XpWvCig+
fBSfFePUI3mJMej+MCPDPwKkiRw8/o72MiFVF1Uno/ZNxful59YefJYEh5f/JIH0s+hOp0lRC0Ed
PA6mfSL86cmErkxzfOi29TJCYEs7DYY9ztHbcgS6zRl3jAulb3gH4tEhANDlN4PVoo4ebZndHak5
leNbeRZPs3jP8V0cWbY9fTGAjKfN0XNaNLqGtUFOIKsKpROjeLSoWW9HOYBg/q8sn5xLJ3somdLb
b89/5z2Ymustpaj4PY3zuNrArhAjEhB2mm60bbjMPYGXxslj1nTWQeAVL4Bw/AAf3UesXQB8rqp3
LbXdcHkFTIIZuXrqKKlosu4BsrJiecWqMpcy0wFjVcbDmf3VdWiV750S+yZw9eTgZAr0F5IR/DFR
cKLTYRaRNHUyMERpDlLhyTp2VN0LGz+u8hYs+pZg/1qJvaSSrN6eDI1nQ3Ee5bilv/wOSDx5jq8G
8bpYUiGl2AhVS1/FDUcqgpKQWpWBynvMtKW89dHajC3A4eh1xhgCE9LN41jObhjTQmXSosPiMsVm
y7h44pyZ5mhtNY77Aw73NftVA8fV9+zbnGcVjSJ/LDffzPO9+RBqLCXfsLts4LYWPE5NPfQRXAmn
KucLfdQCQOnGvWgQjm3LdFOmtzlKDSDnEaxogVsD/ukHefXqX2zKnaRT3irMeHW2Ldm4cbQKDXkT
Dg/fspI03vq4WkHJyUXLIPPly/2qHhSic8yKzIcml1DDM2oLgPu+indiDFAdhkKJ6zMRQaHokpSL
9jZKkciAS3cAj2sdzMuAZRI/8c8/UHGQQTc+LddTAxQk7Am8Twsy+c72jnAj+zsriaYbKgI2KgEg
yoA8cvxuO/G7ToB7orQ008TWgwQcdrtGNDsEuacjqRtMu7PuSOtX++odHR/Qt5bu5qigpXdkM0DI
UZoWZMLljGaw4oRAbqFYq6Ov6D1+d6Cwz5xv0w9VEgKucbR25w4Xx11qhnpvq2xhyhXumk7I0qi4
xtnbjd/lS2FQiJo/2hhoM7G1oDfZ438/Q14ConCXIJp4elc+w9gP1hEo58hWaGW5IGswNnDupcVf
pYWOdtlrGGYdVIWqw0M7+PWZ8AQEhMI+XcfJTST2R6oHUKkNE10GTP0WB7RnTjzN0rP3OHKxoX4C
1WrB6B7fMC0lxcl1Bbe+345xazzgsMlD4dRDhNxpkv1UpBAQ3YzF1zBulIJ2FZyjFRpD3f1aLK/V
aYWn1x8BRnz5TyQN9AIzAAa7Yv+wO+vFAhN58sUEdVq5ZS1eRmp6ZpvmExU3m5PzVsgxc8MWXP62
W0mLRzGi6Us8SCQPkjhS3nIXTJcYrC1Ct1NEVUnREwwjq9TF4z1zqd/xlz2PUbnjta92aaUtNFJQ
PwfaS9l7/iSfI36AHsQzsQcx40fipWxowkBdsLL4C90VcEgWMDvXnOY21Q2SyzGcQYTJBmbHXKJ2
JndqKQFAB43Db6ZI9ZHjbPAwUXuRhBSk8o95idiI4/8Da1bACfctNLMoJ8xTuwsYO6+tvinENY/9
KcW6NRpYnPm5h62Wm45d7ICcuJ0oyC2RoUWDndTiRId54N+vvvNRF5TxwBwHcK9Kt2rEFX6b+CEu
yyQ6jxRajGfA93mLcriJwrkeM1xBeCsDR61IaNNbkCEPn60lZfo/eJFBhX+vhtUU4VxaFdM47olV
ZJgM7W90ofgk6FNHPJSmoOzjsoasuD6TZIuFuZls5xI42iCN4d3mX3ksfgzV5LLZMrTnDH8EBR5t
r82d5QqKls2/A666nHQ0pVwdde4RYCmC8ZZLz7dVW5cQDdeMs8uEWowwy+thI7xdpqzQiZULd2Im
zHjV7w0TjuC23fANzqXZhYhkkIv78EqEpQk+SlG6MigLuLNwCxVfiZAPcwtJ5RhXxoaxLa/OTwVf
GSGjItpW69W+nRGBJ7wify8e8yU+7qZesaKTzEHLImGvRMFaJGW9Hj+EfGjcPjLATlRJe/845EJ5
7aNBLUjkaTu3jCGpC2kwhljc9sPtS7VFZKcMGdxm1U8u0q4SFYyQU1/v0PzAiCm/U6cXNLqlu1dp
IboIpSKnaOkBAyRv2PITTONM6gVzhpmswjWIlxsgeRGCN4xVXnBqNaHwEiJCgQBMFqK83d7l88cy
7Xx+ZCzmtoHJiKWtH19om1mM9luzACGnN8WUK3J94pzgmCUOC22xhgOc8a8BDVaaBk/8+8T25sO8
UE+eVKJLdu+Juzfy1ZZYUk5SdNMvvR1OZhOU1Y9Ym/Onsu7hyckbNNvndRQ1Fwm/oUT/S03v2i9w
1Ek/C35lzvMoDzle0xnhwkABvBdieFwG3bTmTNonn0kSsaXHihvSmFsvb5nBNW0BZ6bzj9qluZWE
SamOOUgKYNQ3nDFt3AbYsEF3PqpCDWyH31391zVklxbAXTTDcLWfvRLxjZC+iV8arVRbc7ryZr2I
Wd7CCSky0Y8NfSCYX6rTnpsug3h5p2gBTYJZbwzCVQ/WnR1kenTZrFVCMfIf19dtnHYZxwp/pxiS
RGXFoc1t4/thyjX24GCYVwhFNoC6EWdxHfMHtiCiCBmpf6nEhlzdS9DXgXD1a3CrmWQ7efDWUMTG
A+8n/eVTB+1eb9g6IBxHxp9cqWFwcKKQ6KXONCRejTO7iWegkrJiybW18Xf6VHiKwVAfyf1GkN2j
e/VT86U+0jL1prXK1wwFiGuj3x+UWbjo70Q9QxUyW3wlFkpCUCJupX9PtEcfS0LD+1ECncifxvYH
ai7IRh3D9aibw5BeX0zjtaypj+VBgzTaT3E6VNMY3nJCrkWbvKZ7H4iZvYzQMiYcVs60Ofvnve0D
TRa4fLjq9JVJweYr+LPcvBX3TK6L7yy5qJv0Ygc/IPNPIDdwmXVum81RtQRuSDzBboqgFXWsp6IK
5pGSmai68zlPXuziiAObgdTlsln0vulDTM4XVvc6KA0MfNpVkpCD1X9+oEclBudjyKNX7pFyK9pp
EEQgSxYIgIxjjEpLRCGxy/LH8aBocCKs1sC6loaBgBzQsgVK9GwkPYgRRyTOd/JHjZRmGz2Em3IC
aH44GwBLo1BmehvmZJ+idfLbe4r+9L1U5j9ZIUa218F4nYLvlFq7hil/4HESO0bW3KEL1EBd2XG8
MuK7+fK/uZuhsCrUN8OI9CUlCXMiXo7MPf7R4Mhhb2ZSB5V4EIe1rxbdr2k42HBAtGCO4jvwRVxw
KQROpNQccUnmNTEekjRz9e6iwNaa7Etxf4GEmGb/yhI3o3Cz8fv4DFVJdj+7MINw005qC+QaR+XG
U7fq/H/xVaKX9K0hwPzzCKXpKrXLbBjv/cV40RyGvL8PYH0PoCUgQKeCVKaIs5dVSJGBWBiE0rhs
+dx2gagXOVSYncEAduxMQuxWRpuQxIenfGpScOcRasGoN81aW1BVeKpksnbFTgGqnPM4RjqZFkTJ
j4naFrpQSIvJxoZO30MBldVVyD62+p0M6gBugUN78OTBIjNvBUFr524uMBCLPz+D0fY5J3iwAQOW
Pmj8/Vbp03YlBULy4gutTeYvoRpV6rSbjCYEgrScHiq/G+Hzx18h4BSCXLNz7zCbDCASDVR1KRaI
HfAMp3Fb249MRarHk3NR9JzYPxsOyVXFCwumudKTu5gRtqpFUo0Kg4+Oc/f8Qa4MBXa+a5k9HLVg
a6XQqoCz9m5enYzC1JN8PrtkoigB+sRHyJOQ00KfHrV4ZAk8DdhaYkVYG+ZGTSzzPTHkfD8Bs+zk
mfKpq/+mnc6c4vbjwbcZzloCkJRkf6GPSwOkwe3r/rAF/7zcXgSzsgBM4Q5hVA1lAKdZ4eAG6xkN
g6CmrpQSGPFFOPE5DXcXPK9cCcrBxAxxsgJhs1/H0T0F6fPWuMpFZRFSQJThcGsoniJE2aQgrAg0
8RICRzmDrd3q8rqqNQRvaOfAnvEI/7XjZ9jcoC9lRM1z1ba8N6NM923hcrDgzaM7vtJqEF7I6a86
EKNpQ0hQ3jqPtfqAF5QvqvD7HhzKL0iike2m8ughEHxMkHi/L2pOXB7Mg9eFPUkjbsXHhlIdlL5w
bC2w8AdT6sG5tkyq44q0EKpRbWG55/dWFR6p2P7i868to8H+3gg6ZrueoaaOeM98Ps3VBSWL1E2t
ag44OEnPt1aQIu5b7z/YQ5BEigerQbk0feZlVdZOntSI8Q6FlEWmChUBQEtodhpN/2fS205wlbwh
ZlOYFa/5vwaJf20qPJ9bKuId//e8/jBSES09jeYAFPfjnD2esdIpTK0dnmuEHUCyx5uLkWkn6fek
CdXIKTjt7/VFa3cmKeDvQhmb3+9W0HXVW++2MPzOG96Dt9UT8cDYotgvi55dAjhcAHD3dnhdhzxy
OewHvpX2XM1bK9NMRxdeiDbRZEW1/+3S6ea0ITELHEGj3D5BjTi812nLBkDALbzA1LSIzFNT1Oml
5EOER192KVNPpNTOa1gwgGC2vCSGS1e+w1+8S/YixXLnnNT1CTV1fdUW1hZCxhUsO4rh8XL6usnE
n8qMBFXUV4FXXkr2h2vABqmRaTqkiwk0pmPZqiIkmo9yo3HnnPaERXzsynIHv+KsZkYlyl08g1o2
j3Te9rgXc8wF5wydj0qxICdbasgtv6HhdAixImHSk5MMcy3jq4zHgIJ1N5edJE8rwB4dNGlMeTjj
v2c/01GExyipcQLrBqiho218oWah6uCeRgsv9Ck1bx4JJ1RKxBBx5sidSq7XvZW0hUtvI5m2yKaO
bb2Iran5vB6YaLDs8ve6ijjvnq/qbS/oE0EpbGS2Zz1YgsUZhxLAqdAOaWxlMuNmug0DcnH73jcN
kMvcpfXIAZ7+uSvVQxSaKI/fD7zRmgqeQu6Z5PUJWcXZ3yC0IOGwX707f6eELzZr+5tOF7jpSxOX
4Wpgl/q2pTkw/dv8LlaiylvqIQOvoPgGL2UZbnB5dFo1GUZNXOaUzkI5qPZLbZGnPqLJszrX6lWM
TAVl1kK33o75ZuhPMADMHEh3jwqG5f9rMu+imsB3xwvqlWMLnSraia9LQmNGq8wLeTfxjK9OLvYJ
I6oh6eeCSKedmnkbN62qYRueZooUlR3PByWLVOIREJFuJsz/mI3D86omSuHH+aHL7e9Pzq/1qEBO
5mjNqMSqiVMmx4wOph2X9SjBFnDCOAUTxbrJsAV20ztMaLwZW+6Faec0ieLNDrNMTflcTiy7awm9
/MrKMqHl4/LrYzgZ83f5lLa9RnWMvLfp13vblhgL30T0Snykk3Q8NtR3D/oWnCIRs3ZsPIkKtcy4
9CEaeYyt3dWqz3e7u+AqHgWEF3awPiXmstf1y13pWYY0Ad1jkUIGtpdRTtkQf+fqmACCFgebXfSH
ulcCRE7Ekmtwr+1aYxNpChxKaAQqjyxaouhEkNDOfeV6mtHtrq7xVwx5LgWg9V1prpEcS0DRmRgO
ycwrYQtA4msfZloqJQDuo/rjcNwm7lurtuqeZ7f/HrIw2zO21NwGzIgKNCzgPCq1T9lBl0QuOO/E
tk3aNZ/pxPKvZ+f/R8492NkpkrdvXVvVuuKcXCbF0aAgk7laoWxqF0GmQ1hjng3pqKrKWfRv/t5l
nkdOOwgYRkP6dpE1PaBA5WwF4zUPqcLjbBC0LAxkVUTSAzIFwUuDnOtH8uFn+gXm4onJgB7rUigN
iFVXs9IlVmowxBpZQKaPMg24Cj76yqN6MqIZoT3Jv2zgIwwnSuOzjILB+cGlFl/1DTRkkGTarrIJ
FDgWsHK8tGkJczNNuj16LGTcijRU+anEgrING8eYy5MUGSlqTb8zYoUluYTnCnD82rKn6m9hsc/I
WtZKeIyfLte32BpRnh+/oHH4O73EHzeyqLHzpTPMopDke4wR2Gr7UC17iCztdgzZ7Whj/TKmUAfv
0MSMGrGupgg6/O2BPMfRRH5i5HbuJpEOrTpDqWFvIHz5DZozgx+mucgda5nNVYqR3yoq7ykugYTC
UPt9px2GcfHzPYy55X1PnimhJcOsNJI8BEfhW3E4PV/JI7NTmOUhBRMk+8fdw3UWuAYhX16/vtdG
dUAuWG9IHLNxrcSCBFZUOT5YAcssaikMV5OW7yjiw2hu99XJZ7HTWC06HhtyK8EIX5+2eq1ABcw3
e25zbPGITWWdT4mYeLIOaurdlIa+bP3m1nlVzlDvlFIWYPzCgqM/T1IrIoG3QDaHQp/JsIiR9//V
hawvqjDquBvvVKtmdOzv8VyOhep5QGgSbBrUhaJu5nliH4PtF08xo9LuA/7g4VCT7TaSjJigTfGt
/btYiFzlkQUVcyA5zCflHDk9t6zCdHZ6UbFhXhOjR60mQ8aKiwtx9RCL+R10LCjvG6WBhy3UC/6y
aBZYxx3OBaAo05TkDSeA+PnME9SBcEw4IfyQkFOP3fL+8IaZS9rbZdzsR0wBKR/9zoaJkpPlSdBv
BMKqBs/PRB4OKgX9hnUKt0nM1tNn2jjfPUK/P1RNZ1cUUw/ZM228xOm5dVs8Mguhgb1UkGJnE50N
lWCtK5fgRlav/9fyIxISFPTd9wrDg2Y+fWQjdcEo5I7GS2Q58TxwDZ/BMxcQsiJe0MazPHEYM07+
JfyzDkdgSpmXwr5ib1mV/tC58DgS9DPU5HEoMS99WAA2tr8dn/BknefFBSvE2OBV4erUj1c3zg9+
PkCaKxKaFK5wgKyOFHS/rtI7TEPVVD9uJ5Go0OE05WbaF1ySB3+fta567FDhlBFQJsqf/FFiNk7Q
3Xqpuc84NTxoUP2LkPosGs2QTnXOgKD8+u1+h7Yqbnz0JKqqFt3s6yJNXtbfx2Z4XuORpsKOKkkc
lcsp9ZCyRxiP3hrDeob4SHxo1x4jwI97OOcxCosg/FZnRcn8uxayGPzBBNqPpwJX+HUZbAC/mPoW
D5m9mtzefO2Rw0XEAcs72Y3PwF+fq3mClEe8U8AQHn3njajY5imvJRUAcw/I51V5/4RTToTdz1EW
DRajV1tInH2gAPMmkIvAeWDPmvIIacxnR+eDQd9WK2hzUP0ht1hKMOFOZuyWqChwrGJlxUyZfsGd
+spSxLqct1d8gMb+0HpemAwpUdWyfNhiTBa/qoj+7bVaGKKkDPnJeBs6JaVMyZ0j/AI40qc1H+c7
ON+38E+Lg8YiWKNYR8p7OaaBJPNAt5etSa47zu2KhW5XJ6hZx7gQG0BBTQiolr/45Ish72xBwmp2
6R/FYPNMiM/tvAg0QdzPasEO39TpIPo35X6uP3TWYIF1Qnw+FbxTtZP1l9a7gbRTyFkYhYIulHUp
mMvmCETTQzVqYRTFm+2Zo9LtIwaazIJ3eFkFSahgG/n/oxCSnuJMUdF+hnIoAClmY7mzPa3E12dv
NUGZYovkDYl1slQB7MofzATj1l2cOADdHD9UHMWGJL4+fgNPj0Vg+iqnReecLr4WXk8UPPahXlM3
eQyenLcoI1JyQv0WVkCfqJoKrO5eDQEsOTS426Ex4P1my8yJND+07VPOVSnMBdpT3x0NU4zhtCiW
9tfpBsDEj3d3Z/0i1XTX2eTdaLeYwqkjW8s8H6Brq84psmMvGnBqllmuHoSMijoVsDmiTjh/Hvyw
FgpQ0G4lQdUVaxXswOFUkqzcYDBHodGb0RyDbyDbTohe+DlbOvQI15k2ld9O2zMdQuXaAivZkjXO
w4YOyayxJzChgWShvCaMkS/wAGSMmO8GW+2b5C3uy4BZafPgi8pnbaVgAudxzLyb3jM56uk6Z1/q
5qEDQyjd+d+OSZEj/vEePRG9KTgLhEjkfHvqMi/EFOsqHQwgm3dJXRTdvC7ED+pZ/LxDpRN4V5aZ
BNlUEM/8Bc+gG4er6nh1POPa0Dt4QzHjtEJN7fih+g+AZEJZRPCpAJ4HZs3mSOGvJwG5wM5/J4k/
pLUcW00vmbI3wgqqUAKX3y27zzaaHYUhFyssiNrOk99GaE2nKJE3PJo99QukAG6seczNFDBFsdYZ
l199VmtR6TMpcVBhuC8nZk3Dk6XQRHCBdkSxjSGqSLdJ/QUv9OK7/5ERXGVrGl2Iirl60U0f7Yzv
ylCkZjsxtotZqHP8IRHwQkjmsggeY4DxN+z+OFpI4lFk8IRtwq1bYDWWlG3w2yeWqm7U0awoMM5y
qKDPXgGoT9++vHFsmiCMFAiVOknaRtTMNziYuf1MAKZ8vp9WJbXwAI4etDgAEGDtYdnmgcSCPdgN
Fo8nxVeiTm/Yt2qcANv6J/D8nqiOuLRYqmDHhBwSUjqze6TqEG6AslCH1u0mDOPOE+gE7z4NzaLG
aU6FoIfqSO4BZdBOR7/B3dgjumKKn7gZwh4QQPoA9nCtCrkli0smxQk2W7dFCOjCnG9OgYdf8IcR
lPZ6yCenEx5pWxiiu8INMJcydn/mAFKX+CH+TsybqUYob16g8X1aSkqFzcKCcq8CSBBD9lfNImez
CWVrF9L/pVWwrFCo5243OKH8VFter9cYVfDA5gyHpYuhd6DikqXgffuu4bAunL8+m7v5e1R3Na0b
uvw8J00BO/prxnKMIZuzdyfnTasOz8rcP+eaZhy5/CvCeRYs8n00++2wt2rZRSDXY6eVoNZBjcOh
DKvkWrO4pq7TVGWXlMw1eq9IxxnJGw+X1qU/ub6SDIdcc0nNP54ewn+Y1/uyE2++y6QkcCwHk5B1
hZx93fs9HJee+AMa8Zhn9B1DzbpW5LXQ9a3ZugnrDFIR8yQOQZRMfvgzBHEcbrYMD7j6LfYAumvC
FO+fjVguzHkZW5E/GC2QDvzDr5CMfV0WsRQtXVSZQqHd37zjaRkUTyKXd5/h+9poTC9p3f56XH9y
pq05dRbdgGLMOTgveiriW0gY2ZjfDOlOM1XV8OC+rQy3p0dz90FlU3p1CxjwsChB4xH8ANLIana0
VmPEMQ2FRfMNw+gbOFS3bnqDYx2V3khHc4odvoH65s/8gLiBqTgnsuEyaSX7ybZ8u7dKGCEnmP5G
8mMY25uEdwI7FCaINvdKHEaPKU5FRtf7rFSO+glbKbyIHQHnEQOr93P3gDejyzGU91qBfR8P67Xm
iK+rgd6qVGCQUglpuL+R4dEfWrgzHwkgF2ACoO8irx6nOxq6CC73JYaZAaGUH1bV+lS6kIWehXy0
T84wiDV8R/NCcZvXQEBTxQ3v7QNAhpfYJnicxc7PCom6gGTEqZ3T/ONUatHeKjuUw4Dl8z7Iyq5z
tZFlMm9zfAoq553rCfPtaS4BTC2zjD3DTwRLF4fk+Xp0WQKXmWM/kEm58+1tQW/gVHlD7+E+fat9
U/Oe7bak0w/VCoJNDC/34HAwq5BX8hw0whGTPRfuF0jTj/eAGHR1WuqFegUMyz9htpm9n05exWid
/VF0mG/JnIFRHax+rdTm1eFjSmvYyNHXzuUQVhncA4Dvm4QlDQEG3hiqbE0kjknhk922iCfXSSMz
s9nmEhZby44DrfZy6PywapNwp3vZm4UjJjcyO/FzDD1uLcvVG73gouxr1o9XBchxdRhy9MHdhGFB
ieXxZL6noWGvsGFZe0VThyd8E31niJP2y6GB08jmypduYxJgl1hGG/L7fc0fpuy9vtiikte9Pktj
oqqTyocdSYKR4zwWhQrJkbrY3EgLL4c23+DFD0lEcPfA+ED95tjmQEdm2C4CXojbcCLf/Hs9nesQ
Y4WbXDycHYc3CSaN4NIoRmTvsEzmGS6Dwt/CuO0vGOmVXosmyjEtKEvfF71IRq0oqQtQVnelQnin
LGLmfDDtFTuH7LxNb+ATs37mz4FC00ZDe8wmLMk8Eavn/hzT8BVDFvD38Zz61xq1eo2Xj+D8Scxl
n9pDnodj10VvEAmuXgZ3qhFLtyn9c6apQsRt1/w5hoDmxzsqrTed6xE0JLT1aoJyKTh5bw/IBCwJ
v+OuO+Rk479CRPS6J0kzJezAXl/gC+JV3DyoZpXDzmwH9xyjYiGCb60nohTmUS+82S/4Lnnxp7pi
YKmz6EFYt9IPc9bVV8ZjBz649vYh6plC18FpHpJ8+YEKWqSwxPnInaX/uxa1ZDjGRJYr/rsi6poO
Y/Dq63FGjsD8dxPqxydyjsM6FkS2yCRyK/NGzxShWUHb01wgxAXVEpR+kbysc7+KfUdRYdg4acAX
w55CLQE8J3t8fyJuSzxS+UZpSssn1hMdDWI+LYTGyDwry2Z+st8Fyyc6tvvWFUxJeJxv3mAYe77n
TM74PUtNq5Nt28d97xg9EesDy4fGX+LWRxNgt+EkMACBqtptbrugx6JVIqJHnyi5Rjyguioidlhk
s7MtVjga+ZKnPflocSVlHHne/S0dgcvg1NzFdP52CXGSIZiWiX/IWRTZZi1LGnhwV2A2xvLg9pu9
3V3byWmEiYDgVFWNoDHUxTGqxx11s/e/Bg2muy/4f3OpiDfDvfgkIsJVJcBLgRlE4G9uv0V/8QZ4
Nw2DIix5PERasUsmpC937OoaNIN6DJ2QfihAxNXLHvh6hKIEE3byAMyks4KsGyOhXM8jW71fmIdp
0EmJgYGZs8oQH5SUZ/4Vfbzu1lW6VHC4ozWSuGuEfNW1jKs52Zr/1HlNicbSBOHE1m0DkHubbDEh
Lfv67LBvcFeigt7THXdSZbNiBVEFuvtorvTp2HjEsDydAgl3SYm8dcUGZHMpdD2LTZCZZVgrScxJ
B1JAofrIzapOWhc+JOpguOQNy11qWq105TbAtCu8jef9VTO9Li6/C6Vy7Rugz9Xb0bS1Q3VbE7st
TJoJVtZ9Q/IXucbjnrwBtKNEskIXQ/iD1uKsEcHkMXpae0mcdz3ZO3qRhfZIyHS19Iw8yU2d8chy
xnEuZ91HhMvG4mTrY/x2AdNNAA4QBmcM0EN+bWDdrP3T7iCOZgI/iBKRZ7YMs0u4dVypgNnnIOP/
8QG6XOOJP8Ea1MJjvb0TMKeHC8r5O/pG9Oa/BW/wxWnqII+RkB2bhmWVXqQzz4Fr+zSaWnV+BTBw
x5YQH0TpBFjtw5mQaDGwziJAlvA4o3a/VW8a8dWza+t0wPKYnwgTMcNUoVI/WyArsDftiNzeHeFY
m49AE4W/RU2RcNxlgGdDksetjFRqS/yOmZOvex6teURi+FBosFsstHZqhMeGE4Ra4RwfU6FXq1Ng
e76ZkwTe33n3eQDSX4tJBJpjGGvsoUfrLix3UMKtXBxpa20h3A4DLhEN3Db763HmTBTRkOUSMkNP
BdB9AtjHhYYCkvqUFMP2lWQLYNt3OSgLWVqKqbP9/I8WdDSeVSikXdJ7G52DVKTHxngllLImvY3l
vapqObKN3udkznXbHOz2G3bx+VCDb8nWFNzYrO4kY/lQe6sRj7dzYCHDrn6UwkzscdhCS2j8Elm+
tTG4jLyE4gxKwCi4NY7MjZBQMEDwRW8CP99bmz4+Twab2BnRsL3iG/hY5G02YEsZrPaFG4q3ZoYk
eKvrmn9C9ceJ0SCnJIxRUgdmt+JtHjSEuF+H4wciSrAQLu7W/WhwX28O7FMiO3b8sDqdiJtnA6Yv
uJk685joowTWIvOYVk5bmqqDTb60pAed7sunQ+KYDOcxKYHjlloPxVgtp3TYh9k98lke2KzCdoOI
tHtobyaclqfmzU+20JPmQjHaSgirTJNAwMpOTVl+stlUA9qq4qgW/MzdfUMQ+I3ymZBhmhnSYPRs
h4BYeHOsO5il1IIYaSWyEMAjwPKrSc4lHkH4Img7MEl/1/Gs0lWb8TTVM48M0gvHJ5l/qePrSrOB
iuFs9LWa+a+C1UAcolgDNAQXQOo4znPN1T/Cn7VG5YLBTfb9byfYxWU4VE7hZIdm/QoPkzCUcvRw
R6jmgVlVcVMTU36+1GVpUeqTD22y4/1XrhYa2zLgRl7EbpM6onqRMLhdg9sW9/EfggmPIMXc27xC
IGGExrcLEkGTuXFjhmIVHXTDDCZsBDpqKipSeQUjfCeFzv6oItjDs/5vRqdmnGoGNxcUNuV+nmwH
PZvGV5WZF8PRtf2sDGqSHGn97BPLUJ3KlKZPMd5pVEXbU9JtiFp0vRsRfRVYBHXyUqMi58sWzsa+
p90OCNZce32kj/u+vTHlxDbo2dWRhvh541kiO6TUNX3IG8VNJ3t4dNO4xZtVoP7p6hQOmkr0Svbr
1omvP3/YjvhRE+15qgZhjAcrwISVtJmBlNKdmfdFRGcIZliraBYOhzk9toULArgGfad22owNfk09
LwEVKiEe/9PXR4BV6ep8O6dXdd6qhVt0wpNAY1Mv1jHXLpUuF3M1ChPQotl/oFY0PtTnyQebgbBU
hGy7BBSsfofbp3E5OPCgdnDRSt4mtLqXJmxX114zESe3/CpIT31o+MqPmPkMHakv8km2janmOZan
GqLDWo+xGRQfQWfql0RXHkyEbCJvOa5UIVzVwByc98d+5MD1/7X49K0O97xOLzwRrJ6fio4aYWt/
NZ29DNjGrGg33fMImClLF+4D6RgZkqY5fXytfagTyfZ/y+YQEYg8NonkUyK/zU5fUCX8fmu1sE+U
Gl0LSrU5Jy8JJYijfdigGiFTtixifZU3aFDnJ55ha3A1pQTKmoJFdxkwjvz7NZzm5QIX3uxM5+y7
GHkLHav/+AN4UCBrJBzXCL//MJ2hpo6jKdLkwSwuuBGYQR8iiIZDOKy2qS9vc5XOxBuIDFJ8XxPr
t2elu97PMaAOHQvHZkZAWJUGI5KPIPdqWQwSAtktgiML7QwO9yZnnH4vybubC1ZjJa/wsGVnRgie
lug+jtEP9JJ+WkoQXvkt4Q5ENRE2iT7vip5cOVVVCJ/5bwEojaWuVRo2A3QIRTm1awsi0Y7zHzen
KFXkx3zJb4uC/4hGCP0ZT//jF93RsybxGrePD6CMPsyVMp8xnCCeQDrq5K4J4PwiPzrDES8gsElH
Q3A1JvQIwpb4qzj3+ynWSVfdQ4UWdWfvbAdgjwAx/kG75Svx8Po8Ymr1q+pwErbsuk14XNVaRcXv
StFsOZkJ4X3xzquH9jmhywxjMk4xGq3fM63KYlCkoD93Y2X7kKl1Fn+20+iEImGs/Lf1KzzaQc+s
4tZz/PO+jCEc6pggQveOiV0dFYAr9gnwunfhaMFEKTv+EYK3BKb7feTaB+5S9DU+PNVYjeGWBcI1
7V66lgDsxe3x+j2z+3uuMf1vrlzircL3J2fzibhgW0StcZMB5O+aJH3/99e+VzPztwGTlvrUf+zW
KLRmxVpI+a201gpxeBY8BLc4US9q2tRRV4HhWsA2Kz+13LSbBrpscuWlMjBE7yMABIkS3GL5yAyf
0KnYgmth7oGCehgBKkUZUcCrCKlLia3kfXo4+7ohkNsNwHHuOe/hWyZNpE+fRDaIBoVK/Ua/2eAf
Zqiw0VI1s81EUbVy9jbZTt6PCCsAwcUeCCYvmDQ/IaRAyIU3sQk821Ec0Vl+lUQhudZv7lQ5af8u
62VOHzpS+smxAV7Ta9HGNa6n9QPLXoIB/3dSzNas4RK42Apr+u74IML2Sn1iU+qNGCo93uPUlejZ
IrwayluMkURWMNYSefnjcWXACDom/2Ar7B8Ewv5YWaZkxDjqjF7MFeHxA2IC/kQ7yDg+oiGPZIZG
yRJHHr5BwWDy7NmwuOywlKmoA8TklAa+xFwAXAY3w+ldJVSspp0B64i4/Ev6rcRxN44TuZHn5bny
GVUiuBhwUmfs/YLNtqV1+K19zi9BC66Q2ZnVD/c/fYxKxwi/tBkekZKPfa4V9LODHmzRm1F7l5Wi
4+M953Rgz2Mhp4gZvWbcP5KTD0ccCIvEpU44QbDazaRTx4e0M6kfUPV0nnGAMy5RdYeKDK7FJE8d
8btQ5aYOsRauYkunl3saAwaqpDshGRZ/glfzeKuUMP+wvk6T22yeQDraz9rHpJgUGn8PxXnWjk1w
ZJn1CkxudMYY/krlcWZUz1TEGbX2ngmAF1e7srZV1qtPDCXAe5DW6LjkRaGH7R00/syIbAkwiYKY
fWwuRs6mSX7z0LpbvAQBDDRNJuHSqTMij9gsXrkNz3TvBXQcFCa14Fq7vqSqCys4X8vZaQrPPkho
CPquWeAJV/xqnxBBd9bUt60undl/o+FwoobvQyulZN3UPXThpwTfz5n8r5i9qVP6UAa0vkm57b0t
Uez25hspBDRNx2U7TbhT3JPQIjU3zokRhw9/xez+lgFAGxjea2Id5Krjk7gsuqPlb4VBS9JstudM
XJhst4KH9UljkdQQXx6IrM4+XUrvjaJK3s5idtUJvseS34Uph5PFbYuxlPtjhXFAa8SbPK7V6Pn1
i5quEjhnRovOJs1ksJ9hjyMy828jqeofiYxS4o0qSn1gTgW0d0CexUeNfVhOnKjdHYf+xKym9TKi
Yx8F/hSB2ltnhOWaBO4LIQDPiAQN3p9qBpFjpG51Pqr55lJqYUi2UuAZEEXcm0MFk9ggoHpOAGea
m8eOGs4wwLwpwKTusK7yeAy3/MFrmpnOr4N6q//rlwTlvTwxB0MTN35Oj5CGN6DFuyOznCK4nMzJ
qKSMf/n+XxEOStAv9RL9XwCxjYyoiE14V4osWdnLYf9myFnfBRvkFyS5+HYVDsDYiVth3+n6LrHy
o6C/8vigSME40iUoPo40OX5QE44nZLIgdiPgJGISI7sHSrpSmAwx6HJrI6JELfJ/Wc+rbtizL288
riZDZhCCcdhYI5KZdJK4cSheJxxLhxUj/y4sp7NYEroIsbedTp9Egle5J8PS1u+2yfl4ug/6G4jt
Q0jZBLrBiEDlum/30kNRmI+TWVSWKkexN7yfn5+5F4MldFxIrUUPvIukQ6q+xWVUa0YUDlRM4iX6
kR+ixR5qVio2w39PAVtkr61INavgxoAxe9clPEPSJquqZhj2fcrUMik2+8HjK2edRpne30IOXXMM
IutvDYuXnIH6fnwkC6h1RabQppcTwG4NiFWDEqX+RBGraswGoN6W9S5PI7v4Kj77k9WCIDWkiqrx
tDih0nW+imAlpIsEk9G0afc4/aT1yJor6vjjU0Sq86ZVRA2A2TCmUUbv0Xwe4ZNPdvv86VRrYWjI
37DqOHsac8qxwivXDOkmu42wY4hvWEEVdHlemaqtxZvHIDuoB3C3CF82+h7KGXnDKLxX6nKbvh48
gFCXl5Lz2re0L8xnP702VpkreMcjH0Cy8aSox045MsusY+QsSHDUqXS52y3tZVSjt58EMVDbdNsW
ZfONagtIAU7PL3Bl9v5yP8PFCycd91BKm45i1Sx7nYywLlar3D1wg3LiX/nbJk8sdZJ+SmIS0fHj
rW0xOyK8XXvphTjqlXCgb5zEjlTOWC/jAE99ZE3n4ZZ0/QLRjA5qQwGzWB3LZNYDxeEsV2f1u8k0
DXrndzqAPyBAkDn2U2flRpn/VqH0ve+GeJz0EObOfb+dpOAUdIzzUY/J2wQYIF9aHHD52ecXSwHd
mpmzvM7m9tI7YMEg2C5GQEAsWy1SXQ08jydByoW5rsryJtoUtYNIOcPHWKviDvmsfAiwjaW8Zciw
cL9vB6Idw1P3lABPZ3xT2JrPzWQTJLiPgbkhKKMPk94erh1XXWhiYbltGJQAgr8fUEGsJ2yUhGQW
U6JcQ5CCUJL7zo/IWHxoOpcetnflVdG/2DkcpXwoc/5xf7R7SKtyaq+/pH7tCV/hPIdYiksXAJFg
Z2bw+D7zTiGErAdtt7ln31IrK3GS2seaGGmxDlrSvtGLKQYyJCPh2Yg4zanq77GW1riyAcGmx+C4
oRKHZBbNIDrdR0grNeURj/sMpO9/3wobg0gEgS4HhjiybxZjd4ozc1wJl56G6vbYN6MbO/2gDi9Q
Im12RJVmbg7SyG/E8hxSIIpPWDFtzOu8flYB8XZrh3NsHkrwtvnCiD9x2NaQaKSbAYmy3P5qKo2t
0pR2+fFFChrxAz/pKoC6tMFHnxu9EKv0wjxeECO/4xsfOHrmjw6Q6LFx2zY4L6DzxDoXUUd57mop
y62Fwng0JvjLYNyva1BQ57FoTK0XWF+Eq6f+sfx3Po8H5xNyF2GGPVa2/yI9qebfbb6hGBEVSb1R
1Qx/Oq8nlvqSV8gb8QMj40ry50hcy7I/47tr3YBKown3yzQYvFu7vDnRMaIQ9w99krTmYBAzHI9o
aif/ehV/ohKRyjZQpPO63R2VtliKClBa3uIU2oPHLVRmmn47gX4cYdIrr1p00nOr7mVnJGsf8OWx
ltXYBcNqO6cMl6FDXMOXDgTf5i5b83vTLxlg7ULUpvYYO2A/L15WQS6I2MCstytzzzBbwRer9coC
mMcTRe+M64hCMsChO+6zUcx19Ocbob3loRpou7oE3zknb3VaZKdoa+9M1UckAGTJuRlg9WRX5f2D
qZ2UbV1kl6MP31YM3BSh+D0XiWq4drYnLcpuZFPDC414L1Gwq52AtXNj5F0f+zQYERU86swR0Thx
lvJLL1Ivofo2Q9+NSbWOyuJVLq700w8X5NHUIPtbJZzu9HzbTiZQIG4LeoAj+SfwLkjpjA/M60Ao
woeJXSyulgF1VXE3WM42tr2yvHCuZL4yfEQ9vLZk7qXNXTXZII3fBVynAdiGCxMEw2bNj/VFUs02
n4Bi3FFH5AhRcfwU5ioJTf2wjtycGd1X2097fhjXtSmzaXCrNG3V0X5rZl6/m09M33kYGJR5vzZj
pl8DieJINY0SS09og1AiT7IFfSD4TAyYmQyl2vurIoMGom0DIjjrPQke0Zy2/Qy2c00o/1uKixD+
e0LY11Z0IsDfluRBlunYyHy4xNeVDq422ng6VjzL9/80Eyzxrh1ABPqT5KONwv8k/FgqeMpRst/m
aHMOeYjJxJ50sXIGGRiBP8wMBke/38ESyUWKy3e+sRGQieUtpHRdSqAic3gL85lEFDp9N+Zpmj+m
0m3B8493GHPPlYNSKGcgx45BiOtxM2ZY6p8PYyf5wXbkkjyn3RPOWcpBgqSD9t2OVR0LeYUGaUYe
Xh/P4jNgMqRLPmwM40lWY61v9U26Vq7S7s7BclnL9nc5Cr9pgvnwWIJ6w68g0eZCGj2tWxFkRnDH
93zCebUuk4YkUSXdq5HNyVQ7fiwhX4XMC0XxLerM8P5EM4KJSTciq0U/DuH5Clnt4Jkvq4FHVlm5
rGqQJjn/gehGjdUTBZEn8XAd1cHoGqIhk46iJiDSpuwOXpLiQzaTL13djgnI+b33OnmsqFEJrY+g
uFX5+DBLr/X0Og8cNirRq8r6IwPLkHoL1PPDaEsd6kvuH1CnTKRPUaGKa+1+ChOTt0H567eplqUL
J3ZbsvIU994U/0KH0E32p0tvDtVPkmm8O9+xCuGuuRDqdJY5gp0wyCnKG60atN3jyaWbWMK1q537
40j8uoCVbu3qiVuhezn0BLACZN2kVHCxA3TxkL79To1fjFQbw591GOcfUzQVinor+NpTPxfrdpJN
M/mNGYQ0AxANUCmLph9ucE1Mr29XKF5wRaudQwjfzdpDXQPt9WEA0MARgSOCHpxY5jroBU5FlUPZ
9NUMS4RFuIaqSUQmIiEop0hnNN8HpkxwCMWb6S9gWP2PJrIULgHOuXEUfVM591sP1lZSHmiMbGDU
jMnjk6yB+zfmaGwpuadft3FxSLVVU9bVkJuzmqQJnD65yrwMjFyfo59p+pjPVUs4qWeFu5moh/F9
ymdly+fGM2QkLOY+inz2PZ/xwqrBy23984+xHfVc8Pq/JBi6LB4jhlfRY3+AIKB74LE9Ty8ahanr
4r/tuadhqAWP58sVzkOlHI0M5shoAavWX8epOBta3ZOhpXkaC5jIH5VHchFwGI2O03qkAwlizt8i
5241JwK0UM477QTmhSrqM9hxjYRApy46jeFdJN/Ssyw0LQz3UuMpJ095hHvtMHVpDfwkT+BfKjIm
rMqD8mGSNeEy8bIz4bVzIqgWKSZ6ROyvyXo5KwzrGI2QXZ/CTHnX5/gWBvgs2ZPeLLHix2J6Bkdq
j0WMKC50Bmwo2n1rVKtcv4KK3GxA7XGHdPAA8Mc0kbNdJ3LGOtyAmCTFhJytlYJTGkD4mUB5v+M8
xraPRsTLbSdedYYzaU1A+uy1Nlf7JxLR1bdVgZMrfCisFbmy9Hc0qfAn1qDAHBxc4alS3Nd21Hr3
C8J2nUbmb/gH3tUfE/Ss3M9kz46NzkJlU8SaU/kHhu6IFpchxzQKEvRkzS8a4uFkliDmGqiXvHIC
0EeiTGe7pZvPmgAkqYcHRHLTDHW6A33fSxQ57KBtM8PnB2b/tidh8yUmvQUb5qmjHYlQYvmDtkc4
UG6Wo8FGaDJtHRcBB9FuUwO95ZulCiYOV14wDLI39Oo7v9JEjDQvAqT2KEzheUt1P7sdwqoZ5Kaa
NDWPyVMTbmHW5UTux+wdJMYBYppaiH8pZ3NyTrJ3IPEL2ofO23zNb5tu00sV94zpxt/j06nZaU3J
HRszenWFyWBKbycP2E5fvNC5mx6ha7eYZyPQy4EDKsUZopZYydv1jCuvxB9/YlL3c5z4PK2WJcFu
Cv8phEZNP7Gzq72LTRLihEv9nx+ombTET0mopXD4gHIFecbMINHU/M2M4437izuSL5eTxDWU7FPM
EPTGs9FIQMYiIhi5Do2EweFEnpqP4egYGHmlzr81kV8uS07gpTNCME2uooK450zJ0/pNLlx0jBzT
W0bhpk+yKknxqIepXjLp9inrTQrJsrGLtNRKB3g52aMeULjualQrbRCkxng4FslYc5WmCB2602bX
ffomYIwQQsPfxOTKmMY3hcEGxoeYZnMZaIk07Bcj+RnQGtcYHvva3A4WrJBUUmaEU6S+X/KBVEtA
mbghOKXmc2xnlE00AzrB74zvn9/VVx15QWE6Y/arvu7WkhgwFK6YeULgBi+64jSR3rBcaocsRIcY
DNwA4/rB6HmwemShlc5RD1Cbbk8N/PFOhTBa+Q6FXCRq7/N7t5MCD0T2pnsxJ3nU4PMWWkOm3W4P
6mbpYza9A5g2run4I0iVG+o1mXLCPJ3Pw110eCyJdUmfNdpXuL9oTXctZo+Qa/Uwb7ZFN7mVt78A
LmOVBvKDPDm8foPUmUOgjctR/qCGc8XGySo31giuGxZxE8x1oFMd5o9vhDfnqUJ0hCTMN/RrkqYT
P47RhNlAq384yvv9b1V8amGOLnq6KRP6eOYdNfkAiXp83yeiRItn1UFOMWSfK6T0a6A0M9sN3YK8
bR2lIIUUuD3HoAxykn+nt0nuOTUg+g4D+oB6dhJDoVSmS0In0kv0rYxLat2i1aygrewzvS/nk5mc
+Luea2aVTq2oAuRFuhC1ez+zIXBa10QRoGo+B9hx1yEl19KQDxtHAfbd3+3NkRa7e1kYJMW/hZzR
nos3F7gZxZY02DXV/0VZsNf2N3ZNE90RnlL5MFWcatC4639rUyeasKbouNjS4myKxz8/Bh7trX9l
z3YSnNAxqc53KDDE66xzeOzbgr40MfnDePWKxZe2HO8n/GqQZDm5RCGNdzwu507MXCwIzTFByS+t
5lQMlJiRvk6m2Boor45uz3vBtiOSBgkMrFq9upOkAhJ9U3l9+69SPPN8Wu6mw7op7NlsRjRpTc7e
UuTb7Y0cadfIlLCNtdHIQsO9f4b3q5OJ/9gDAk9RXImPuTcsoYWax0hY9+O36DRHJIB9WIOtwg+z
IYqnNEqQla4PSIY2iujWLwS43TD/WEy6hqENjr176ibuaryShMsU0jNSj4PI+9Erna0HuwP8y/X8
5AUlKdm4giZlQo8r8kz3PaYQ850rXdMFohNYmv6H5m5ZMrmjrtEDC9elQI9PyuZ/K8slSORXwU/7
ooQXj+FxaaTN6xKBnsz9NJSpRVJgrxarCWCHs/Xql3hKZx9vID0J95I9LyfHVq6gErzWn8Quoz0v
+6+Fn2nLv22SOFzdX54m777MLbT2iq0mM/ojeHEQ2nq/ykUy/fgnWSvBsN+5Zyjt4z+BhfAhEBG0
m/iCUFHD1pfTs5x9CKfTTS6PB9w3vmJpqDXzB4ZCZV3/COMYBj66Lx/WW+oGX/JOoy+01esYyyGw
5XpbVlxn47TEV9stEOBWpINlNq5Ptbk2KU3O+0Zs2Q7n4AOtlUACU69jsY0VhwxOCcrmuursETCF
kBPcnVcGXNcQWNPYebLLVMiokTGlxCDRJf6VoFI0jHiQ5kHrEDZPJlrvXmqvaa9DcK2YHYBpChzB
sYIM8tMnpSJQLsdLls8jlYqGLY17KfM9kVz0q/5sAJiduhTvrUXjD6cuHvhlW7mxaEFtscwVRiBd
LorgD1P99VQqmQ75lxfnSbRC/EbEd1nRhpJfjzokHGG3tA/Mjw1u3OIK82XoSkZXVNDoGPwiOPmT
BT4+2PWMjCbaNB9bMB4CNMknNhd1fp1yZ443cGzECULtJhKhZ2KVaT2f54V/RcgnHvEF1B3K8+ji
KjYYfxBDSVG9xsViyBl1TQye1LH5xyo6A2rLeogH8pESKvz1XapYFzImi4HnfSJZK7Oda8ZCEGtX
HMVjMf5qLh8UXODQvimCt4+zPOcVwuUDvViLrrPVwYsIvciGMIxx6796pi88yMUxpRuSPQkUtmL2
vJyM8vohcPEzCP6xXzJ8ExLRMh9yn9gzSowhAJumA7C57hJz/NQdIiQN0WElD82Bkj/RjgI1lmWH
NG+KZI2ob4JBulbo0N1BktTywC4u+L6+q0VF0g6+ikiyTy4Dzw00nBVKJxtbbuJYm4bTgRxa0gIw
4IT+l6hCNkOzzX5vZ+TqGar2tBpKaIoxif9e3CMb35tFEz926D030jbcwqupQg+qiiZPBAODnUg/
dRa/RHcNjwBqBppg3ji+ibFluOtM2BDQVPm+kcPr3Ag9xQUHJayhDgDbr4F82CSNyffa0xiz6snH
DaDBfR2LCZyXB1QtU4nBbwcNqOZxZhUL8YzWimgiSfcIuFIdCDqtreKyLWNzyvzLyQ4PYo1Z40ao
MS4rz8A40jOND0+bTdzsTUcG818eehm0v0KkPNCYApSGwD8u1W4svCA8wk1MCAliuYoFLJdGgGng
4cOGpilGdQef5GSelUhl1hjeeNnTxU6HOW851YKvrtH/HhTYFnYRE0/TTCGrh7i7PakAjJmjiSeO
pLADbcE3BCB5yL8DW1QHW+NETY1BxNWl2fVRv2VVVouYb5NNfZneb8BY5v49h7bfrvqUAk/3TpYd
c7Tv2ygRSQ7HCQ9r34d0Xej6ZsoeWn9cnsVupUmSD8mI3NHBckASj7c+eYEPOGY9NO6ujXOdI9rV
KVQ89/XY1wues7G/gx09SaAvQHqyd4tJExKWqzfKBNupy33gQrtE+aLS9Q9REv0XQwjmA5Yy3Zll
knVc7BDyCkho/LkvcQHDFOUhQ6dhBzNfenR7f+gScYtGthAePKqhx3ZWPDnFmCUFPhxfn/zNJF28
swgSNAWm/iiwMeX3j54P927iUTeRDypYkz5UuQPpRLOa6CJqjQSGW92Xg4n5oY6oPgu7+ihRVVNC
lNj6eWdY9ZmY2Zr+XyHYGOOBZKBPUJRMEiSCk2FjYZH+MYlagTQKAczy3AQAYj+ZwtOzUdG5vQvg
s4D/KxaA7yJgPHIbgYuIwkKEI61yUQEEvZr0iTsSesmGxs1AIHKpKMtPTm6t/ZHHp/H1b5qvCzi4
SWpUfbtfLKF8nzw+PsaX1gqG7nBU6jHEcLTmlSu1w5a8BMvWLWdcgM51y5jJYsBq29CeC9PpqZ1Q
94Bp+2ELHF8tc0RSflnU9y4BsfPZZiV/Zt0hJz0uckBGPprmaivEa0Hufjh9oLMaxBVr6tdIlyMb
cggYvsYq5YE/WhdCC/kTzQIinbO797AuwiPIX1VYcPp1RJoXX9mVJ4i/6DJHOfHTmtC1ENec436c
AwwyOungMOHW4IfTAFCz10hYOlcbTV6TVMBxc245krZybGrmjsZ0SRcmpbs2PwtIUWTfPYK/yuUR
+r6W6sW7yE8TwjNP9W2nzuLK8CBnD6gYaAiYfEY1JKKCyZXt+jhBOJf9cjH83ooVs8xmSKNJehMn
gU5Ws3p/mYCjIcsAevFG6smfYf3u6dXF47WiZ/D+Gy+DDHkYirFPqgpHSBYvwBTJCnem2mEkyIkP
Z7LbcV1p+OT8zkcaAvxqD27NviIRvANh8OdXa8dv9k1Jv8TfEYui9eSP5CBjJuZVmXBJ0nryvo2R
kWkgj/p7g49eazKlqfnAnAfPvT5z11LMorkxoC0ueWR6FjPIU3uY5idvuZN3ZcizPnVVN5qvLpB9
8Vf8mD0GZ1L2prxEhEqqHDKrEuUFVDix2ZEg31vvqGCA9KMQZmwaz2BNgr1h3LR4nVMrlrm5wxW7
yRVSTT7G4lNVwdC4QNp64iQqq1sR/3N2ntY/hx3364FI2pgUtPT/dSbSpUAmNJ61eFbWeL939lPb
wZsP/5p8VFocEYnLK8N+eOuIGNc9mPMGEIbWq0mVR3Cl0Mqwji6suD0OTf7S7PSgT67ElIDvxu1D
13qnCHhXQkZwKJSuN48MeRISmd1oOGUL4n19LSmsw/A+g9b7OMhqKnKkDcK8dXrwYQ1UiDPlvvU3
Wf1qcnSC0jUZ9wWsn8eEiEuWvUAeNAMRW/zaIVcS58hFweAb7mvQNjf7W5Al1M1cgUsb6AAdcKHV
21/iFZ75ui7LTA+RcInhsT6sndxgQbzNR7VkL8Ja0x+JE6rApsAepiwW5rm1CpGOvbnf93sNpnYu
0tgi0MefFNvW401dpK9lkcCAdn6lNNTrDxK7g/qyLe1/+U6CfWiAeidE0C+MUot54ACTPEKGyPi+
elsoebC9RpqnXfllRsI8JHpQIrvw9DALkBfvk5nwPvZi+ffnG7p5gxiwCN+d5BE9/UU1uztaWCgE
sVrqk0Ng5E7m8CiuZX0hqCD6LX/NkabrjpYAUDSCk+nBkgthcLmgZpXI9yxtmiagzWn+9RK9rzOL
VvaieV4hXSDYeQVHbuH0SksE2xj7kMhZZUqVcdxaOiSZY4rH29kfJkC6MUmBJ9Aa6KH3Zlnui70v
6zmm2L9wTP5yrQaVmuFWkDBsiTVvyVgJ7NCuEpwd9C+RoEZPeZ1Xn2gYplit8gBWOcIhWjIu6IoA
n05xrNdKREM/LdUerXcU7LA3cBhkvutDPvERH1TKs+PfCWkck+ODK+zR5//LE3zx8YTPP+QdY8gT
ggzIgypnScrpuNLk8HC0y1nAU34sFYBgrL4+kf0WtK8eTZ9ZivWD+BCk9VRZx3BcoiA9GfXJ4vK8
MPkdnhgOlreA/bVSmuScVK9i6w4yoS/+btRcFlxcgTNAl+j8rytUEuALweNXSw1E8vRizNf/Xgam
J2+RUN/lYZXY+cTINr504oNmk/cPzgwRp6J8KqfUEd0i4MSGd8Rl9X07PCFTm1ez8LMbEubpUmeP
CC9dGaQX891c24TvR/mmGr4FfO2+QgKwZYEOmEE++p8LaN/E/kQ5YXJhJIKnMBjwTyB3O9zidFQd
DJ6JWl3QbUN/haaijip6ruAHeERPuGqIm9lZ9tKYpLbzQf+IUf90+l2Ei7UJ/4u8krAkqXH/xZfp
dSzEWXKJ5RdMhCPIG6wNGmEWMh7Ohg7kUOXPlX5vshjv0hn1siCJfWvZJ9aHG5zY250nT2cspXcH
7WQ1sw906RKHaLTk5ydPD0ghJenC+WZ7euqipBbW0Z3VWamUWbe7py2SkRMQzDqiNHmWEgr2d29d
+w0stYVHFnY3Z8wvRh0bJoYZeDJR7ct8kcKMam2aW1UCJj3NHAEe7LPckARZoBcz9Q8EX/H5tr4G
6pqs08D6nuvoi/rDl3tWq/HPtsT/QuQgPBUikP3xbCLv4OCC99Uoiu8iSEGU5p6lh76nerOdvKTv
YxySTyeFATaulrT8UhuHLOllGmE8ZL9AUB4Bv2qH8GWICPNrixSMSzz51ThuhclLCwyKEgpjT4HL
2rMJQDcz5bSxA5HEdAOoPuc/vJARJ0520B7rJVh7OC5lj7vXzYIBuyFLvQnQkLbfCLlUTjPP4gKg
XQG4lYY8X+g3Vpj7b7YO/H9KtLPBFx2zqpH4PLkR2uERt8nBjCpYcrnX6SOTDbM0Msc4SP9uK6kM
sGZqxUL4Ti4gD8Ikwi4pFX7/ge9O7Ql92aYwe3LftZktgAHTkO6u44hA2QpM1Q2STgeiUXYbimCH
Eo0LFZyLgyyzc2buVhOIA37cqOk6/ztpAU+nGHHcpAYKDS355kiFyvExHVgFwwOZQmJQJ+Dx/x7x
ZDAxAGw4vwOGN4biBznlf5hmXYkAffrxKIh+d4b6+VBNxAbu0jl+hSo9KNM7gM3Yd+iA4q+ZDdlj
8BvK2kK3nE/uc+HGJB6lDeXmn+6xH6y/Xn/adnOFA7MBzrlhIqNm3FPa95Ak5aNKtAABqxcYavcU
xi3JeYN2UQPs7yrFEkRZVou9y55jqjSSSFLObylpi6XsDB/XMB35rJ9C0IsqiZMqmAOgSWubHmlI
apt/LR4xTW/KAVx+ZpI8De0VqxqZcFVZtm8u8EGFAUDeTYZZFWLIuAbWQQNRAd1RhwuEEjfxz8Qj
6llDBS2iwRBgBICKmWjBK6OiU2pPFq0KI9CA4MhGyTpV5BYU0ehRolb7FhgE3SYwa5CqAo5INpcT
znelMtwZWBJdy/pDjSu5/IWlhR7qbr1+L53FioitBFLK5WAlE6iyytncSNxD83r9iasB4BlVeFK3
GGpjwArz0tlW2gjP7fdDt/gIomkIIlgoNAKO/+mp6mItxFnDGgohfnlkbJJWPJ3JCKrc6vS5tYga
gjhrBt720Gbsd84+f3ma4Snj3rDUhRKFvObP4A5CLqJUrYNbWvUVVM8uQ4l+csok3VlXIb2VY5j9
ENtlJO2yHPpg2UIGKg4q/HOsMwLwz7wQHB74gnVkqI9yJ+52PogZPBVbf2QFcU2igEYmiiEjSrAu
h1woMJ/xKGivggtNQxuy4M/DBaYnUkG/s7haYq9WMfWEJeCYadL6teZVIq/+C2hgzl0cYANycAFr
KhExSYOF2MCpAsV5cQKdM5EXenjcOavhepFDg/Yo4YuqD2AcsZVL6pFuj2fKKLng3BAcgd34c9m8
YvnK00foHE+U0cg7hKOB0vD24lcGPgSO9il9NTtL+w5uvpZdLbJVU+otPRUQHTDJyvCp/1MDE71G
RauZpLuDdfvml1o+zxOwTH4OezTfrj6xi8UFaUyiNDbFYeim03rDEVGjq3BAlP5TZ2DvbpX65wWM
oCE6HpLtvZYHH/cjv+NzUawSAxYImLEY1+j0D2NqrXBqjemaDWLD7bEfUgne4noyCAMm9JNBVx5H
+y6hKTmntHVJ0Z1Cu2Ltj+PqiLLN5OOsyKLuPyztFJvh3vST7SfRcqS4jz9F9fhQ1krr6ot6UWRn
S0aAqmcDYKgry8UzpInxujvwwOYouTah3wZVWkghNuO4DbQXhrFxQvkATyIqvtXvV2LiVfAM3jGA
wgApcI9IH44a631ekQTBL3DZnEOKzTSaLzccJYeqxo2NaYKe6vBES/ikCYRbEU+ijytxPO5xcZ3l
P+F+fdMDQiQYwqzg7GxoddMXt9UlKgbfFfYRelhgCXqFQmB6HEBt9ypZexDerVJisq/zj2ySk7q+
J5UwkZLmLjsg+bqq0z58kJMsHBmsvdL1t3wCYsZVa6mPWWgaVUMwlr7JN54IA4EFLp5BQjcNRmw9
lh81ObuNIGn2obBZpsX3xf1Hyk0Fx4YY5lmZ8vnnZrXHwtRPuNa/1InXcYi9GnvBguwAtNTTW/8P
JGI2SYtYnrsK74KJMRPIBmB6w6DowxCGNAH3ewRHlPGVA6mDRNCe7LCsKRaA1CAdagEblqPZqBwd
0+gbPQZTkWcnKEdLWpOPpI67hb6uVuwmHqTgAoMYqrRQtNy9ufDp89C2yTeXLs5ayvhms+Ws1k+w
wQSZztWH2jslErn3v8w9n4F2RCIdMzj9Fz5wiJnjIRTVhamrCs6g4DsgJk+DxLWBzGMo9K88xb2C
hEivjUXvaUJB9sOff2BrB42ZcTWDVx8lHEoG8EU9GxvEPJsGKXWCtSSaX0udZvzKI9GYesEG+YmF
L+ZMnmsyb5PoLRXZWo41RqS4w7Oqw7QjvV+R3MjCgSxLM2zyh0bMidRJVSYE4CM78ZpQQWRxCRE2
F/k8s+5Q0UR21IRUBSN8fNT7jfHxlFn4Kj3EyhYM0ibgxWb0Zt2dQ5dQOH8gYxqNeWoElDcT9B0O
XVSV2mM7Befl0Zkfw3l9Mf3Q6jqJlT+f+19bwL+SUBVqutvhBio1rRuHdRmH28B3K4pkCv8JNFvc
S/8j3nDSsB7TtV0jEKKujcXDCGxlhhO4QfQip9L4sjpTNOzfdR57sdsfi0xV/uu/r+O/YI2l0lri
JX+789llzCGtjCEguylMMThLocp79FiWN1lrjiwiESXkXG3+weujQNPRrmr1UT7AnMADfX6Ke9B2
bgQ1HRmock6LCwcmwJsEj7pnIZoSTXarAqOzqHTBi2WQEuN6vCB3bATO/mYkqcss9HZVslcEPczB
LzPacB0SA8IPteiXqRnjNRKWZeapkWKYyUTj8PTTGOfMkOHxyXcOEZd0vkNzsCssekZ1Hp7O/VW5
Q3Qy3XlB2t5JQIKYZOVfDKLSB4u0m639SMFd1AZ8dZjCC5cMakjdNiGBFF3Mbdgm6IEXHk7lCw2p
YsUWBS2X0Zb81LM1PUGECTASxMq+e5xF+YTrCPGKkw3TRXwZKG6AnX4jhDDUZfHEq5xUYDXxZ6a0
gO4/TWGQVWCQ/A3LMdf7dqzUjIzWZlvZ45LPCHDjHOGmVf5IdzyQoaK864VXrDIi4L16XD02v5uy
3YvaEGQSXJtdeUkikWzikAaXLgIlY9ceDZOkLGnNcPIcQ3I3/+K4Xr6gXNxIJVKBQf1KN4DZV4xV
6PIYeCUf1mREsI+iP1tQYq+BVKniqyBLSJmgCcuW/lYwubpBC5EGRRx1r9hqPU89DIypxk2fUvm7
qjrBqm9tEREjICudULZ1QOBM2V2HKkHlZ/J6VYviiLGbo6hW7Ezt2oJ1DtEtvRuPPVPpZp9RTwI0
sU01IK7yNvOjp+NTWt7UFW9Phrz+KeefmnBvQD2FjuUC1pvICpOtETLpz7CsMqxtx36Pm6GnCgj7
OYY4/SiFoIvVBQr40AZK8EY3jycX43BytDjOxh8xpg33M5Q401R8xkuKrRl7toU2lYvGRY2AsxXr
8QS5FuM2a2A9hOGOz6+0/rcWBjZv/2weTYIqGA28ELzAZa8UpPsTsMiSFLEpyUonSDiFxQyIpqQu
uk1k9NpdsHym1Ag4hiw4kwyOb+ICO+AXmOD68AgwA/2Bv9pha3isLh1Rsn/WH+numln4C0d3NwSW
yZrHGZUFKs6ADrFWfXkduyza48N7+KL5Tj4ifVMNVO01h9LAhDxzCO7Rvp4A8P48I6zmt1xembTJ
g5rydgPsJnjeXohce9aJeeVVjz+QBcCSZenjkUPRoKRfvLE+kEdJIo31F3gaHQ45wg86qWb2FMmL
YhRMaoayV4Fb/dlu9mxgxui7485hQ2rwAPUtlFXcN1w/nHntVsdxJcjtE4j3dzESdIGjB0X37RJk
3CxU+du3BWT9YmY7Hba0KJ/lcMGTukMt56FfY1eG7FLBs0xLfbpB4opVuheQ+Cq/N7ux3tUvCtkQ
ZgRzQVHwrDBKHD81GacEK8rIv5y+vH4fF3/QCndp3yI3dClkaJaYGH1TZUAkho8iVJiHXh0F5/1c
/YUh4Lw7UL4cg+TnJkdmOZyWpwPKrfkVHHLuoQtBTjcNnxRM42mMcp3aW9mSUI0ObKFe2JE10zIU
22qTO7HQoPtX0J6s06rktxg4spw6p4xJHhFPcmm9nx6tPAWR8X779yjP8nLZ4/eMa+u8vMfDxmha
24VgFbFZDLN75JmQIzpHV52g9mGtgb5SHicas899GWCUOxb1IJHeQsEId3rUtXksi3QWzml5rJ6e
RyPD+o1UyoCvMpfJq8BVJo91FxkOOB17L9bUroVCq+qk9VXmChqL9aY5FoWNDB1+kZuzljh0jmH4
NA4PzDjiTzAr83e5NfOfjfiDU6vGhllFLTHEuYQLK7N/N3PpqIAad+eQi/17b1KMeR9SH1vowIcv
w9Q7eViyphU3LFS9bXOyU2iXYzCtucEuQ8cosbP77lLnOWQwAVxO5+rYcvcqAML0VZgX+g4t9pTq
xlP3ti04lMYX75Vcc3l+bxdGduR1ITgX5a+NhPTVBnGy3aqb/iSRfH8Ez5Cr3SGX4kqkl19EUyPP
ZeGb/qHG+8ZENljzuWSyFYHeCOz65Worypw/g/zha6HFItV1PUH91Di0Z2T24ul871Jpx+s9hpn1
IVqXrDcma42iNpg7Kei7bIkea2VI8wwt9ANkB2bLiVWwc0g09GjYrd6NFpl40tRTd1nPuaJ0yqFB
Sllfoel4z70VhYDwcjWmpm2KeZlCcDPhA9CpTn9n/XYoCS4/VxpBZFua7j4d6Q80EmnePF1gI1em
uOBvc5GRj4WauDboriPQNQ+c04+dIhaG75H9JRirX5o/Mr/GzaKuOjpOqj+jJEmgboq5668JxCQU
gInBtJyfh5fFvhuoD4ks+s+a1N+WhpdyHQMzsTzMxZSZVXtJ7V0EueQ6yE8ihhNJQGmKAHvMNjlr
yYniEWwDUDOsqk4lVJUsHTAcVCkPcAQO4yiroj6JHeZH+EApyz+1tJEPpWL2szvYSrHkvSIcWVJ1
pVHSSRxKcOZgP+rKUPXzbNY/0T9Tp7m4dcrCy9McOIiDB/zDgRZs/3ZDpHqSbITBZbkE5JezERR9
xcftAndQ3ugFF5+jwrs0/0rvfMrrPjwuhms+JfdsmzZ6wIpotzzindBqDdbSpUs0awG4oH0doXZl
q+z1ukzSqwBC36pOMyUFjMQ1SAWCopSAcjHP28+VFfNsy1NVKnhQrtAC5sXB11jWxzZbF7XOLlJ4
p4GlxmddnIRkxp9JXOcopKt0SmxcDA+DMlUwMMghUzFoV+PehS6HzAWz36thgE+cuNtoc+hRDstX
EesbhTgeKKWSjdOh2SDMWTlUzSj7PBMr5Pbg18BWYNog7KkZ5Py9WL5jc1mnHu19mFGS0q3ykqq7
BcqQfpKsAlUtl2Q8ihc5PGIw2nxW0rwH4QgqDDAo1isxui9kM0Z3IR2KSSVkqRK+eTHxF+S7WsI7
fDDcwkr7TIDYt8WE6imcOo2pwjUGCglYnlYiBLmu7cwWryBgIogrSXJnJITK/xKBo6ichtVQF8sa
h2/QH0edcDw5kBZMwrlBxLr4wdZA9250Qhgv0EuA0qOWg6UfECHBzIUz/Z1aWisTFc5n0R7864nD
E2ZuVCPCxUfiQUzp6gHvG2Qt7iBFkL7FVGttxLNvu12mEEVPlzE/jYZlZK0eXsXnNqlax9d9Gr6a
v7lsB8HO5l/1dDrQTX60p9zMc9ZLo26LijZ0k2A1Aw1hRKgDpht/bLa8Qkl/1ULdoAo3BLet+M6x
FLV4NmpmZEsA9bv90cJEWeeHJc4nAJmlgtZs6NcaxXQdLz7ARWfTTeGmLrxpBPQKLNuBMrpRjNIj
pdgMrH2aWeb8Z2fo/ZLAbkREHvYvl2AdlyrZK4L6BgyoqERB05GeXe+Kh1g2SoKkdeWsxDBTex/+
tplJywaKCo0sgLd7ZWb998h5A20NnqVAH2d+sh2hkpooNYNkip9mXcsu+usOMuv1AVy/0BmEX31G
Y/JU9WsySBQ1tYCfF4Tlx4Vp5aIBafB+lNNADJ58NoAd2iuY+k9Q/oQTCieD54qtRBY1bZg/L0bI
fPrWFzWl/V88Gh/6gdSa1HQ9INbU+n83TXqFu3jZjxv2Z4pCi5oEBBUXCcTmWPOTLFHcekCKXNq3
dnERXewPHX7aZRUnfOycmvVBWQsi+C6UOtidNcTW+mPoWtOer1qSHgPd1i89KkAXtIElp6Y19vUi
R8dbcwravuqcD2nIkF0SKcIWanzg9HS58OzjVtgO/DjfFyYgYIcoUtAyPRFsU/Od42hh+pkne9iY
nqMemyzs+N7XDerhhyB0ALnDxE8HBQN0NzyKLn9X74LQqOjOPOvqvhQ+sYdYYwqpKWBbtT9nuphu
Z6VaNmnhCibmBrhSa98tRDA5rRjiqMHY8Q0vT41s5kAfoRoSdP6w/c+ppRdo+Rj8QaO/bjds9Vc+
IVAytPulKMWq4XKGNE9ZZcfckC134QqzY+Z6z7FuZjCE81N/LgCBOr2hKF9p6PVUabSZPtG03Af9
O1RgAZP1iOa3DMYkyxmD+nhydQsTi0zcbuKRqqsRxxHg+BkWf3AF71whk9JQ3GyHNct0ZS76kHVn
Kh0WEK7JG4khKMxEvjcZuW+aLNhWUncXYfMsRDIHiFQe4Sz2ZbprBYLwxnl+32Rb1FBbTDjsVWcT
Wa2YCTno7pAd/qtjM/E4We8bAB10LqIcWs6gzKE7m3gmjIKOAlznsbbB2/oZzCR8k8jzvhzuYRGg
5TlbDLsZYPkCUrc6wlZXS1G9koi5o5a3nEnE1vRq6XOvr1mmzSJY1B3poFVr+R/1LQyHAPmgdjvt
YkI3SWr2OFeEjT/KNf/ve9b5gnxNW1jhI2dnrxsMOy9AZWiry0JNxX1Hf5jfrvFdNOR4y9JvOI6L
NwSh8VBsVu8w9/PgM9bcR9YI1iszAxab5CGN5KQYpaWkLmQDPrvzZN+nT6f6b8Z5NmLaGsk+hpaD
ycL0AhTx8hves5WdQGdH2vJ2ePqWOJ9UrJrpHcaYOF32/KVkPqICiUePNsYYYLkEWjpYHVwCT6BP
dbJ5a7x2y1YFbLicWO5zxIOaHvmbadsV7P8itveU7dyt8UnnSFPGau8KmRWunnLWjkWCtz9BN6kv
tY7dvEu3fsXxn/DIJADtSF4Lr7m99/o7FmUS86PQJpxryks+5jmBT937ilV0qBa3HvSy6U7Naw1R
CRP6/42qAZ35mmpKfuzC+ANHCui57yLaiZdzqRhlQ0Xx5ZuY4pTs+GfxjpQTBjZYsj6nDbNQUSre
KCjBPW+qFnBHxt57f3DUfsBFZSHFGatWO8cdYRJ4hGW9LokafTujYDimQyHilrIsXRN7tnioBkd1
Ogeu+nVCDIKlr0F8E3dCMmRkqLOwbQ3jenD5f9GDZJL7H+RtOwVO41/s6eZ7KcKVqAAIFzNpSV4Z
It55QTZRdUunKObkn7Q/bgMPL5z7aqN9/OrgITiGXUiq+Zhs+mL8O8UD71240ViJsngHqDqu1Tuz
RUE0Ew2S61jCaXtNOB1b7lG55hVZ5VAmXN4wtMgGtCZx64mR2tRDylM7F12YhSFetsEGAmrYPS9f
TnC+AELDJcHbagGu+5xSLyfZYacxzXMSYejsUByLYgyGy8Kq7nnlsh0af+QQxdkL2jWXpnFFLfBV
qw2qNgryJIyk9PGaDkvQ5kwEuxqAgoZsmd6m4JPcJpUf/GI9wlz0szQJa7nPf6dsG1pndhLrp+xy
pVAUzH/D+t3GpBqgsT8jNNqOBF+62rgcHqDaMf7vAtB4U7s4UznnT6Zl0uzwU4Qc/pOrHQDzQjW/
agS7Bb2Y1hyOlxFNYF7vRDAmjpziRh371HYtc8e1kLadXB5lSItnwgZ5xWydn41J1v7wl7FYrLv2
YvXs88hIETHgOhLWXjTYmEIWh003l6OpIukmSm4NQ3y4GoOXNL2xQkK5SyMfUAyk2nQPqEraY4y2
Cf3KLYi8fAq88KqXZig/17GjfHjD92znhviGF/YCUMYQkLZ8VAjbzd1zkUM97of4FiCnBki/v9zg
BQMvxfz+MQtE+nbSMFzkInlGy/A67B0/Jya4FjO+BtGkwj0QVnUAACubGoX0dpZNm4JxaPl0t1YG
CiQiIJgBWYGHk9zt3xsbwogdOYcvI7E0e2tM+YMqFAR55Q3od4m9MMBlaFW5L18Dv0JkorugRsCa
AJgfyY/+I+upV9qPEGr9/2WuE/Wdl+tdp1czNAkucPAoEjrk1+cIndOVPoenN0NlSUlyn+LHBJns
SCbLQSvagk4pUYfW+yOmBEGUyoXvAz4oI4JxHLegoorgGdj0lPx/L5p1hWRsOml6GldHoyJeiHZ+
EsC5w0j1TnjVseu7DglnjWydvHLima7/G1AUQIeVwkwfco41tT5So1wNZmVjTcvWVp3NiDMjRhGE
lXBRqG1ybn/qjbtSGH8Lio54G7oHJl2t5bxuiijBb0ZUX9ZVsfPrIV5S8j5BDMwl5LZaacx4pm2I
quwFlSsOuubtC0lPp6Bvx4HVSaeLY8ex98X3ymr1xNHwtT92KqBbIm+wbmCPGXK7shsrwsyipnLn
X8ILo4jSYz9a8RjI9/cQ/cQQf8nv9omu2BEtwk3Kln0QUeFiRqNYMziiCQLjy5r8qgXR5lwarcX7
WsdkR4cnJG97SIAGElDH0fN9iClbZWyUAPoiIs36a5wjxCNx118NmoIwi9SUpES8MHFMYEtQpHzM
9qxaIzzr1T4HKWTIZNvK4lIj7hyIQ+naWdxB2Hs/jKkMzKkY2owbtmP8mXIOzq9w066oIRuODOH6
i02+7AekyRIDiRkY5lkrH0iRVh6KdcE+mHjSt3MRmkNBLyimtrDCvgXPMBe6epKoffihvVrfWg8X
UWGfmvNOfuCd+bGvggwRvBx/94SFMKDH0eJPCGqBHXdneYD/H9c0ajv2C/Ug0+ycbDRTIrDOHe/E
iQ1WxTP3wqIZRltLz3u6ZNoTKCz/uDJbXcabE6nCi++7MTWx//ZaOe1pqmrgK56FJGMqwouOcSDV
jUbO25sz5ZDAz31v8rdnhIEdg2HvtNKTnTWACvojM4aqn+wwFarzQXdCnEJtukNBa1J2MNKlNADl
kMfTZepXERzechvAHAVI1iyGS10SUovhrm5UJRxIF0jg313gq+GEle/04n9SH3eBdPRrPq7aTenG
iMwxMFxtAkctiUzCRhEr1NDENI1KBPXRch7PQOlKaJU5NZwXJXo+8zgxtm0Q6wQPWbaEj+B2wSTv
8OStST7s4HwDllEWofN4M7X7nAjeZMu+4Tio2bXZrXE8SaTTNsLzgn+ZbUKeuXG0Bj6beqqUyhL9
72ceYleaxy8B86sQp5AcoEyc5tNeWp721Q29HJ8o3MpwTBVuoqjdRbSPNYtL/VcArDRF33j642rR
ww5HPIGHT7DEUvhbg5eIkj2zW9l09q2cmsH3572pgqdh465qSwpREj4WapQAZcc6hYYSrte1EuAa
kjg3gQgxTmVB86vB8COT/6wyrlMYyDplHMlE2oGzbPFVv51ikUssUJMZrgI/Z1r0zHB+CpidhUwy
n3z6Te9arQlRlFJVsQkXYUENukVh7S7N5l9KbD2xKHHA6W+1fLa2kp7xW8JYCu76gqisFQjNAjE0
cfcWuFPfk9XOALcp0yJRk+Logx5uldW1QmQxVXbluh5p6Z1n2DNM4mQvDnGldzynOX/td97XR/dM
xb+LF9lt7EYJ0PaxTlmoFaG04xx1AOUx9G7R6e7koopzMdIlVS9/xNHxotlEAIImRQm0npZQGSFv
6UrMErlvqC/c1d5gqkM0UEAjfyHgAOUnWpThJupHPhchxMwsHJCGRajEo5lX03+QJelKlzY0ebXK
MWlgduONxv/rdcvPiLshD7/5DMft9neaDMXn7JaVHIjUg7kBEyuH/mTCRJWk5ic6uCcCFCihef1a
AtFxUoJlRI07sBzg5LzJuXwepsdw2DSqbQJTT4M4cqzUC7Mot++jP/bpT5ujd4nJBn4StwB1Xe6c
VthZiAu8R2Gy92ea9fhNUFF/GDWimT5U9zuiQmTQEhB4UdkwdhGZRtCbUix+yRiRLnNzTXLsI4NI
mifJVnNwnM/H3yKVCFdZgFlftaGd5p+ZRodUPLoMCXZcH2x+gIZPle3x9qImtSvDOtoVuNMKmsw6
ytuoBe/XPiNr/WjH5DzuFvtOvp4X8ge8hxSCzvFfbdIxE5ubkNoiUDo5d6tFU5bNpWtaJnocgjMa
9KZi8dYp4rCr7qBOhkzxOSkHSr4iXkrEHTN2Ti0pkAdwkWoUESI0Xn5vxdtYmgA6tXnPZNIn1ppj
5N/kc6UZ6adHz3pPxdrm+xOOSRlUb6nHzHl33v4zBVJsSOzuKYoquEI1/0wseE0AcqnxBbcInbIN
wVQTbq6IRXFw7F790RQO+hhQ2bQwiNPxc5kZ3cal4tYC6ciElZGPcoP9Yl8W9tB6AiA2QCvoHt8g
z+wb5Qb3cI9BT3zoEtX4goybqGHeDwMpUKPgfkoaFIRwamanW7Yy+U+wWIfbMuMRWU9ehpieOWoj
ax/XungIWL5aTomudn1ylI74gnPD6sL3e5V7Lhj/y3Hr0dyjD6ElMqcpGZx8SLTNSaNe1WxYyVqA
0Q79RNhtm3X7Bc2l9Z6/HljXrw3JiNeTkaXaekIovOr2DjH6LS4kphbK/q+5+K74hGtr7ujApdCd
JPLhPoyhB2QwO9AZzmg0E5J6Tw//mzEP9GZsF1jTlvlR870RmcQMliWFnxwutcdm5YX/G9qtkIb8
g+AkgqlqO4dvne5guorhohBrk0wC8D2SK/SsiSBsyfq4u8PpemtjmY3tC5tqjjMH49GG4ItetrSM
XVCLiKaz6LxQKvUMPJ3JhKlpOwFpGPOJuVDYZwz9qzK5nskv8RXTH32jdX/jA0sdcl6QRHrUcpe2
35WiqpfOb8LkD8yfrZDOdBw+9kYBPu3ZZ8NXGqC36h+0sNavyRW1S2zqKs/LbEB6GUB8v1cxnMl0
h1hkmtxWYRaJ3oLNfwBylqFh2liiBFjPGTWWOsCJoBvuuG52CseLKyQS3Tn5iH3+QuAuIn4q8V6a
paVdRh54EDyO9gFINuP/CsOdmCw1OLmwAdStkejvplp+KYV9C7OFRzESUUQ4a8CluhF/CgUn6Hk7
blcVtioeFK7WQSztfJn8tYDHJRJ+Wtcy/4ndBKHxNVmy6HltUjCWiqgxeD+pyqGoCLhmUbiZ8W1n
LlcARq+dzr1/3szlDTMxbWo5II5dA2yfZ8UJyLWiDH0ZX/lY+PTfDS5EABhWIr7BXt1HIGJAnTbx
KsLzarqK5jmOm8tzp37MLA2Z3F7T66w5ZCBn0HmDzqww2B21pFVG3ncEN1E6zFB21lHUJh+MJqgL
6v73AlBjLUZRFEEyinNJwq1XqmdtU/Cl5NGvuSMMuPxWZaNWXuojqtDTxGixJObAq+RNfjXLzdPn
RT4quegsl7f0ClBRmY40g9N1Eqwrun/vBoO0y6o83WTRI7zvA8Fl+0Pn/eltQlC8WdRNMUd0HYZC
P9YTlEl0dzb4QxXA6Y0GZTjnEyAFa3ps5DoM/edOhdeONaJUkXLcK86Q3bzOEfUPmJs9XYcoc7da
k78GRSkm0bvYlLlpqg6BP1b+ue38/t4276LIqZnOsvhD2lI871/GqAUo4FFWyyBY95O5Vw693/7Z
UlWC/ORuU4DO24UI+ABeGbY5CHHdjJHn0xLV+96q8wasZWrp7uaZptOpuCbJReWbj7kHNOXIuBnI
C1DC2wuj8f+/4xqdvfC3qJI6QXZmtxzhdHoBLX3i4NCBrwuB4RBWzlf2fLDXQC03SuQMZuggxpTQ
tpyy4Ujc6CXJSk6ITUIRmz6IKDBslWVbd5dDJScdVkCvJpFsrG6/mZFs44o6lzufqDwRmalTbiD/
fSXaEWEARhs7dAUpxjrkcFcwzTTgy5510ZxtYkywVXDBX+mwQqaxUChpKQFddJFwgM0ggn9Y7us6
3PEC4ZjtTO72wcvNvEUXwDdevEIROHx7svdOnPiN60qG7asU1qa1K0pmCAvWzcFPsncPM+x2YRAK
SddzO+Lwc7Q9gFOik5kXBKAsBLjGExi4GS5NHzxvlcWj/PvQlrCOam9lq+xezDtB7srRd4AJ+Gxw
0P+JJGKlcwQj3XT0B6XcAn+6vlOeqebJHbrY36GzqPcCPmRvI6b5+OW38dxX3nTPu/CoBqdCUhMN
sz6amzHAJccAuiIyfnhY2Kp5NGvFLh3q36OZTh4jxhKB7s0GlFpkLMeLgsrN87Dp9AvbgezGkXXK
p3+BjLqbhG+KIMWUdNrLgMpxXR4GEeiNOPMH2qupFSQZwViWKFkPTlxRvV4ixYT88A2F7HhFuoUw
5W3o6RhMBPv9CNmJZqaoyu96lKZFhGjzN3hNMengwYbrfEMox48rkySqiJcxA0TQ7HTSNzXDpfDN
89hSKW3fXNbcnS5C2tK6Y0tLthysiKexoVJ9PnDW6Rqt9jL3aQIilN5DWJgFm1+spkcW3Br1kLiM
aingAqK+SvV9XCNWsp2b6gxZy7c3aYEIyPLoVJCXf1nensAqIwO3cUSe3/5/msmCwPbrkXpQiXJz
jWrR2zw9s2xxWcMbmsOHTErKeiUGtOdYga3v2FTDdl8jYqSnmuYPOsqjKN8Y4yIaPCb4TFIkpYyb
tbA2jZR0a1rE/MjBz+Hqu7b2WcIIXWOqTsSKLrFyDLEo3NvDBUuav8toXntVR1suRWbYAlu/LZP1
ECeN8NGbM6HKqcaSySvWcPjIUyZgNdQni0cj9ZfQMrLrCGxPttFXAotHu5zA3m9rRRLf1+qhYJnD
xjEas6HdGwzmmcxc8R2FfPliRiTyGRQIPGm7iIIusO/dSSG4c63TePPQiDleabLPUaZYuGlqXkvI
5W/ZI30DU3XGqMkb6NRSuPfkDEfuJqT2escWwEbaG6140BX3jMeKUSEMByhia4NfBpH8AOwESDrt
ogpk9LRlfmUQmZLJBdvLrROLFbYVnZEOjw00nw+PxkMDKXGai1JjmIgiU70IEU6c+MiTS1JU5wWh
m3MZZXqKB5ddhQWq+K591ClAbf7y6uCRV3aMZzDZq9JkoPFjdbxSWi0Z4n7aYV6PQ0ka0vCr9Qk+
w8NwvOkJEtRnq9S9GPxUT84mKii6v4bL9R28k9eRmb0J/BznENjyGop+Hq45eJ/4+otsG3b972+B
EryOSKBTS5YFMYL7DriN7RUfBa5kkYwG3lIEVZ8Sy8ES27HOayFpI9rqJixnyNT8VTXOQVHa8GL3
9S1cAHrUcR4/z8vnStNLUxQ2eBajv4M996BhttM0rsBUluAGVxRJUSGG1/unHgQrJ3sg4XaWnqp6
v/IvmFMk2bIYv65NSh381RbTwlarr2Yv9dP8JhE/A0chTuNFi+xuTLut/1+TCsXp33PX6ZbmUYA6
zslPXmtQsuwmM+zsClNP3hzb1Ca1qrAheZolFVcrULS4T476ptIrhoEuC9bpt1e4tRpqthcMQ82j
HZmYpX8uaGYWViNiTcy5ZgE1XQvjb2V/RnRR4ue9cz0U529iN/1IH4pc2gjnLJmyO+P3GqmA2krc
aoKl23xIrInVERaSs8CU7fwwJLUi/I2qbM5wvasOy4dF1wrfhShLOcX5k1cvNQpS57TyRLnwv2Mu
99EN8syXYryMMy+971rLY2qlyBMt+zpseCba8Dik6ocCzW7lqYc0pSNgAUzc8rlww7ydNF1Eu8L8
WM6egtyxm9B3NG6lTqLYacsk9zBjkeR7Na97De7Pr2gsdmxmhnRAHv6EgsyQYe615wWgy6+cFsXJ
fVfJSs1i2dOFPUHm9N3Hy2x3J8Ydqvkiz9veKzZ6jVGOZ8/IAhsuUzjHRSu9EViLDe88cO3cfX6h
ack0v96+VwQA5tH8+r1S4I0N6+PkuxEbGCxIOO5jcUuKsna69lEjUSGgLpt1MUCrv2Sm6P7WS0Ka
ikyjpgSW6USYj/5kWn0acTFlzu6u3VQZTTgFJB4KMAGCoz85Ltz0PX8eYkiy8AnPmbCGD8RfqHjW
zmqerkiET17i1pmX+L5RVQVORJCya227rIfsvfV1Oe3jHwu/5gXqyTiQYGeE336gus6afkvL00fQ
4uwchhMZ8jDqZu9sHYZMQ3ssPorarm7k6D/IR46peiSrrX5Rcx+Rtn5uiWqN+143zxm2KImYG5Cv
ynXVP7p0NUAktC8/s2xn33zpE+ujUzYV4doZXjvvDwELMnRWkJ3NL4oeCFJdkvedrJn2jp8Etwky
6RUuMV57cqc2NNSX9F7BqWygvFgE+MtE+Gngp10VVHgBy0Zy7gxB4bU89eGvziKH8vla2u5mpi6E
yfb8HzLJ7GajIr/rtaeiiAHmFmXdoTVdIUjsKP6mVWBZynbAYnDLfvCbcpuBbEFSchSuKBj02wfr
1Gv7l6Ez+MAAycvH/roZ/Suqw6e10urjrMrq8syLN+FXBseEm4wSfnwyY0r1wmkD02RAj4Vsb7Vr
4PHa5sMwi0xM0t+66zbGrYyj+t68C1uRs46GR3jbNLO+XcVo7Rf08cVmeYPQB1Jm+c/EVBdnRsYj
MJoBq05FF44e5NIdaEMIeW+rCZxemJahIOLEkorbucNNDe/ZHQLcHK+rINZBFQN1KUEvEvuUCpe5
Foh2x2LfdQ7FNw/9+YSfvyV54nfPkMeYaymFuQ/6yD9QG9OCiNWegC00qa1uZDqg3pNeciOUzSoc
q+aok+G/4dvl7VVvrxObiyp520Kz7ifb01B7oEWLaSXwwzZMFmj4kLKS6gU5cIPmb35MdKX9N6D2
M8dEFoDtEIWWdBwluGIl6fufK/6WitHkDcQeQDX9FB/VuoVGORfJnsud/X07lfoRSsoz9hSulqbR
LN+AdpMln0jvJXoBnYfw23nGrP4a6Wpw88RMWClOR+IUzEQ55Fa85aUZDc1i7cY1xx1lF5oc4rNW
5kM6kEEwFJ4B69g3ApWWN+DscQ77bPtFyVFWiKlkLaVCsOd94mkGJgfCu7jgcAJ+Few2y6Ps9zSd
E0H86oMmDzz1D8luctY73xZXC9GwQC5Ga5qY1neB9SwZpCUu5QhMrYZ5oAEAgkly1Q4EL5dBukks
T5jRGXg8jqqFo2pFCKfgmloYpkAKJpb7PELSKLtN7C5tnq9pM7o6AZ8nQ9qYnIJ2+se07hMmJrmZ
6l/yD/qn/UPTSJC9uUs23zs47o/ObAHBYZCFSDKEsgPrTc2TWGRK+qZ7MpWZoitf5naDj1z5lOfS
umu/jDpXs9aeiNasU2QNiHrwPsCh+vBMhLbXm6BVFtoGh9QPx5JmZ/B1nII9tydvD4E/GevB1vvz
pvVK9fHlCZZl9p+JJXD3VpLuu4DUhVAX+u+gYOXx6TKZvDgitsBDkCwzge+MgvWuk5xYHNf2OsjY
6AAzcONue7nzoZihU6Lk25Lk1Y8aZC3LIL4nSFIgqP/bZfrX4ti6kegAE5VjYRU06QOL7nytniR4
+zXRn1OieVNzvvEJNrWZH7GZUu9YcgqqJojz2X7/Naq8AXbApSJsck5KmQimN6Xyk5qm3Rl0ffD/
8qeU/YPRJZ4wruOHCnpTLYqk1wMSjkAgWaLv0ibIAfZM35Gh5HDkWFOxjnNanFwvt5b7jFAf4lzV
DEJWLI5HmrVwrGHflxn+RypIm8w1ne88g4HtQc3ZW80Z7y6YYlM6ztWeL7j+4X6TDB318o5tJnYo
bHJA83bQ+m/kyZwPzZeTvooWbuSO6GrK+iBrfc2O4Hi23l9HRE8mM34iqdoVDassMOhlFDLwj1pe
/lPuRNjGJ/ewZPc5ckspyleF88sDE8Ejg5+nyR/9BmeAycmBFl/nIv0jcV+t5LGti6XHHt8x5x1V
gAQ6mI/X9aL8Kzw19KEyMuQFjZJbpqn9BwTEULQUQrGDSj+xmrnCVWcdZr/uedPPqjsfi46tVqEu
OCaPtnFssLCJ+YHJeRDX19kaKdkSyLJlvCnWE6bPFuTH6bFcRa1XfYRDuopQl5zfFHj4K7jyLX0X
/qu1uSJG7Hef7W66spDheh6F9brDEJsXmBmKkTBB/XhmhZw95udO5E2yV7HNQYlr2V/Lj00ssexk
fUAxGyQ91x7KNot9/4JBVz7f2nP4wKimp/5tePLCR8LrneHjMzm9eOWpj9gPe4tUc7gfuWtTz6Gm
BXg47NlXmC2/Zv9T/Qz2n7kF2beW6quOlNlIKzM4Qn2r/rhM1lw6n2deYSG+6O+gt+muE2Owxswn
IeyqKZXvu5iV8EhVmAzP2n/KVFz4q3PXiFI449Dq1b/pY8IHvFojJeTwFwIKReL0LuFvYuv2xId+
Xdg+8WF/iwUh/saIxEq6MxscuPtMvS3klkzrQv8pbcMbK3ZA2OzrH9UsKoaPD5iEWZpZdSUMnF5+
CI8cu5/wFCIvPF/EPEk9Gjd7x4Xt+o4HjB8nJyTecGOH3oOUXpJGM89ov1RfOml0OHiuyGLOPVX6
jSuqPNhVsfrg1Urz2HAuuWlDnJcOwX26+F8Guc8U8xN2ijHjhQf0ql0yEtBacr1G3YFjgDU8O6Wc
8cll17lU6vtHqgmrSZiw5gic7UPgEV47fPj11Kso8NoVDp+i7nO3Ilj5N22P22+gzorLkU2aSrzR
BGMIjNQkplTsMi5nIA1PGReio6jRQeAozuLcUQWVx6HMH/YnFh7tX3/aj0RieGM1Wy0xt+6VYHzy
DN+GqAeR45edyY0yk8vA2CXUQssq1ujEQDuGX+DnHASE3q3DKfTZ4VRYfwrXOSoCrIuMKgCAYMNY
9+q7LA567qm+9fEAqvJHin2JQd6joLA48mKEHe1YHJSWnWDtZC6MAtsCa+5oWwim6Uu4+raXYENB
OllVx63VC3BzdsMM7xGmCCwrjWmn6r57tsoGC8S2RleTd7xToq2BuCIiQBgk94oLTCmEyJL+oF3U
tOixKqUNIsjqCMHVwf5+THafXCAY7EoMyjg9pWR3TQpZVm4f8JV+pzYYVbTeuAHmYRjXFh7Yu6jE
5BqfUn2WoUAj095xZA40tH4wHuJKFjeYgni+4qWXrDpQ675Qo2TM/oDcNi0wz2Bbac1oEVcjwwB8
hMz2Ni5TlO4LuIqt+G/YU2nPN48TjvhN/ksIoXHbPlQv0mpVVn1Q5pnKR/hKWHSmlPkVRV/pjJEp
Z5GjCV/cmfvtxproVQFDVlc6Oa8pmYAkGe0tohh5/e0nzk+gzitCo30LSk709MBLMlpsD9dWoftZ
KJqoKjarIyVwteN8/DeI2qyq4mR+uhi7V2ikmy7KV19msGI7Miwwql5C5bZwwaK5TzAKfT+Yw9/5
OGGFYKPNpxcd1IqUwzo+VKCw0bduymjLrrj96i2W7CqAfcJGMNjoy6xj/3GdBS4YxhjDGiEpcWqT
uTA2yCvOUIVPbbZY7T9FOOoSIca21WXAJfwduVw0QpL+ElxovN4UP50p7fzMzxA8zHiLhkyLi87V
MQGVL7heTD+xtnYeI2OSJr8HfIUREvWk/PCRVtu5ItQx4Nu5f2mevUzhoAD8BNEmWL+dLG+NihUe
jCq0mUpOhRNq/LEBC7lqNx+IjhYabYxRRheKOgLMtex5Btr8qLbP42QBpsttAdV38jjKWpv3Bguf
xA9ueifyr41qjtV1z8INtSK2KA09rE6AlIb3kFQ1UTOpAdOuAmZs1hYmtFYJg+YM31wYN/Y6iWNy
o0zSLYKeW/d6VL5pbw0qT8qXOzgf8iuRq83DsNJLqgAKappD04fl2ZZDsbOjBcgQ/sZxTZq2bq5x
HeR85leQk8Hu8hbvWsyBnCAINhVhV4JKM8/jZQDDgW0BBX/F7O6QW76rSSlPLvye4wP0hxcbYzGZ
tkcGzbAwAaCew4WU55oewdUlmAho3AqyDNmiAdXvPKMKMRexzKWkEy2DHEwwi3MECkBHDuj/yjhp
8PGeSoBv8I3eRCvD4LSr4SroXFl3JPeYuchpFcbGt22BmTrMDyU9h7R5Pi3lncJFqvsjCvf+XuJ2
tEDKhbhqfQeiome0tauthqc8hgvptkwExiKMTKzCbiou4UeogYaBCAQ9iN86i0LaBuI1bOgSHjDe
+WvvKNVHfPySu4AvHHZOgz5pddFJbYtYHEMCU5+Dx9MiT4oQTdMTK2NMIL1gpfdwHRqcEP1CxEvG
3ch3kaF8I4Mx3a3XyiQA4tp3wCHZtgPGJmGJ8pnfh4IVQ256CS0bFjtfaHxx+YoUFex2uGE+e0s7
tMTjzTa8YV3Cpz//Oqk+hNzvQyWZlmnauKkVGmY8+k4pclXU2YrhER4JKWmBjOABK+j7306EXqcP
hwUz/UeiumsukqZAeCNXZELze49lLDURPtU9UYhxG0zaNW3R6zv8y8CXHPsgiQeLmTkRsK63gkVm
YubvfWFmXbA7JwXrdeuRLb31wqJv2d3QEDJee9af9/+bo8oY6tP+tTQ6aB6UpsUd4WhC0+SUnYWg
GAkVU8vhGFPvDSBUXUKtBXy9G8LWjJ+NG6eePDojwtM/4Whgd2nJQ5Xt1Ybr0XJVza3L5CioAjN6
91PTb+EhtqDRkEdIE9ptkeHhKXhs9vXMIZZwmCAuT3ylwEViEULOzLj3jMw15kuLySVt34RKMPbN
H6OrcDuVS2uafomW8k5Mf+VtZ11kK4OGovXXeht4xVsF92LHqr58Wm0HdX5l5TnyXQDSfGoy8N/P
Pq5qT5jFJOFmBqnGAzbEd+77YV+n3Ie18BQ+lNVq46QVbz1E+udJoRA9RhfXB1e7K1TuuHuUFYNr
+vvLlELUQVm25omeKFlDFoYAnq0l9hebnntRt5GRd7YxoerBFUOSCRrFVd71+ZEXBTLokWQdUJyd
O+TlOaE2Ku6eqJX2wFATxlgxDYU89vn3AS6JRBWuW0UMC7wPEggREbtYc3Sw0qlSQPTy6pC+MDvH
d6KI1tVhHpFLjfsf440AO0co3nZ1Wk0lrR9A8DvlWP0Db0il/97EOsSh+NeR+d5fFS9FmIPwAibv
TE/7u8YqM+T5WPlGIBaZgGDfMc8dusTcS7+0qwIbIPHhvQSpoBT7TAhN61CRhtCnUKEKanPvhQi4
2lkbwF7M2Bb2ru/Pp+4VIzCGImHna29X5Iq4+eiv0nA8VjngXy73gMAaaDOZkoC2Hxuf+kcqMiI2
24QjVWX5i6LTLR4jNs+79Fn2i5HfalySmGNDvMRiFLX2mym54zH0f4tRNLRfEoY/pnQ2Jv1vAXOG
x1BPuSqLCmSs0iz5mEHYRhuHY3zrs6AX92ZUoMHJvVxZJQJpMdSN4wFAFSKcBINvzocoHAkGntUQ
prqkSr9VEEXh+nkm39MJwZ7GElt7lim38MOmmy9j3N/FvawPPDZ5Jai69Tzh8wAMRE5l16jbrCEB
C/sG5Whs8B/HTq/oKOLreA1CrV9pVSjLlLP0Hj+XBaBlkTD9wo2a/vdVooJ1khaBundtwzuyvgnP
R2KltHiw0GWEW7EmmWomuWPKZ1/tYvOtk6dh6a9FlzfRWBdAORXxiqvX2YiKjTY8EYWuilp/CCPo
4V6exrQJlTaYPWrY1ehPyv11i07CkgcGRj+m+nNAIX6QUav0nuksU4kPA3O8EDESQFEqip4dFbjz
oZi/K2wzEpdQ4KGyP+fnXo9wLEZ1VAeQaoHAbayA4Q56KuQfI00AKSobAXXb7mCG12DHatLvcVQF
3oLlcuJ9tPJ1aZ7S8kJIPNruMEYQw83Ew1OoU5ZMZv43KvnXID2K3CuRuON5Zt0HgNXDgbCW2wmE
8GdQhe6Oyo7uT7OvSf47ArU1yGnzP80C1EjEhXIZPrYQzt7uVmqyNOB2zE1vlDm5Nl0FUsL9Ehdw
rZqLyXc61UxprBzCP9rvfLwTsJW39Izv7JudY9nhsRqw9hqzt9gDTJIH+FAapePmKER/Kr67rJMg
uu8uxa01/1r49KK600TyAWComYofuMH2FhCeehDmAEh9xd8MffkzcJpMwJMTCaTabVEHPK5ZmF9z
zuqCxVgj5u9S7eT08qU8V5EdgvitlvW4BJ34POLYxZGd5gmddHVFPvD3jHZ9nRly3ik3Ms/NnjdV
4LQc1R8fhxj214SrZ6X3JMs1GQYsX2DoPqNZiv/XpXSJIAXwKdJFSdrDPMVPjCevXcE4LZB9r8fm
yrjMhtR7Sn8HhAIXMhblvonLwZmhcHhDFhTwBTGO4b79cwUrz3D6cZYDiwdwIyI0w8Hi7AhZ0qEN
2IXJWrpR7DIBJ/Rf1uOGZcwvHGkWdzu5DJ9iq7BvQKAXeon5UljFhdc45qMAHLS8xLl8alBhFqrg
Q31qFJN4SNKi0LSHVzFyTfKxOaOV2UZuygiaEEDuWCwu2E4v4my5wP3a3C0ceCHx6ZLe+rLBEoik
0PcaQNpg7nwmG2q8ZJ+j+5Ojx4ahu+NXODMw624qwkLLhbFc6hc15Qw0DI1V/NrYKBAxhcIij/C/
vgTCFh18k5tRWeXvwOLHaXmYqtPHkztWWNw+EHtmWMFi/lvFSseSmfR/jAnE8/5JwaX5eSep/EO+
yxrD5AzBxdSOlGUyOJb5lAlUDuNbKgM0exosN0xv6F4QpV9ALt8JCDJRYNuds/gsywR2+USqaHK+
Ei5FFYo3+wPHq5SOjJwfl6+C86NBBGDGBmYpqIEl3BWxs6gcsblX9bwjTi86JLP2cWroWqOxCc/X
stR9Iv0xzzkOr7U1pWynOxsvpn5iSnjP2Z/XVGjQHL4Xj2oHI2rmsWTgtn76Oi7NY+PlCH8AxOjq
B+ZsGOtcAOhJKTNFGJ2ERllJsbk/QfEWRXSNCeulOu3n50FNnDxbkarPkwR4a68LJixQ8iBaHpWx
/y0XPL9TSMDF4lmcgfo2LFuKf7pkqnRKW4xituG6CEAnyoKCtTtOSHbZ8tK1nevBvM/yS3jTmyjz
8KOsqCgM9YSjyif5XsKELLdhmkAj93YErvXbkSzHHcAJVd7WQ8WGzQGxc8NrszJ167bjDnHxLG5s
G6v9zvXWI+Xnw6jHFRt5QTvoocQ+YAZC6ZJBoOTFtGZy5+NmZeqGx1skNwtvyGLzUf1VEJaQNI3l
TvLmYYZHOLbUl9OwodIZkknDF1Z/vQalvGwruqDHQe3UssDpvAAcXmpb3hPdV0QUY/N4RL6ncC0q
1Z3QM6dRpkrjVbsjXPGLpLPJNDPeFGmmbsU3WHWMz4hUdD3OddQPRt2zDCuFM6++XsM+IfTOy4cn
tFcx+m0n7r+SjPu03Uu0BU2eEcgul3xNq96MAA2S/OVuDOHpna9zyvwole2w4kNc8j1DKFoU7M0c
45TNp3Q0E2kv390Xtfj8pDlwxQoR/QUwvgl3AdTZqKNPEXfIaj1C0S0QARJ3po6XnIItVo08+/CH
XAGVCwp31GLkJPqTzraReCtlrTKplIFrFZSrUhp5NMXsdRIrMSKLR3ZYVo4pFSDwDMr15RYWq8MF
K0pAgEShzLrthFr1fs+DXT+AaBmdwEjY9ujXB7k6K0EM26O9YBb79C5LLl6hYzJdOOpZT5Dpb7wE
q5Ru1tJ3BjD5AhbUhmxreL9jfbGnf9ojpffH+Ahf/bwuRtWlB/+v8X8B51VzO1fqjtDQraAkDRst
Bc4LdNJtBqU43X036ZRbY6CXC7Fd2Tg6md+I3mhjp9NU88oN/4j6t40WEfq67s5fguUZJzomLqB+
5wNBv5L3o2IAogquZtSDWWNVqRmf4LljOD/eNYp7p+uRYh8k3BSt67JiAMztDgcT/oTsztC9QKvp
Mwd2j2qIRhipThWr8792FRdveugVwgVxZpBS57+Epy1c3QXV66w7IlzmxfOLKhGXsuWMu+OzW9sj
QDppKIDBzgyYydFI3p1nXP4J4dA14G2OLt3XvZ+2d4d+Z91B13OcWHY9dzaqcYpSk+Ob4+bcKv3B
07tXR6W0VwExzbRfYHtl1H7JrFO0ZVA8REi+uqsu8J+FDaqcujEzkMsrY4FZZSj7MD1kFBlWk/4s
JArrjiE1ml6kLqh/AR9cQMWT1uVWic8atF2YYwkw6f5U8EZhgJNCJemLBQ7CmJuS2nrbOZ+2yyNt
qHHKLbNApzDXIaYGFvHqnxUKjKEx7+5/u8+nyGf2DKCgtwHYnQGBfbvs4UahLCesbhPfuplOxhZg
Uu9UzrCoUxBzQ6KXdcK7HKf7mi6iPfWFgkTeOZOr/rmjG8EZnCaUBXmiPp6ZGvmiuDdVZqCAuItY
PuXItgs/rM7uXNa1XS7thbhW2WOVheY+eoRGO/DR8tYzhDWyYvE6hbpV28EB9hTDuiucLU6AHiVz
J2ZKDAegBI/A5K+1uTn/ZTCrQxrPi0jwG4+2pceI8YgsqWY1cxrxKduCLYokafNQ23NROp2upmg8
0HteqjpPJivpFh05KGIk8G9u/uOdqpJib2AyqTqjdK0BsUkqocnXtRqoPsi56eTAtczNkEmXd+TR
a5WsKBADNdfeCwKGj4+0rd4RyPNslF5wZQ7535bZdJnvw8EcgMdD/XOhBrhRrJ6n4PhGQgjXkRZ6
tukCHTG9WIb7hobNfnXRUrHxzvJ7YtbiuKLkgJoDNaMv/4hruWPQf2RdE6J25QixByW7v8fKXGn/
tQdJrdEttJQRAHsSVw/y4pO0aTJ+L5E4JezP3HCLDuT0Btsak3Uz3oAzoJMZIn4MMOfGYs2NjW1r
FPEih2bGhJoJTO+q1/96+WNlSPrtD+QmfAdG/H9TzzdGDoBCGDhf4s5p+qIdLAXIkvbF/5PJVixZ
Huw6UZXVevZGRK6+UEFB9lgHa6EYS6wnXQZslWtSjtlxTCCUE7WaKQvZmefFdFqJ0Fpz4DTeuhpF
lL5PRDnRukmz7Jk0nxN8/etujVxDoGktSQgAddMWaKYnTfXSnOEIR1LYjgeMATvNkjpAzZu2LRZX
hamKNMb+T/ZrHzHOXrU4fYHfWZAc1vaJjN9lUib8B9GjSYET5NiIM6orGcdcAvYBk65WySH7sJiN
cW/6vp/qkObm0KO5cyGerQjEjzaqb1hdxvj0kM0fDVXGjN0fiM/tXSiSKfOzphwXoDJhTz26uP8g
F/bRbYCAs3HCv9WaG+UP8e9u5546B6WFi7TG1oICIu9MAQ+awe7pKB3s3f7f+YA+Nw9KBoJhz7a9
A/4kDpvtnmabOHqVq/PhHG/Avo0reSqoJKJlJUQN1RfBXiYjVnHgJegFnPLhygMDh1JEUE/8mq1N
6gWgofTJWQuL7whDCUqgTGactjnYI+AjBa+f16GlymWXtP4Dx+DRbjSiwQ+BAvkgyo3JDQUjuHoj
M69lXpG8m7eebYbCL0NqgYTr5qSrPwY6eWgEqKHnIctK1O8oDzeS7K7g9+6Xq1NzG1wEsHriPvpS
NdVdPmUVIBcVc+pSyyl14rVi/SoGJhS2Th+LcJWaOEO77A5plkBefFGudwBusZ9v6OUW40gWnoOZ
N10T/vLQhA4qCFYewl6JhN8D0eI0zX/MQNNjws6bu9o7OeE/YVRz3qjSFjHRTCf0bufXyOmYa60k
eAJ27fNsOI7n0PrgJ4lw5WziIHkUOufDv4PyrS14mNBI6UYbHfK1P4av5OneGAa+Om4b2fRzecvE
+KyXPfY4raLAVwUEx2TgGzq57x21eFAfo92PaRBgwyzQdh07NCAxnR2FT34QbQ6l4tD+duRDJVTz
9K2h1Wgi+wyBnjmDt4bYqUiERnPcuWD/xLtbzOL7/arehdOoRPOOdYsIy8/o6/3qSiH4aZ9WTUZ8
Z+JGxLDaihz/q5XHQ9DhtXrlQ5F9o8smjXAQI95nQeMUL+q23xyp7t7fKiVQJJVz+WceeRkyfaMt
zEs/V0fX8XPmYJm/TNxxkNRjku+wH+q88LwdqasbYOKtkAOgZ6WUAYcV+7+3bk9K19Qgr95Joy4E
PWRMWSOSmApaIydyaJLrXKieQSJRUTm8wXqEd50p9BIzfR4eivSUHKvbpEpZn8c9y5FDtpHHSeos
APxYyGAoTQUhey3J6nxVZrmn5vasTf4NhBsh6IWOnEBOwiGjsZNaE3yeCKvYMw9Xi5L9PbazUHxU
vOq5X5D3PeF6FP2qUQL1lAABap4QJSvNgEp5CT29raTpZL2KULyr94gzJZMQqUtVk367mtqgBTXc
zD7/8d7VmTkJlRyYYgX8E6f+T4sHa8IR0lEAiThbGhRQ9PJQhEXsCPzOJxOR/OFWYCL/NlPtjYOx
rHYLGpDWSoVzfI0+Hm8xwJkCZmh+gwtQAMyj1vJar1+YO45FwR+4mGk/Uvnf6c4KsbcuyRoMdTkJ
lLPQR/Iy5c+4HQn0DQV3Y2aH6O2ezRRXwRWe+O9vdF9GmiIuixnWhb5QxK7q4xue/taOt2JqCpZ5
VwNDSm5sX/Xv7BcIp4jyzvJgHRGed9t8IvlIqkB9oQSSaRGfO5/RJ263b6HhsJkqbzYBIx4vZ0ww
aF4NzFBN6eZmOXrUrsd6Nql0yCLHE/6nXnZSBOlIaOVk+O7W0feJ3Zyw6r+/7yzOMZsxvXGu05Qo
SZydAI2Gle9A9f4KmEYAWNFNK0WigGOI7RVGXYyLXldFIune1rbEK5DNNUOM4/2U1i/iqkfH2nxY
Ni6Lk3HNJZx2FjibK3jEMQuidqQjr5dODfEZWI9oFzQHrxWwhUAUUlWHf8v0ZzZ+U+s0gevfMP+9
Cv9Sq/YY/jWjK/qR6c1UqUVddjP3rqEff9Rrs4Oy4NwQw7PHQKaSzn1p/qjvpKKL57JsmYjDQNgI
2z281F4oI5iNhRcJhXZV8GLwaJcrn+inh98ZcuIXnmkHlW8tC63Ih28dmrihfclJRGDPq/zFF1/F
bEixychU+nLLOerogKuq17gvUZPWOFnLfgDeeffJA1U2KElcBealpCRxT64Jvs9XlOWU8hiA+0ea
E4+lRHAZRwbwUet7/jG650ill1XgpWvZU/TfQJlej9xfX7dCVmOmW5iPfasc47foBT2GRZwzQ0AG
StVtfaCfKSK2vXyQkV2n+0V4YMqnUWaqV0ApVUU3finvz7DXwbDH+fpLVWkA4WFiP2MWZ8U77lqs
gR8oJB8hf5ThvfJTrPAQLNlmoCKdqRFsbS+vtF6fHX0mq6VW+rMvbhUsrXkaXQexOP+dAgzIrADp
etjskB8nlrpC9XRA/ycKySrUaye3ebuFRjL3PJf+kxsK6N0RPSlTqaRRwcojdWC9N2W5r3athQ9u
PHXFGb09DovjNoS0uiyE1rWhT2VWMfOJ89RK92ZH/kRe400EqxROFOAnJ7t+ErkseTaj0KLi7JrE
tchMRwBmabVd97O5ItbtdasVG6Q23hfA0vvdp+gBxBV0bYytUV1tyAS0tYLcR4E5Id2O5E4BekPk
5kERJeIZqnIDVyVeVmknfEaSrYcbu2aPm+iTOmaNdWPAm3PPytcRWQXe2CRcEHiDwmKCAOL0cE/i
6NCAEti2ZCzshxvzyx7MMyXkTe2I4O2F02hW+Wu+MCMjJ4jR9HrDApON1F+XNeUAdSt7Yp1pkXkY
t625a2JJZNJVRc7pMG4isJ7vi0NI0XHk9l/h/Ih62wYlLTSMOabgbq1rC3ztZNUFYDyZVJG+ZkaW
cQ24+Ez+d7+ZolOz9g6Jy+oPydVopppX4NcotglO/8Knm66NJ/ZVGkrC/8EsuJbAqY+JJCGpo9hT
hDAin+Npz7CeiDzYevtsseQ+lixigDqWdN1Esi8WchOu8vIicPtiHaaUqcBB6Y7T16JPrQiN/sui
2HhABNvwGLyM/s33yUZ4rMv/c0FhsebCXM6fQvND/U4u9twVneq73+6e3wEJrr2m1Fn23begMuRS
AUllWqX8384MouZYMYa6SO1xC3hIFTLuIsK1bXYJN/6r4zHby6DpedV3fac1bb6qakVvK2M+zJ/G
Vi6Lvsb+06W3yZUT8n69Ou6Yry5uOGqT3NUEQMrnYnZwsTi5maefUAEbY8LzMN08KK88M2fkXCqb
x2egtjlwzPkbahlnPTiAjDGdvtzAGdxv+7Phsf/XdMiJ9K+KI4nDPe5QrekCZivt4YEQ1zdYNO5X
PLT3+P0d6HnBcm0zAckfs2PbJHoNCLz+BoE8aBCeyRh6SOuMIc7wPeIgyLJb+vshJjHZ91t7BPA6
5+c1G7VJvIFvXyR3Mr21dOc1Hba+1D/RdO2GJ/uD3mDD/y3enir+/PHjKMo57Jvyvj3yWtf0dQnv
eAORYylua/2HT8+ZiBVrzYh3vOAKZzWn8vjFn58RqwmaTLhLv5zkpJ13ZOSHwWql9YdbVZIPCSWo
/9RXjdN0BumCDbIZMIp5FEruKCtuD7bxK4jm3bVCrAYY7HgfvYVlhibTXogKcjiwSgnS/WNI4+0G
p1bUyI32vtDjtJ3itIHGussunmxwLsZkGZZhmHeMFvia7YJV1re5J0oL2Ce5PKKsIIF9cWOg7O3P
SzQdec399RIhWYclU5yCjYaRubpWx5poNjWEB87W1s9A/pIMiKE+6CLeW0nXnvSnCxz2TDgEWR5H
oAeO8GLxRWAoKcEdpb9i82tMdbZV5yCe/8O7fzgQKLkaXZKs5wv44CXFjQo7I6rMBRMGmZBC/cKn
eIeqMOUbN25gVJYeAMJm9D2mSReEQZtkQXnNhfvcdw49jFkdma4PB5mPD76/bF1o8XWbc0ePMua9
iCvnB7VQsVjxSHGno+z0DXOcDEOU1ALeDenserP/pgtVEXTr5/GJ9h9gtkk7KyPovc+uGE3nc9PZ
wgqZzCFNY3MQBOGz10qpXEEL2sSWeCaCF/Vcxur5YbpmHQRNZbfXxpbkfOxfxQEB1V+FjXMBoY5W
D0+Y7pV8+neLFbqb7FgvUXN+NOysygiJccrDqperVEDNi8s4kBfijUwhzwvYSLOEKXTkAtMuqOs1
LPZUPrKD67ISdjqFu43gtmT2+EfjqgKxXQictCTwEWki2tLtRESGM0PO7sFmrDl6seVUrwnlBOZm
3kfF78xk2g5shaJQ6fP/n+6g1ZLZin3mDLwSme/rUxpARrwNg11e79X+H5tHmBQSd+pOge09VEtk
tPJkGEeLfsZ4Qs56kJQMNbbpoBqThEWoDHF5PxlusalMnK7G3WuvViGbsVgyTQYn1fit6XkqlrEN
nsnU0nCkA9NRUBzy9MLPq3qSi4lM4uX/yjdmQOdAOGl4LrBVXmNP9rBV1RpWNxOFq0OIkgYzBPsf
lHzbEyz8zu2bzDpz87JB1Gf2vtmrOg6dwtMM5kBp1V6m3qtyVr5W8sTxDeKZxSji22fIizcEvIjT
iDN0d5sUJk+a+EP6fA3ahAu115nhcekbRAb75VZMCOgje4kpXu4xdgDM0dsMn8sncGRb4TnSKgsP
qxCUJvuTlnVvfreil8wPZDz9U5/ZBABgnu1cE6ZrplbXk+5tEUF5lWQk+pnLeaT5kOvKZg9k347b
w/fDngJTemqwGh1uylBs7QeZ5K0Tu/I0ax2EcPE4avySt/0DklStvr9eMAa6dfpeTP3uXv7qmPpX
T3OBnHl3cp7Uw0S6Tm8TatLv3LqCr3fehXXOYMW3HW2zKSiG/2PGpu01LtgXAz1EhfjjXJoniQcQ
7Ofl7g/2wZivuCu/hYGKhP/XWabYX+K9HASDjTqGv1UXwUmyVtRsV59tVHh1QOe6EeHW5dRdg7GQ
u1nUket1RMJ9zVw70OSWLY0rOYCBf2kpRGyGYw8Spi4Ru7R+ccpxLjztd0bwlYGTzGppAkljrNrK
I3yFzLpPuMSa3Q/t6nwMFOfDLCqZkNlsDl3uKWA+Dl2lnvZVazMfxvzNUu8W8VbqVRoqMPzdUa0R
ivPu+hHcx2jAfNj6Ra1yU0UO0iopppg6zoIeVqv1pmUtKKFmk5eSqqVMruA/WSxyAPuZ51kb1DD8
NbCtE+z6rnJnlKLxjvf/cLD476xNd0PqzSM5tWFzcXg3LVhv2nJl/Vko92k/AQqWdnxad/0PJjeY
zV0J49Mp/il2E2l51MGOIIZTPlxNQBpPRJ9uXVVCeU4/XOl389gfu+9RUZOCgXMWCrqwSQVqfTK0
1Lgxkea8hRMub0yNFuNaNuSjbrR06iIpD5VbQGyRUO1DGl9gAiohofJsEQenDAZGjQxz6GtANugt
f71/qG+UuNjxYiQEjtU2H5L/nZOIySuN+Y4eZvc4K1yXhdJXYFxRDhRA0nSBCijivqKJXPZC9wuB
uTCKUfTxg+tuv0EkRuGZAbMwXApkber8ZprazZiDaSwuFYERPavPJUzO0hJrA+w2LAw0ATMkaszD
svHWAGA/tebI0sTYptV8uQQmHlaeL612DU3kkPNj9uT2CLRQy9xKRvI5NfeR39PGs8u7WmsA0nTo
HbcIx8H35GcUrZE3sOS2li0gIDPjMnCQhGzBP15iACVGb9WlG2hm7KUy5yycGBUONJWYrmBqJ/yb
exBGZOPRtcLapwD+M0e6XrWt16hXjPz0vktffLHa2CnZBgEQ2+3CGTbBaGoin+Lrbx2na4EGJzDv
NIknw/iD1rtHTHk9ZS28KV2mf+7BIn3tc9aEXvEF+iU9Vd1xnQkTB2Rpdudr+g9V8jdfeZ9/YfJY
HdYZppeMg+Q+Un6Arcg4NLP+Zc9jx9EVTQlDQs6jSxn3PUG9ks9SClU0EdfXcWKdeuJPR9+YWZl6
grTxzqFxrKDWT7jVHvvfBulrXzLJWBHiDs6OGICKLgaBpYMmd6WmfKATEYa5NiG5LgWL6w7eM+bm
4fV8D7iXRu+S3VtzrZmGqBurPcV3IfZWhj9OL91J8NYWctng9AILHiBBFjvBVTh+yUnacD2XSjKS
yEemoB0emrgrjF5zcfDcqtcnozw8wt7M1W+GzxjG+5BGWABESg0e/4H/3A5LiF66IdrD5HBCPv0z
X7lXnhfbtVBOheMhSY2kIYvpR9ek+eYTD4rDCPd1h7mARz1nmXivGDzA1vb8lKlxLdF9/TRtUodb
F4QO9WgTRh8KkEMfZGowSgw21TtiYvx3EE4VvzdagctMK+PJ5B2L8uyMicFJ/DVSwb30GS/16heF
Ybz2AIDH11hddN4YCWlhCRvJgLNmFGwrvfTA/3ywkgLTdy06CysDJ/qx90DrSUHIg8DaDP4w7gd1
/eZwJ7Ibm0E32M3TfqPmKuj/girPHkhEO8UkWwgVSzUsBqOrc8n/m4roY/DnSMa9ruxZAmbCh9sp
kfwDl7igdkuNuk4NapkCzUDU0KHYe0bjZvZ3v5tphAyqmkY7NO1EDSvYpme85qT/exJpv7IXQlH2
uI/UgvwcNPWo0dwkZp3as+lneY8eN4NlKkaq43O/DKJW/tOSBqiVOXe4D8JQLDfoVZhjIGeAis8M
cM2M+R4wEC1Si1+gaxJxJWY5dyPvn5WCrPXEObt6Kn4GlC0dsxe3NWdYdShUCTQ+Kjao1NWzJGsq
xVMpVF6+pLcItRVzwtQzmVnsaIsA2XVbqrxxrsPr2vXQedp5ylCftkbTV5Bw1lrp109YiOvA2xPJ
PcLjCSbCB6sS4lyUzvG+xAXABoxoCHLHED7AEgDG42P7OdWx/HVyncY6azgRxiziL3i8498oWwBa
GoQSrpk+pn+hT6LFlQryzekNGZHBSeD+OOj2Zsrcy8smHmDGklhbD/+Do7mQSQH8S/fcOuBpScWL
uJIV8rdhlgoNxPaLrkqPUllb+RRirJFe3Lud4ybyIr8FZ0AiWSqSS6tpTXB8ftsCBhLXUD5ZCnZl
GLRpS4VR+HUKJcCxKO96w7e3/Nw8K7RuUw96zP8KW3IYO1G0XC2SWpKWcnpXkzLGdmpG+lxQVwtf
Z1poDDu8bZqrLlFB8lItz8yiQdTLODldYaX/lsk03L6Lu9bElLv2YvOKs87Kl4u8ohi2kM4aCCVf
IbQFIv6vp3CaED7mjTCYfSHgSnPug5gNkH7ZB4H25UyrbNZlDmtoJihdynnspDhX3CCDIgmCnLPS
oU5PPo218s9XPhK0oBhpsSXoDiTWZJJP9C6VMpOgKbptbTDAsjYOx23fZ//AuwE/XKnrMAoiPDrB
IfDQBFM3Y1uQh4+slQhTGqbj21iXoPuUH+QijQSHGUUHAT7AC+h82DYI7wLyvoQEXXs5C6Z6u5UK
HC/4FKmQjAKZuqK61Xuh6EFq2SQjlW9BQ6jOPT0HDHk09LjvgZTXOWc1y7nmIHJT1hReSYN713Tq
oPOElM1ykNOLfuuAFhyR23HYfjbYGn7PHd6tOz/kkZFArz5kzwM5gLGsWumKv/bKFAH9wY9q/k6r
DVurWFvBqNfMKCK3ArnChUqLCEYvUFcqrDZ54OAh2/xKot8gBF/86LfSGPFt6NVLsvGp/YIvWEKS
z3NNUc6CEmCeRhQV4AV0QyZ4gDEliWV4GSiQmm22QofGvHWEQ765DQ8kw0sWbYGMubjLWQKJW8JV
eHjYEnX5aZt5w+mJ0LA5MGx/xCUwEhrO871p2cGRri4+lCFSptfiRq+ADYOJEryMQvCA8n/ec5v5
/6PCYfZLosPjlsDvplBSZOzeQxvzO/o6YqO3LEzHxVe2ByCnPGBc/HLx7Ndsp0iXLWoxHUzZ8JHl
fPYnZbPnXqUizYxmWzk5l7cu63rLtGhQlA6xYeMbCVVHC61f6ui/7bQVMAT1xLTSb5vqm5MA1zeD
TIG9Q7bX5NjEGl2cajJiVOge1xW5H0zDIEJz/CpasSGLtTvuXRl/5xc9xkGnQBh56ypkfVI4vaSS
05/h9FxcYpIo37XH3A+RY1yDyxXlLfYPEJPD8JvJyxGMrW1ZFCbppEHMiEG3xCuu7wY4AMDsxHNE
3emSnLo47Fqt6wvTJMLV9x9fcXskk+ZI5SwLxT2hnDC/r+lA4DDPTtHRlZ5mCcxtwNKizVH/H0tw
8Bh8w7Y4OtwYyVG8O4NLU10nKHChP5qb8RL/2I4xSXa0fBKRZL4hLwmPDuzEnDVTEg8FIEjcjvTQ
tLlGOq8IMq3EsGy3Thgsh5hAqhrHo1fRrz3TX5QNJkCTfBqkue7TnKp9q4kiqyFHkdLAURKVA3Ta
d6Y4+QtsOSvTSQI29fkjCb5xo+JzNhvxhuaT5cJ4wAeoCVR1wz3QFuAz8HKlDyinCyhrqwBuSQyT
zOcTKWND1hrONMHwRZCHWVnQgjwtj8XcZBsHlsFmFspRtZVE0qCdxFZV4m6V6T9+ZOAXzxQ/8jPr
sFPDiklDUWUm0cHoDa6G30dZqLPbrqlj0PXrPB6c4UenBGxIrRUCFdpqVdnK3pLqX8ax0kJyuji9
SQCselfnYUV+7XAQeNIyLCyS6/cyPxpHokF1Spdvj0S6Fga6utrxb5uDM5ygnbxYwN+GDD2aXaL6
5mZ/BsDlrh63uejqrprFl/EnsyYDxKIXAnSmf23PmO2iKPoeI/BJ+u3yqwRb0osaVe0kahcq9sHp
mH8EFp6JB5zFloHJiN4AGD+tzICYGznX8amyT1AH4DaVCS6J+zdPFXpOFcl/fDzqSdz7f8E1nEFZ
vzRu+Z2/8ZabogdZkWqKzZmepvcyrqFtzuEdv3klnt+TOy4hGTOAuYy74oU8jniE5mLNNb7yc+Q/
A+VXv7kgUQXnMjB6rKYoTbBJEDfGcCQnFHMoPyRWC11UPbrRHThF/qv3UnlDI44r1Z71uLIikMdv
8h0Sq8kgEutZ1I1NXrA3ooSSNqZI8SvA15YkBFQvbmEABANjQMf50kDPLmpxobvDwj8+LsaXk1cZ
W/12ty301zB4OqczpGCGN4NcFJwrlPsgCqQrmWbzj9d1tRoBvmaczLE7x+JGTvoe9K3YK8K0SwjE
Fy7BVWDRPzjFrhWZXkfPoQHKE5cBEpVqtKYu7FC8vPpJEHNrMiJZ/YF231Vxa/GYAtvqjplRrtOg
Cz0CoaOiKxx9Fpmbp1KCuRkUZjLcT8BJXK4y/j4FRTBZXKV1NsFLnq2jQk/6Ry+YT4cUWj6wjbnB
ZGsuzB+8QZjLyOx5mT1em+d0wMFniBOCKJnbU4E+7DyjEGyTlxNfH1aHDUBKtYOUoSK3TW9e0AiY
68OrkJQc3hFwfXUxmKeG/VNPNKnh+syDS2y6W40p/msrYbBZjQv7epf2BFPuLVlaQzM7nzw8Yrbw
5eXLil2PsrFxfTcBo/2pCTL1otJ1x64qKJvB7nfloktyzM7I1rQl6oTZB661YQ5jkXDebwZxOa4s
wxtsm5QRP0ZLq9SQeJebMplMJX3YjRPxT/HWY1HCBGASMJ9ODnU3iq/flcSBxd9eQ57/2TDdTBEZ
2rQTUfiZKT/xXiwhWYxtRSVZAiom57Nmqcis2HnLUPKeYDxWUokTwi14DkefoDrNp7yIJh/fna5B
7hc8jf4SOTdb9ZonkcZdxa0GPRdE9PmKznS3xlVD4Q9OGBbNMP4s/B4ueQljuypBnK5JURo7k0Fp
zGUFnrhZhill+TmL7GF8BEfzeeneVO0SS2wYG9dNaQ+mZiY67bXiq7YrNSbbDtBgeSqubdadAIEb
GaxYGizF0aRkN+YLV6CdpomZM124exK1tD7QEd3kC/sF0g0kxQbKj/zyHA4P4P03Xn0aZWD74iOd
IIHYTXyZ8HyYRsTKZiUKgesQOoQY1ARSPBTfL26tCRrbGWmRU/2j72vInbMwoHAw3gspAIOKmhQH
m0fY+SN/8crdw03X42IN1QWuKwJ108OSogD4rICRA3MBF25tiPIvdFVXvEDkk6fvc+bzJk+JV287
BY9EFO//aSCOdFzsuycyJXpc4NjjpF0i/ciXQIrrRCuqd5YbnCi5hZa8a9v7o8tEA0dwjLZbsyjW
s4xRtL1GMo4DN4Z0Vnce7SI8+BHSyNwYfPHwHLTWEGEV7q89MJPjDwJ9Mnuiil73qyZdiFY3+bi3
jW5miBApU00dnfzjn0xCoBJ+u6Bk1cgxIfDwBBKZA89XrewPwmJfqTVEiACw5Q8ZY4ninp3AT7IW
gIlesHtUmfk8LuPBcG1G6XtwiU++p7iw+rielVVLmCOQhnv4vM/1vxhduoeqC+0Nf0FO66Quj95m
A/rS7mj7LFkY6yl1cHeN9/mw3mCmMih/eI1X/RkZ71PF5CAodFZvYKQtB1MniAF13NzxCjp3aAOY
JuuJZzx1XbE19iO3Tqmy8mOGPKRSaJtvK/NL95NxpnG/xlsSIyDxcKpBi+6a5CVsBGVEq5MnRI0b
RkDnb8rZLSBMlSU0fd5WUiSns0j/ZNTvL9DoO+OFSsZBze7HZZg88zAyFL4mGkeRvRRRthYWhSVm
YdyOuEd8bo6/m3OciznxH0alH7wLjQ9YcJf8ZxN7pQwB7reCT/wmz7I0YkcOsYIyubwKDegDuarQ
ENbqIe+7Tl47TXqabbLY97xLQ6l4JJARbN2f4422HmhlHSozMGBcIxWNtOAvnXzNWHLDSWwZJEz2
VWb71mnz7DLSF3+bY1w+BbKJ3T0JRNA7WmXsSfFLym032/bENr1hPA8vljFMkZ2/Uf+oRsIF2rdp
57gOd58iXbsB6bH8EZ+gT89wctlKtGT65mvzO6Oq3dNXeHFoPBKtDCYwPAaLJsfjcV26PZ0uSFqQ
XWivZjOWbpuy3JGpMrSzwdESHnie1i+Aq+bwiE3odb/dMFIry9PGVnaJW4biPU20XX5VJKzsc54d
RvqtuG52tVyalM6KVv90IcvMdmlz5DuOHlHafNQQRRGZExLIjHUU69vzeRFFrMCaQ7S0pD8ocp/x
aHzsoKMkhaYS7hK8fdTlLhpGP8NpOtzQ0jyecSKgReqXAtLJR0OOJItMDgLcq+OJj6ED+W5/hnXU
qfIlN3YCPhCNXRT/zeHDMHKS1+/krVvKNe3G4DI10EouT1nI37e1gvHbA1gehF++u3daggFkX5GH
LJ63twdlPHOM62A2XYJLxOe4HQ+wN6Eny36DEji+7oHWST4ZsGmkss0I62t7CelUtwarqh6hoZVU
0AliRe/02Yw+XHtO9mcjGLg5BRtRUttTtjFPUy35ZOc3p03q9NI8YIhb7thxiVFr9r0+T8eHtJxt
Y3SaXNeC6/aJzjqz7qs+FYiANnxnQsfxPvKpRlwLuQ1jW8Rj+EVNlSZzfe50aOjO/oGOXCNSo0kw
vPkNi5FE9ebD+A3DEgKu2YsyzlVFTNtYZhn1CUTNGgbsd1NFdtuyYGrlq7vTPBmQP44aHnIrJYU+
2NgDJArUToXcrnIh3+OWCFRYOxj43xw2ut2dUVTlVywyhxhToLkkshXy2+76l+AM1mSzHDntuGJ7
aWIWCuLieHYXNaJ6ZzcwkwBw2WCY7wIKvEYl+EjQhiDO7lWakL3UzK1OSl2uuGtk8txaZBxnI+HT
MGsrYBXDisqnivxWONkJWvrWjFRltXRWqbI+FFT6zJIqWeV1QVue1aK3FV2DMYpvURzylRTMxDpz
SPzzoLjsiXrkWrGvuyg406DO3CL0yM7PiSBgsg2aow/yWYWXW8hgjp2iGmwOmmgjw3GjbnikmZ9q
J8vYoaJ2xIPJU5t/KgLNgeEQNOw8Yi8RR+AMaoc2r4420KwukxN98oBmM1lVvmaXr7GQjT9OI8hv
KG+vYJySWNnp0PD51dGyWeFycTQ1wWcaVyxO4iHCxliIdZzvYR4jxYpQVWYKMLtNT74bnJM8hedG
K7etFBj9LSNeRN2U0BShqI5z/2z2L9qL3oRM6Ie5e/AprYSnkmd0KFForXD9LTxTNGlo7Ni95aXp
Pem8qPR/MEI8GaX5ssUfJENmWzI6hWSmi4loXCcU/jfmBv2Uq22JYF5aHo/Z0NsqV4Ke4cA1q4mH
nECDHttdelzYBFjgTdwjoCmeH61UyVuSRPFLlFVBUM3IfmbBE9gcZxdm+Mt2QJh15tRrJAwRcoA9
qO2zq6x1eZZ2X3SvTx69mK4KUfj3cVSWAZwFId9DV25MGNR32OrcMJ/uYja6sv5xQDN/wXGwIgQh
MalocpoWhx6nZxNbgEDTVv5F7IUPM22KvGIINyYWGELX/29WoVaxfdQ5dY00ZbDm1odXTkQ1UH46
A7iQwa2UiNh8aBBkUau1jfxsm//s7kKYOO20H7fBkqStM3su16bqbCz0EiaxfcW5dZt09nQfZlC2
rrYzzawgBrJkp5XQFNTSiSCFOMgWF2wpKHQLm+6spLo2oFEKPI/5KOEVT7JdcTNIJ9OjIIKhpGue
JV89uxiCnr9dbAm5DGBw+ei5HDeSWhqdqOHnp5KCMvAiyOkCpRFq2NyARBlOYceE+CCkRtEkkS1l
TXJrObRSZAYCPnoM4eASkzNfweGYELEKi5hJmrUthm9ka5Qrpy+P8576Tzj4oaM6YW8QunarvCG6
aZhBS95+JuBhlLkaqRRTnimpT6mAcsHhujhmnuDhyRNSRrCZeNMIZEk/jtbDC26+bVlrJSGC93ZL
CTe244YMrSx+bBzPqwbK+oLOCGVBDmq9fnDckuBnaJTJzX6ZzMsH3zS4cYk5nEbPWhnDyGNc/HEC
kcLUdwwkkYavOHHbqI4IjZ9hh1sJgq6uSivBgMdRaLfH+rcYf27bMhO9jypbSbJojnOFFAdRhSjr
8zR5UBWFWWvzlIu7DC+jNCZyceUFPsjOC6Hw6GGa8G+6hKUrcpljYn84E20bFyHk+T0gEKPuuWbu
nZ6Ca0KdDNPZ8gmQkIVZNjEn9Qlj7k7I0an2Z2HKXR6G4HUBpWOqTFXw1fV25GisPwX2f6Oo6b0M
ob89nk9VUTKQ8fgpsT4QkgY95nytT2asU9eIEkP9+4ZnuKAcEC3qGKniefvUSYufs6y5AzX/o6a0
EuGlVziu3k9/+eRwQYk2T0E+KuAbHH9NsMU+kRUhz5n5oKk1QnUyo9+wdaZgov1OUhEIqR7pzM2K
MjLQWenS8bGg5PxFZfkjyCaKWs0PAgRvWxcyfzzm9oionf0AN3f7qPLo0YFacLzBDjuXgZZvcEvC
6Yvaqc0tr1Cz/Mva9KABhpHk6UCOE4K3EsDt/gK0yIlyGqBXbs5O+gWLJPtIDQPWXFkrFPPVwETY
db7hhtcDsaB8Zo2aJFdtt63tF68213wcWw9KSH8g6ZPXVdccAXL7mzKuvhcTNHbvbLid2MdVle2Y
Hv7adcGDQ1SnoL9tkDuiol4QLKohy5ymQYxn/3p3p6cK23AW9JwqyOrQJK0gpP2LPNrpE7eZtfXQ
NfY7FRUoJrz67uuVYIQG5XMOscAZRMrAVXmrsJiUEKSbozb7VhN6RlWq+NccJ8CLm6zykkh7wBBt
+is4VqllIKgUIily0GrMkwFhw27VZ0n09idounbzL/KAXuFuycweuer26d36iKoR7Rx3RwThZZjN
yY0jlI333w7LqSlX1WtirxVxeU1FNrlz13SeEJPQzKAzAujmkuu+ZP4cDv4xw43m0cmEelyKHhzg
yECjjaYDPNteUdqjMXe2CGhblrkXscHQwCd4mduwXzmAetVyg+7cuU9aiu5DVwSWSsQf5/t0VKQ0
U94rUoXfYoLe89CYqIU3/mYs4q87mhOAIqLmbrcpyTiGrJR7FuOwZMIMzhpsD/NjhpaJfwRotT8w
7Wq9PoXrTg+OCz2qJCIhJxJLx6ug85bgVk6yIKMOhxmkSKYROB6Y0I6/eZrqWZEP0vzvjRZ+TE2U
YqfiOO3gpP7if3hDMD2HB1JqKI30trlhYETAoqQan8xPeZYAcgLNb8rdZT/YANCgV2WyCN0SnDXA
q7Yh82iXh7GscB+rzt7myoUoh+IoOQN/2b79Wc2GuegdF++u42QfsWrQYO+/IlNEhmVTOO2CMdC1
ie1Ycvv/FALHjj4Cv51+kE9+lh812Sh39S7vmewqjVNO7SerWXkul1M/TCeNO1AiQ+NO7znHRz8e
aqGyCIX1iWd4Ig97VLr5csaybXzqyL7frzcb0IGTIf1iHDeOyPdlskE6E41qN0RShBdS38iWtv2/
CuszwYcSpYHxfY2NRtv25XK2UuJ5O6/YVmnXlJvrO9qh02J6PU+su0ptbca3oKIs+jpMpAYdMu/n
G4+BhvI0DQ1/tCLmViBTFPTxrN7Gvrb54tuQ4Q4POQH2lqgzSR0PPJcJUq2Ur7Fpbu0VPLYDb2wN
p6mOeep8vCK9kf9WEpOz3PjPSNOWsExeyaG91jKMFJpWu3qJ3n1FodAra4BnLpCqtYqh35e9c5NZ
GJ0/oq8icHB6kAw90/cWe5t8gcus5b5OBO73qQBTNv5Wy/UST8TdctdSuajm46WiNHo60XJqPmkM
bg7pWhScPYNhvlxEjEGAjV7S1wEQGHHL0+QkLgPJ1KM6ymzBWiFAL0iVFyPFxlQuAk0/wzjijI4U
QNfp/sANrWNO1pOYVXidaN7AFzQO7+r4xJNh1XDGyxoP5UBsDsXXRmTQ2UHfTaiRMNb9QgwX0di9
biSmG2TaF5LsZatIZQPKi6gxDLj0U4JoYYr1CONyHyMmIySOs27/VlRmhQtA8Xm2WxL5QIY/xiHq
5N3p96cnUJb2cY8C3yEbxovy4Vn/BxeBlaCgQCpWBXfl5mIBdvKe3W3m4mst1X+xf96HgwQqFN0d
Yn6aNj1NHsBiteYoO+vab14pefVXpqLkHS896gtL/GW47JUUzdhaA9Kc2Lay40AhRXS2raWAqY7g
WL8n+ihN4ExfD1jW3apxOLyohUP6SxohLeJx16QG7M/HcS6xQje396QnqCCtzDOZbUFWiztTo7cr
WqCjuLz6YkOerLHsq45LaZ4wJ7cR2QfWW0x95M8ReslZaqci2azoIalUBHSzVcAEjwg+nQxVOekH
IZFQeUex9xpYnIk0nQyNLdF/LrEkfdfpk3R3fFa8cAXSxrzqAPLBKBksfv69pPa5eQYMKiUpGFit
GAe/O0knWrwnq4ekC4Z+//RpXj1jW1mIv2pwipHV8FlUVbXMM8af7Zh37kjRPi9utGf56+G0eZ4+
pKjJqoyhN3EYVjKGf9vkv/uKsAHbhK4mX3iy7tK/A1oXS6LdEwqA0RVdR9Hs64LjI+bBwSWhmENM
Chtdum7IyuoUk2/iMtP+caTs62Pq8qp1axzZQkJJcEswgRccp9P+Y3URz/GJmq+0sREOGzOjpVlx
PucXofC2Gk4MGT0MEWrSv9sdM/M2izLq1Y8IPFdTpLyjHrdak1s57RTh+JptKexiJ8elrVn4jxFC
5jVIyTykNddPEezbXbGeARO7oHQ+75rWc+buW+EpNoDyyvomNSnS0wvntRPl9YS6ZqoWwX+5gnBC
1EJ6fhe9+rwcHdM/dIeApaFBzGVYQxrSBD6oKr2tvgyZ6QjHpCIjTH02awe9PjHy8cn/JENwHOZB
w5CMiDIj1kKYZjD2eu+QrOFvNW5F8f2RV1hwjP0gK0xKUQb6tMLdfj2GDYfgWV+LHK6uBKp1Ttu0
DWionGTPRjOLjLCyK42vysaf4ysDqIl9A33nsGQpQJUk+JE1xgBDi8n8qzHBxA1hSNytMP5JKMA9
wsckstFg0H1SLS50J0F4VaWLeHbMWafs5GM5uKRz1/j/oUcCQUKmmzNjnNdxS0XIbObtLyPSKbkR
+qPodLfMjUbFhlcdYI8sAgvzj0g+IMQ3GAnN1/S80QwsYHiaYfr9HZp59cBqpCRRN2w5VB50oupj
n/ASWLjo3yIwqaNv2m90vkXDy47Q5+NmiX8a1WKVq4YOYHkwDtl7ChXup9ocC3qj/OasQc1vQKZs
IWLd3bjRS/Y0xAYFXAb08IxAseyauKk4SjZdolOUAzm6f88BRu94b9YgSFPO38QciCUriLSS2hao
KDT40CUGuyLnfw2kasAfWw+PShsqyydOMlGuohlZ1rcyxeLB+qjhf+mEBB2JrOKHytpbDIT1R/2q
LVn3scNp0qb4oQQTwZ4/TOW6E4z+MxpmoAMIpgyELBoYgEahuJKbrMYi1UoQNaTJiWmml1OdpONe
TYmN9uUQtMJvhi9+h8ghEXnQ6nlk46qxTj2rlICMVNA0LKGr9rD2g3HH+CKxDFQW+Lt0OAdb8iP6
neCMlECl1v90W8COmNFS4P8ruUN42VKdXSSavUCYUMDzQpllfCTMOhOyd8lOtmsGYBnP82A5ioCU
GHxO2hEgHpOkbvTqDJpgpl6bZSizAQliOL6X0giC8P65l++hES98I1Gc4k1/nZ4PPeuVkQA4dFqv
XyYVQvHTA33iJlHetg5UO0+Nuws6Ro5IuJA/RFxXRXUZTtWgMkFv8iEls1rH1cTcKJobTEKN/pqz
6UxxENrsZ4nnnJeECcNqurIAsuBPh72WFTNUsOO/s5n40qIQcyU4Mnhs0HmNN9omawtQS5DZxuHj
wMkDbI8I0y6vOmzOLvudHOM3DIi+W/J2roaX1bQwDHN2aGKnI0Vwexuov2e4yzq0WNEK7K2okga4
OiB1TKR54OrZc221r4BcQ7vA8H4leoyfvxQ1TCi3+aYmuhO3WTRVKAmMIeNeDKwcenvTbUxNj4eL
wLEDrhgznOHbs53Cy1i8xuFGI7S/eQvNX94OARxX+CRK4FTc0+BU78ZQLHL1PMy8iY0U2Vdne+M1
3SFBrFu/hdoC5vGS3aGMOU58qoIyjI4t3dpqonOf898IBEOzpU4DjJwn7UMJF6ceQvXmZ42cwziE
CkD9804nIgAwhgfNajxawIBKCghVKWOlcUcCRUeeBbyv9KkhcaSa7DIpzw7zVdjomvT36Obc3Kp9
CebH4XRmw7zr77xYEQMHRbs5r+Uf+4rozMQtdq65cfpGKyYxekJfRzetCq0qJGFPwUtTePxqKYUO
O4g8XgU74YZxb4Fh91KXxTBIyqWulkUHShuHrAIEWIyMayyd7NKneDin535jZsIWtr5E32kUag1X
0Y/6icxEzu8n3VNEmJIIkSVP7tKFq1RuwIkU8U8WbRBQUu2XFMwpFuEGokEzj9hHFlB8Fsb/8jW+
GI/CpB/zRwX5Me/iIxpHoxQkfcXu9PaJeDPU1+z5hkqbNrBjnEOzJat3EBefiy76qt2VDToG7811
YyEZb2OJfOslB5F33SPLR/aND12SlN9ajizh2ZymX3HbeyJP2zDlzOgfOlXHpwFuNqKEvfX0YW3/
cxtQFSV8PTS9MD1DjomJ1XDaEcpy45cj9RKu3CYOgYW94KXWFxkXS3J24rlBcoLjil1qYpr6MflO
qujab/70o8Pj2Zy+ORpiWFX8PAbSVkdniNtmNOcCCumv5zKhr7Np4w1G8ybVfWEUyIUYPmDGnVqO
SMw9ABgWjon48wrVWFuIXPvotOit+SKDNF8wgQdGRoNyJd8Z+3raSpZsji4h1K9/K7sxBHVsPz2g
bCPfVC5jtwrP12pwWxgL27ryzskOao1DsQuqcB5Z3y2qoCVfuzQs0jwBEf3oVfeyNygg2NnKwiGd
EjFLTqI2c+6WUP5BMnqg5xPjjViJi3CHwg125BsBdZLG+WiEefc3lwF4Bau6ucHfb7D051HTIjWJ
gogHP+J0E0Y1+bLQinSGw0eLnJYFXfryQUeJ1KdZYsPaOfSDvBhItZd3GeyqtDIT4wiU9L8JZByV
idVSq0KblpskSOxa0Orp/cEhHo5TZD3bopDNzsiTa02yo91oEQFeL+Vwf3pFo+YEEpdHGHsn/LJC
EOmFP2LOMon0J9EOzkpm7EowgyJ8io/xyYEt8X8HabElDq33pbuOf5DM/xIipfosl0ofeF6qXzCK
xN+K0Y6vuvk+dNn3AHakEocakGr52/3Pj/XwTY2NXCwrsjqmkBQdPVWVvFAHUuidwaAlZmzGes7E
zhCS+1W65UFBR0cYTDw6HUldUW6/DpL+vPzAzZLOYv5ZAu4djqxlCYVE05B1EMiKDuw3Nsco1kND
OjbPkMxPFj1aXfnT6BVyoduGJgyW9FDZP5HxnwcvSJF/bum3szKVZD5ZXNM8eu44Sg30UQazMS3w
lyvZQd2mQ4aeUuV//T8akt+0tnYW1j092wQ2kTqKHRBLjIyTiO/B6alr4dv3TXS2kXwMcxPiEZee
gUJoaW7nPDn5YjV2QCGOa5X3qOol7QhiHIr7dfaGXTz1pGVF+Syy9AqOEh7EacCbObaQufNR6vkA
eIrhvXUvnMdoqrfvcjJSywWu5cZOEKdzUqzBUum9h1LNlOchyCEj9CnIGyPtE50dvVKQECoMRX8D
vjYuGapsFzxnxcZ7N6VhjmptSZ0Fu/DJ2p0VHeeyMUYJPsONKjxXk54zKp+IKCCf2ZLUppPqWWmp
W+LhQY1ABO8DnLZ/8ssfGbVD+5MNDSFuFByc+f26bVHEsOqc7PAYvDtLxsWDDfyaluc9Mtq9EMuF
QEHodjaMVBiLYBs/k5IAhTgZFtdUD44obTMJ1jnwUe3uTE7032sxBXy3xhqEowQZtuBJTOciJu9M
5MfoY1bZTH9M5/KzX1QYIkrXs1DO4QwN0fDn2JAoh68fJE6NPNikjyVPnneW5U+B9P4R/HqAlpY7
Marbvx6Dh912YXOEFUntfJbp+R3K7HjlXS762XVMExtSI1BHswoj8kUmMQc61PmwaBkp2DO3iU08
gSa+1uTM2MDqVGTvEjKlXKXH6zLdw/v16nYo+NJf4jagqpBakBLx/0vIzLBiyjsEbu/cSRbOtjiJ
MN7aYEST9RMTdIYjO/VgfJvW15okVXosu5HfITqpinI+5u74TKfaZXdgH51jflHzzisdWqNtuJ98
Y5WypMcHkG5zOb1iL3HuTHOgEXN3iTTb67XnWN60FQXISMRZTpVKlz0TU/1ZL5Wg6pIFm1hHShU6
oswl4fDDp9yZ07HqgFHow6b59E9EDp10m6H8w/vlpmy5e0w67MxWJVQRHakqsT69QXbJjfvn4TJ6
+OVbVNKD7mfLKOr9obg2mKxeRY2qqzsfkBLgRkk7JzlhouTPkQ65BicCvlJEOJhqeCWg5XtysaTt
hg00sR6tGHzkAB/F5ZpGvLcHHQHAzcPdoIC0K4oHZLSgSFUitPU7+YBSx1Ij1xKHXxAWX1lJhfEh
Xq/zIrDv06n7dwxIovtJ07NX9RrBMgbJ/7dL5J9gDQvkpqgm3GxgZM0MXYmxoSEAKWsN1QcwiBB+
KCp2MmrrqI2n7EBCCdxSoWfa75fJG/NldoJ67bVxouXNikIs7kysnUMnHNPCTTD8I6UZFoTeylN3
JISPM5DOiYxErrutxw7Jj+ZUttqO0uqCeB0vVedabXk1BClRmaI7V6Zqkn6MPz1a/GrG+fjWhS91
NFnSG/6wouRulDAvzRm6oRvcSbRsWWsn3etdlCguS4/N6XHzgwAB7fImrzWhYDJ2AOSs9JuwiXkG
vxWbUcm+56vVxAK5arQbQ2IvtMibbabGnihFxlEm6/Pg6hpRPNR0Bxjo08P2HtGcECwD51F36ROi
iWVotsJ9ZhWdAbaMAVonEKg5Yvf6ZxpLFKgHDC/MTyzgmGI8udZCpRcOo81zwo8erxfSJJ9OQs0a
4EJnAg+LD2tTua5EihITNu0ndlljVc76y6dXWf6kxkXdPF1LWOjLgNuTjW+ZZWh5BTbgL8YI2mOO
JIDJCpI3rzyT9jVaBCJ/kSrBIl/hj65nw0KhiD8kOjwPUyD1NfPAdduR+2SUL76mrT8Dln1iL8bX
t6bxrWcJE3u5tqnfQc/xCWwbdYgvyV59Mpiv0Fy9Lw7UV1Jd338hTmZebpr+8BPw1fGO0MG331XJ
zKN0cfDDEeK+yotfrRNHphB8HgbeInG5Jiz4A+3lWF3ZM1RxB8h6SdLex1jmNkv9MRnF90lREJFs
/XVBdcsWww+H46WYsRCpQu2EKdcBPKHNDXKQOTy4iK+U3iLoqSkQxJjMXb2gGnrkkCUCc4XnBH8B
y2I53JcUSI6HGhywihS8ERpzXjLgXo0PuNkKJO5bmpbket+EfFlAjv5GSt0gbKBkl0A+hJIid1XF
8WSd/qAoQCv5I21/4ZAv91IXzuLcvk+vIJDhPeGiilpKYMC2kWjVDkit5Q8g/cub6AeakiFzNB77
xBv5gqYyRyKeGBNAsTo++dBRxXMlZLJL+tGnIEL2JKoMLQg5LTJ9tvIaSUlfTWyDffaGA8jkRwrX
0TDsIewFuxLX5W/hUMp0BaPsntjl0J2NOqQ8eCvQmdW6bfPp3BOqaAHTe/kWxZqEgIEhgq1u2taV
gABlYO8zAFjNB8s9/VK+QJJqjDM6IQFcY7Jx0T80+7oEigMsUyzJeONOa4yvJBZjxJZFOSFsIHfk
Pp6xu/KU6fQs55FFwZibKigSmWqF89+lkOP3oMn5/oh64PDfZQBJuxlUDCjxpYRV84LNfxMEXyxy
w4IOjgXujQD6gXaKnl7T0FJZqAZT2XUfNZh4vyuZTB4/LJ+wbnUv5g1053CJuV9qPnjO23rO3FfM
quxX/RJYG5b04j2ADyjV4pbjPFG+N4S4KVSxY2hwuEzNUTOnt2EJ6C9601aGqxdPcoiM/u5aOpNB
dxFrTq5LWCxfD00zYkz5tXWzGRjCoXA2lfk6f+I7+HEWOMwjrlpSqc+VRAvO6kRMyxNgVw2Ob7WC
ZyJKQe9EOMWwp+YPCCyZccB4TKEjCkAqcgnAJfEp5S1P+AbFfs1CD6a3HcN7VID8/Hj9FJjRzuXj
EPw7m91+5Fl61tNous7g4ERDEhsD46FA3vN/4owsBGvL+YT9j45emKaV/N9J0NVtww0Q3+QVigi6
SEnxeQXqlT+x25gynWxdJByMH6jPdQNj3DewSc33WdTDZYWQWbJdr2cF8d2QfdsC9lqK+SNLZk4q
+vI516OjU293Y7KZ72dY5HPdhlqfu6NRf3dKBGJ2yGsHpYpzWzKE0y0GPv2wv/v3hy0uvcbv7w4x
xI4AO4EZd/YVLBXV4cf3Mt6LUy/DRbbJo7prX2wqpztPWoJtZJDbRpOwb1aGwp0B0oBsLyZD3nBB
jGmfuLHlO3CGwqfsPjcbDQgpCIosqqq2JsZVtt2zHzr+9YJwzQGeFSidsobmFyhcrAnUoVTjyIIx
0pb+UlhZyByful1lfc4m5BYPsk7HIqhWbqcC2Fn0kLObPG46shO2gTCGbTMXEpOl8Hl4RKG0njPc
lay0c3kZJoRPmzJ7UrsH68P7b6We9MgSka8Rm6WlKm3KjrOAnrKK6gNb3a/HEeux7/DG/vRj3Va+
KvfO675SY395IIDBWKDsOVkOoX4Z5gDsO2+Kmqtrue1YQJbnsGXsR4nT2TgZE111m4wMGi5CZesP
QNKHIkQQwoYoYRGD2/uvZAcBw6hYuYrzTkihDz+cuPgdrUhdKiOuZurphNTTzIQovR6Dnpv7Ha1z
Zu5iH7SGsLdubvS55XjH08t5kiimI9iwIs+Ig8RXuGgzb+mid5FBan4kJtPLg+LQmOsnLoqlZOtU
ijNH/qnSJCJoFkrpbrGx/y/9yFyjAhGjZQtrHuwPBDe4zadFd/LwFmp5ngQoZdaB0BduUGfwZG3n
cFBqoMieMv87CQbCzTbpe3WSKyWlvBVTePyI1TackzEIInfMcU488D1kQXGP2iit9LCAUaPLd7ah
rWrs+j4RPdUrsxX2YvIz8waCjf4FoKyJnBPNjEMONiO6NEF5/AFyKZx7OJZTxcdj6sOnbYQYpwQc
KADergPMjwT5UdF/DM6o+6sO46zVpz2TfBm6zAIxCDUqU4kSilVA5VSTa2I0Z8l1GJEg/UJJvWiq
p1BWyh55s01OVXLYKGRoyNJCpG3tUX8jW53gwbUh2mWhtdLubteP90W0I4BULzfPPaysluDphTZH
zOFGM8rluQCnm+txn9sQtzB7iKJCT/MgOw4XzqjiNiWnGU4X2HZEUJpNS0OCQTtIvN2cZZ9L00kO
cG/6G0iB0Qw5uZsw/KEg35xrPQ9wX19CscibY/DESQA2oLpeSsqAQQma86xi1/G9us32wqzEtlzs
xgmAYUGDiABNsXfvW1ylXy/K4r/JTz0Pz9nxyHUxRV3ArwFj6tOfO7QayC417NylDPlae8Zenrkm
74S0Ui02ZQ7OS3Z8RFk86wNUbedWP+CPaTwiXjgRnobtpkGC+crSM/sBsFPvLdgZsW/E09bPCmP8
HDTGQTNIDpcP1EibdpNflGOVdfj1seNtaC2S8MOWh2Za8nbgqBAb01QA+3TlEBqivbnnQ3c2ikCU
pJFPjq3HAU33bWaB32KBv9UNzxvFasbxxusnJUdV8M8XtLTmuzMpQyb4GLSpOLqyIogeZ5U6+1SZ
z5YAbN2xr1vKelG867G4pKP4+rbPSe7DE8ySXBcuksTz7EcIRIbNPKXyfLoY1UM2T6OvHPN3CF3L
2mtwhMZbuXuIOFkIaVSobI0QQSrMtx07G7oIytr+oyaTNzSGWdQdzp6yw69WKf/iEqDHVpyNb7rt
pm35GjW1aU5cP7T2aQil69/l+Lbh8ejy25HlIjmKAId+3ibZSL9ORssQAlY6ekqklVNqkvjReexk
PZF8bZ2KV9BCBnpxWsQFSAGDR8F4StimfQLMhCYJ8t/aQpGTosIrh0O9XPSYmVLsXdUDSZ3hc5kl
P6/1k5wPOWLNBtY3Kp1zivV+GmvSl7Qq8N4Jjg9POBGsZSJSt73DmfzsORvE4xOnAKvEnyHWNH/n
pNrltZrz9mzg+pO+BtJnnqL4IY384MqF4sGWXAH0Td6YCVvQRNJkyNQlmOc2X+caVr6tnY1G7GLH
r7ElKU6AMGTd4udR9wanATos02/cHP2sEUI3neAqo+8t2Qh2ZHmsTVc8a9SekiT2eZHIA18jX/bi
XNBXoO3fTVsyexm7pm9B3KTRTO2Jfd3DE8CinzTlyqWezjtm6C8mMXvKfu5y9bJAX2W+GmkoqJDd
HOw7ApFWVOsW83JJuCfRV9AOXjaOoK0BMolIgiHEV8/rdzINYBZJKxZl0x2oq0QEQELTW6viTKXh
hHzwvI4f70xfAqZ29AnM8c3zdJStKSc8s0qyXG+BA/siuNB4PxmZQjWlnkXHQ0Q4ryNXsyh93KK0
rTRURfhG/3dygL8XYT62bHh0+trYFDMS88usSSc1L8H86+5f7l7Ag9ghEP5BABhWfN+f56zU6B0w
iwMcDhaaHsDPjeYT7hVJHThHkQMc+B8/0gYWJ5iwdxlReM9a2SB1hbcE+10/Eqe5PBbTUIke+3qd
eIgMcuWq/z8QCs63NN3iSIbRCqpp6YorV1D8UGLcaNRRtAGqnAKStxlZaR57wFmTp2tFZjGfuYh8
kON7NlirszkPTIhrkn7R1lHd4ZseiyIMsclmXMtBeG/KtJ75bgf+DZbHZ5ssORgRKkgFrsWsm5GL
08VHyIM4ZFtlO1G7Pf2SlkBMA2rbsv+u1bPFKyK/I0shVh+QFpXWH+CEKMg3XvureZUbzC/LsBwE
4rBmyxonjWx4zUi5IlJ73tyZwoS0PUjll7Mzn7XkEnUlsHh6pgyOoJdm7/S1xixJeOMObygnU0Ad
t2IgpFQFV9z5cKO4xANT55hDWv+Mob4T7irTi7boVtXZqzYTFIFQYnJVS3R6KWbj0tHnXrIe8YLX
R9K0oTJkHggjRWPL1qKITwAPcYL/QnlVL2vP6dBTZm4s7nDUfiqHHL9DnTunDE3Rk2DmvSCuV4Or
lmuZ7eew8aBrJSgsAxEUqrgUbQA8/RrhrxSmkMMKIbOjDN5k96GsNNBcOUAq0mvmiBJmiGrCo8Ir
OV1MoFzYkS0UTlFd30eaWwO53lMvgZ4aiWeTEWxpyB6MBLVS2cg1rqaHo/GAU3rVLFzhGnTdQzit
yOD755HVEyzosfb56seyVJDRb6K7+gXWOMU2TVJ+mruSrzcDHKJ7SorQ/RIPG9fPzikItETlFvuA
sA9MGDK9+Q8vQNvfYfAxg0ZAD3oomBIN83T7TpRZhC1eLY9OnTE7Jc8JwQ3XzDFXBoZQoBq4gle4
vbGsHV5yZNlLA0yVMOwRWrDACfpf8vMr2ZuOKnnmATXKO9wFKAqw6evRT3XoJteEoU971Hqa0z2H
2/elsWmVzgmNjrlLY9jOCUZqrOm2uD8q5qaTdwY2VWlm1shk6hgOsTT+Hbi/sFoafPIp1Z+Xq6F1
PHZkODSXvkZ3oc1pMYP8V0xZ4ad3FVhl34js7xqEZ+PVCbujwf0ujmFxcENXBcazD//GDsf0B5qP
DyQ8w5vc4+OVvV6plD0HFH58xW3rx8OrxDNTqr7sYyH3ASm8ybEd0BhLrHMVYJMWj5tAol0kWW03
kL4noW2n40YUZc7w+sVaRziRzTy0J751c1nt6Zz06vObazuE81/VR4xgKidKBAmKjCzLxKCwJ8a8
n95g8KHJQxnW0EkmsRjAMa2MkO883M78apIT2/mzhXksNgxMSxPgTJqaoDq7z8hjt+/rqWSRs/bl
mSb20ncHYG9VG/egKCB0Vj7aufYoWrDd0iN6JpF96ME5L5mCgJkQqRNcDKHGW0kxno3UR+uEJJX/
Nlz8R2xR7JoUMekvEq2X5fIrr2JCRE8f5WJceOr84pMdIPIgE6QAl2HghfvEbvFZL6sGaXrYi3Ky
0WIT8L4AU1ixIYaf9vopQ5AAxAyZe5ZXbYaNTjy/qpNoEpZ+fGWusoUax79v8s3qLLf8CZbirzNu
RYzR87fkGa623N6pQixMI6J4IhH6QUBgRRe1N90PwqPlc2+O1/zuZoFMs1AbbZXs/cHEKod0S/hn
po6DNW/GSboEEjX64UHSY860ffUN2rTwtoOSKLyx2PLdrh3fERN/35d8DPlGXyniL+hNzFAKNQo9
FcQpi2aS9SDWsNowfRtudWTSKsApsGME9GA4crEaRxUc6kCi5CHrPOH1mCLKoUs9KGF/4nsEIfYK
c2iMc/o66VaYqo9g5tsm7R5KXEmNpO2K4xwYe4RRY5O8C2AOioK54Hp01Ov6B8xJ6JlufgTVd5Jy
NzeDY7H/TkZB5QWA1zGPGmRygDRxtuhtsGrO4msW10+Bn2CaV4G67nEAiZSADqhBq7Qt/oifHEas
YOcr/RsAsD8Gd18EZa5V51xSfsj/u3dOkCuvxmCgnfYGnolw7dSH/ciO2g24hoiQTO2rLhrEinYb
tOjoursWqtt7w3sFyqMrWIATw+eTwpKuFCBBDsza59Y03LXRe5jqx1TqLNEP91qmVYwqGtSz7MkU
6wnvavThzFbGqOHajm2OISgXZfLDjMz+UKwjQt1RbVh9Rbz9q0Ak0OI2lZAYVQqUI/86bGyzQ5e2
1avGweCb4rUGHV7tu6y5HTD94CyIT1oOkuflabGXdZ9/Ib2R4yGPK+Ej0ubSSM5YlDRWVDP2OmzE
MYCKX8E2iW695IaCzsBpt9quWMK6BJV59cw2Z1yGwqqLGbmq1Rc3kk6wQ+hiDnB+WaE4pMYqtzXf
HNqVsJAl42KtOwgNAjdYCKtCB5rGpUfo55kfhHyHWjc/YwAvUNLLRpJgG4EUYpnT+UkfUnwOZPJu
PxXwCn3yynY65P8BsjlDQiGVCClxl9Bgn/dC93CkWLWRXX6zo+30krUzxr7ejAF85t2PKLiY82h5
7PDU+E7xNg1a2Ss2EYwH4sBurLQEgIBNV23Cb5MWgQEnXXZ4AeyJgo38DDNHvdu8UmpnSWc/+BK6
k9FMo7QFMaULDim56Wx3+HfitS1uQwvobc0FqMF5cspYZ/S+oKt9leQh+HoA7h4xYN1bCIv3SGqC
YSmATajUyGLo9YQJrEjrpxNK6HVnqIDcX1NWI37EH5HMY9zftvCDLLDLVox+0QPrmNrLyfXZt6d6
miVAiS/rwtki2pGpl6QfC4/cE4PM4sPgzLpqkAtnLHy8+2seUDKRGa+/yDLQsasf7WIPxXhGsDTL
XfB3aCU91xHa5R9rdTA0iEAzUv0/7CHYNx4XPB/2Cnw3s/pVIFwy+ZuuIdeT6Wp8CtoUYLjhGVLN
zJm4geFZqX5o74sBgm3EdZFiJVW5mGKfugXbwg8skgQdQQ6m/DlHrfSNZOVieOeoTEIlX6eRM1sv
quZtiQSBsWMidLUzNtwVkD6nn0aUvOd5Npx/OffNdB1hJDqYABagaUyt+2zr5z6qbxwT6YcRytyY
cPVCDxMZSdZZpUvI+LI6O2vZcDSpsS01YKgnQ0azDYFF2UVNZznNshGaJcZRagttDkguslABlHq3
cc9f9UDla7IZ9D/cQ8T7yaOMEdnK5aaQQrVX0ZeyMidpp+gWGScV5ZFBF8NnpfYq5oO1nxCEbUV1
IB+VmQUJWHdULFjd7OVmmbV/HlZShPRqK3Z3nzWtGeZnYHDrCuZxHkf9+tDGRwdLB7w2p+bZsotl
m9s+ATszAmI8W0CJcEQpjp0NV4M2Ficw10p8fmRqTYVNC8EiSitkyxh0nQ+O1iB/X6USRDeXKjVk
VQEsBBYosIGeekrus+ZX0q2wIWeZ3OPFKrjYq0iHPwE9l9EZ08+Vi6JZ/BwexZFKutzAbDNvclLN
8bBoP6f/OTy35+0vnkKGy7B1jUdOwQUG6thBEimKRAReqbntD9w17kFnsi+z0QryYKcAPcXslJVc
VrJZMetpqfP4jTsKzQQe2sf1nAkBZ5s40l+sjHYqr3tBLtCbYgYzRDrHZQQUUpzvrfck0d8u5igl
2ItqKU7eAz0U2mLc36830OFRi8QzFpJglHXG6t+LOxeTr+uWzjMagWnVYO4+SzNrzccm31e5Anaz
Iy9tQ2UQgfvqUdyV2kSqhYq4Updg+UMI3x9Wvnpk1wRYy5vDI6gBORY0VHYA+OoCwX7iLFF5adeB
TskpZnm2WDohQMoWmXz/f3EbgQJyQ+Vq36WO8NA/NlshiIw7S6RyNhj5iVfFtKl8klKDAmgfi1WM
brbOfgSV6m35a6kjPIAnzD2Jx//xDfllwRP9AU5DAVzKuoKz3B5cSJ33SFLJTNEcDj9Chia8QcPI
pk2Msx4unovsigq81tjdif16e0cXcGXfesNo6SdASjg3LuQWShPGN7X28wz9Wv8R9DbIWHqyarap
dgqPTuoIODP/lxF9a6Z2qOpljQX3AjrY1XohNwsD9I+iwAsqC9OR1pLOVH4HCzK/geU8ad/p4L3w
l4PV6BN1tucnBuddH23NeDQOpDV2PDdEHcDULY0y8grCPfu7KwwJNI2eObhbOc/I7XO7Gx5VOyHE
3XfOJGglIRu35Hh4STAoQfVXGsz9DgMWjqSa+13+4WPoDVkhGoZiCGcbaeyGnEbkN3asEmbNN+fe
DVXiwpmnOY6VMHkCh/G8TVQ8URpARqq5GDY1Mih3x9aAAQ6ctWly23LU9LF0Y62SUr/SleQ2qoNw
nCfth5G7t0i1+ort5yToxAIquT4SY5cXnXDDOGumLU0mSg0d6XGZJYcLyoi9K+qgesbd0NNnGUxq
uSSjgpdOfxrRm3gUyGGlgJlKAiuVr2PgPZcmlwTmY7qJx13V8xgTgSUA2X/dGfyGAiN4z1G1k3QX
PgFXe/VwIjM2SakiJCioP5LnY6YoND/YYa7O5n+4i7u7YFk28q7g8fXGqnuKH4zkzRBUV/WISX2I
UmwupIksnWc6lYkxwG896N/EDdNLO453fOfNJPsWc4rco95Xj3XHAlFLJB+6WEic4qJ665A+3VU1
GNrDCuAYgHy5hHdJb3CFVnu7Qr5H2NWUpGZwpuOgYcf+RL7nrt0M3kmAhUs0FzR7zKbACzaSegPz
Zr3muf2o/9RzyF9LrgWFawCskIWNK238uvC5xLZcCk9kDAUFzgScfmKBBejcqhoS/D353rJrgoXL
2L96BhPhoUu1cvp/i59goRmquhiNxIqPXzAf9bvEv9XiNNEzmYLiMZTcHEWuxE2QS2H6fBPpId5y
y+MJFey/78qZKQIGZa+ZU+Fj49QtK/t0tkuZDPyJoO4G3+zhxgpL1SqvR5JNjc+LMQi0lxIngyUa
pTVv3o8uo3OnRkqW2DiKEizOLWxmri846SWIJx1iu1FOoS9k59Pia+/TNtQ2cLedhTrnT3qsrw+R
WiV58bDXRgiLHf21kSq0Hlwxt0gaF09HCTBJXkAGfhF3TIZvTFc0NWgg3yKylmGGTQbOJhVoWkki
2oir2kjmcQ5rAD/24e3et1wx6ttWVsozhACyYV5MhgGx7DAs4aThWClRNkw5icVwauxmsqBXX7VK
AS1g49pKvw/msltJsqovwN36JAbCFuDzbP8LzrKs+U37fmpLU4gvo7XpRw8jf21hr7RLo1M3PSbi
z5A4hv2ZRVVX/0vTk/MrS/f8syFtwVD8fy1yUAk6F39hYuaN9FHWkyT63UkGb/GbHOiIaPNDhsEE
iGys97jjZjar83H77W5U0WLbVj1hzBw+IvBKgazOSliB/6B4lWoM7Tc4knX1dAhlJzcuQ9QZz7Yy
sCoUe//UqUv8WipXJ2GMIus3N8ehlEnqTDXGpIQ5OQraPtlDP9vVEh4wdp4IM9L3u7TOMbc4NVfq
XMY9qPJ4Q5GI/ggsVVaritjGiAnCPCLtmY+cS5p6pGBNgBfOMhhSaFpe7KqMBfyY7M8LTl1jNGIg
zW6IOQhRLjfjI83FmD8huNQ9lItCJKbu2gOQRnSm3fQ0kBRHYS782yqdZM4v7nwmxCHE9pgvzEBa
A1UxRdyizcf61FjD/o8cx2i3bux03f5NYVxxhl3+xcMCwk6vGllrYOrXnrtbYq9nfX99/+GxYnXk
L7oszTEf4Jh11Gy8EKtm3e472r4Dr8NDOj8m6uvNHYE9ISMWzkfFnpXQjSMFR3tHfCqMCL+OOM4i
7QZECUcjfPedceRq8kSpTpucJF/b1fLafxjsGWHCk674PKPzyCfIet61dqZ2l7jxzEl1NtTm8TW4
zBFRd24O9ssxWrXkERYb7Z44Ye55ze9LLEc7ENMLDbZuwFkTWc/7Lh3V3UCEdEdpS7HfZGf3TVvb
K9eePvIsVfiPxT5Bh0z3PbaTsaVGA5jTo4OKTnMMky1gWNVdVCUn+ClO/LrymOc2rAq9J55uYq0M
5IoDPEipuEcKDfcQMLs+gA04VE3oIVdGzBSG2H+Rzj27Vb1OUPbjOOTJuuSeG0WsI8Kyrj+xFStZ
snObk525hV2dcXah3EyO4HAckCnYnXaaSHKG6GzQKAtIBnc/nN+NwIDFbROHPLPp5DgCCmUiH7Yo
0DGOGXdjjo2m+63THMjtrkYsifagDrrC4vj6BUCkY8yJ6ejW+DDZkh7Vr6t989/9dPIPzvpktJjm
uR1jNigcty/t42v0SIgc8yDWSJwm4Wvb+d84EJ+wq6JgSIqseC8YHe1xiEbmc3l1DRQlntmcDLg1
Ns/9f/dTECUYTpUvzBJY7sumyR5Ve2BBugHwTzyRh+d+oenomnfecQ1eqC6/BF7A5Sx8h6NULcDu
yLpVnNmAh4e1oM/r09aGG0pOnAhOLRV+8Rmd5POszTOWScU+YcFOqkxlzM/v2KqpTdh8clD9jFfz
ndBad/IVJS1doqF5VCS7lxFNzdTDagwtweA/SEuW1MMU1Ou9jv/nEagxKwPtEqg9olAinfAVPFTc
CrV0ujl0BueJgbJGeP6vw8F8Pd33KQJe561/f1Lbq70Gunf62yHjAe+rnQ0yVgz+ZBvAPqHp7LGW
vGoW0uk5/BQHrtij2+o3++xqMD+/Mjw07vQG/UfdEltza3fqjNKBG7W1U3IIYdlP+b0r9s89/gLC
niL0Iup1RKPPh/6O88D7ezfvyIOL/cwLjhPq+lYfEMEHANbsbHx5Lc4CcdLoNkW09MUmm2ZHpizM
GYd1OfZzsRDIY0j3dMbJZl2F2zn7W3B2kKHIecXoTdcFZp60XFico2vhxyze9ksm/gsLhPPZ4SGY
wAtMUmDj7kOTh8oObfbp8y7R8yoXwWESD8zqz3HaPm0GVuA9BWetWkdZb1RpInPIFk6GsiRO4T66
ssEvWHJv4/9P9v2J7pD3PDukTGVz/Q7g2yhdRV4VpxU9KE1iUc+ImYxNzWuiQHGyP+pb+OTdI69p
xxPah88yiPLNdLikN9GWZYvyvzSL/U/z80/O0HXhuxI/H+Z1TCTEWrImY5Le5zOENaPVMGIWUlZU
D3wFiSP/n/z04tu/dnmLRG2yUAKxckjXKQsPPHAPDK5uzZuFe6jaFyqZ7ghZEeABIDuCC50SEzGR
VeEIL5InCcdncg3rOrbTPd4cFMliE4sqqjZ4GzAVqQa7pJTuwENx8rOOvrXRDaMYNRuTlkMbcaw5
HNnw8vM4QbIcS9iSpbcbZbwB59xy18t6C4eUknTdpuMoerl+xGqSk82aGU8nCunCdxHl2o+wt2jj
JC1i0NCyL7Yr5CGsaIFk0+aujYkQAdMG3clrWSjs8tjn84NO3mgYVeKUfEcV0nMhYPnkKMDH7EoX
Mrcg8AbQchaM9KnHwzfuK6G0wIMnshz2AtbEf66JNPlSUYbK3RjVskLAvdZoPQaR13eYEtPAFgwW
w2g3sK4lpp1q+fGP6hphF7g6DZ+/fg2+J8/zmgviVzXnQ6eWO7ZULR01yv3TBrTkYWcwFkw/hxBO
Swicaw2bakbTh0kFKFTAud3Qj6D9ZFajRo/t6WTuAlGFxxWZ0Ck6Hxa/kGDpdHxRAGNTflaAdv0e
aPq2VLRtUajBlgmF5t/UnYnqKcK7TZLSK2MAYD3iAv0lTMQ61EkPtsJPi3QLCDHTN73r6hFaxTXQ
OhUERfAE+3Fncd5PhVlbsbV9NqG5tgjhWgpdypnk5BpEeetjTh8/rnvdhG/b2fuexkgue/tN4ef3
p2lRrPuzdQYJ0WueN6Vr3PVba2/aJ2PpOKmieejHHAjXplrGYiYc4JlKF8jkX+vatMlIRuUWX05Z
ES/lvQs/lM8MRvpEZyiaE4RqJZ2i9wnaBQCOhw3YE/uPbDZatx6dU+syP2rmll3irVoUiLxwsZHL
NvmzDRLmwrEM5lAxcIt59d463VIFJjER0u6gD95YC2JpC2PRGvYqC6H+dvUlQPaoNg6C6oQESkTj
nMW0jZYtJmJ5x7EAVXGebLIxPBRuRMEunpm9amdIhfaxQn6jBh8VPFIo/3EPrnlhamTblG+jkcpc
FpXqMO3KcmsGq4e5309u1Yegtyv7YF2JrUjStURthCqx9ouTk4ddkRCGIxc9ZSIK14qYD/zR/ut6
DDIGKOHHu0wqLM5brBTlC5MCmW4mxGIP7XZ9mAH7YiL9Frm7OagY2xm2VZmUGoYF1DxBuY2S3OEA
2QtCe7vFRRUSFNyKpl5hwnHigL8xNhA4n810mg6r/2aKX1W8zPWDuv+Ox40ySsuHzUF7zQ8R2k3d
Fl+AbZxyUdEpbWs1ZqeKHiHwBF4wXcZOX7kZGEXT65EXn+JopcrhEZgsuhesb9w2RJzcWBszqtfA
Bkp5pKGgVGoyN5+/JjlHoLPNGMkECyfoywKaUzBmLw0VAmrZ/mebzzOR668NHGhmCbr3U1SSxFPJ
GGq81TBjKGAsKxbBDMIDReMPA/rDK/wFVoQ67unLgxM7gZmiOGy/fkpmgB19zn8mrmjrlL/RuIL4
MqIv/HL8a5JyuDPZiTacikqxlf8j9YM3UYxTTKw6m1QPpuGYsOBSR4+cxqmMDb83HknWxwnoRNqo
DNVprbhZ7QjASeL8PVQ0JzZNWv3iMTAuEuRuyfl/7LuopGJJe/UHDNvV2yVBEXjg5w/68wfrcj35
Y/uMtdQtFR3Q49j1aV28p+heUkeXgbB+v7rZhvJOPCl2ssITyLIebsqM7KpnHCVshaBoCibH6wUE
BFxkO8WJprTZJBpzeMlrmw6ALpG36QGa0U3E3QsLgcZwSbxuS+7RWv9zlgPv99z8hnhd6/V7QGE8
+zYxoRexdhibpcSYofr00eNwRD5tIuI847kmtqCdbA1ELmF1kXdNrH5z1OjP4jbvp/YV3uO6KNuX
93hisSxaPq5vpQZyGIqoWxJo7grL/XaGkAFIO4N9X/s8wGh1NcAn6AJSL9SWKYOQ2PbR7yPs5ZeC
bj8ZyvXg38iUBDEfLcsTT2I6AsmxNePhshS3tALUcuAyUy7iXBE/96sBDqO3vo8VtWVNcD9aAxGk
BA/YLzd1+nh6VxgBCZ3tkzoKZL6ukwj5qwLsgyPrYgEVQLVEWcwRy14ZK2xMJBYbd+trwxMC9fXh
8t58crYPx7HM/rYZFXV5mtKtZAXyKGySq5SpUKOirG8YGrhb/WwqSPWphlLJ+iB43OrKTNFLuHhY
zQ11TypDr56dCCMkBRhH9Uz99p8vgALoFEzpU0VcLBM8FNh9phQmi/aIm/F+byVQhYLGyNf99B0h
dsYQ5b1KYnnWf+oRhgcUQauVvx1MlXCgqydOrvBSvMoWCE3WFlS5YBcNuA0IAO7HHsl6sSn3DCSq
sybIYqPKpDnxjWjKncBCCfv/x1PdKj373NFCzkyxIXRld9pgqe5h5YLq4aImNxCezvvhkkPOmRce
4W5zpWaZKEes2pTHtZMcdyS7gCmxMxwdDUJO9BS5vuisugUu6xJCxqDyq4irg/b9z78ycGoMghr9
RjTISSDHhFhRCLpVh4Gb1s1KpaPtOH9ero2PrwLdtfa4h5mj1s/zlguuzjiEMNj0sAa5dHZWGMBf
4zHBAxmnlebLYiU0fd4JKmra+YKo4PATTQdVWrDlrdB8z5kE0zfcOCNoVTflB7b8Tt76bQZm5/p6
Gz/RXeXONsJuEF+5t3lhEW/buB20GgYhQDec4aLKBaEQVD05b/6YNJOcQiferZAvZwWLymMPOjII
ew9rIzAXoyAsRh33n0O6ASitBV3HIWdvplOkRjG1Dojqwhclc/Ak86hEM5cF1/XRBNsRS3ih/WD6
mN4T+CmEtRUfn0xSjvXWvj/9pRY1mkpbTcKlj2PoTgEsBKvKmZ5nhPx8v7Qfi3oFDvyj7fFlsXPI
h833pEonwHT+ijnykOZCnqOzGCFJyvS+Vn8brzJQavO5K+hhSdSxBuPq3i8knXUip6fPE+SYWFj7
0S0ITMmg3STC9fDXg9OAlz8z/q/BBj+4gk9e33KQ+/fu1Qb788HjNRt9SROYRWRW7PeZPw8GqKSx
zQSVBP1eWTMqoW4MwoB3TeeiHNgfBSsXooOjvEf4USpJEfHd4Imt8aKGk1wWmVhEBuP4LRu4br8d
oG5IfE5F76OmrxH8yTRKRI930XfB35vGYFKPG+BwmH5dX8srjD0z1R0fvaX5BnlCAmQeywXNWp7Z
8/MWNM2EWhCMzfEPN19wcX9WCIflZtHkKQFDV1/tk1cKcxJgAcV5m6RqOjFbzdgB7csKFQoTy5GN
02LP+7/ADs00rTSgDesDQVI+1wSDn8Rsap6vYq37WT3gRpHW5aR1GFrmrAcsfOYDCqRt55/pkpqR
z7pVzWODRG274Y9I7YV0MmxBYX3Tu9BOjGd5xzUfgtmQJJTkROHGxha7r4ELLobrh7nvHRpXhyyb
D7PWLNYvv+Gdze/0QbhO+l5kqgsRoOGk41/WnwYv19sbLQAknF865X99nfN8cAMtn+zSV+gIWhMf
T8p1UfBQnGSn0PvYRR5kX5muvKM+y0mDTQ3RHBytoKD/+Hc6YFlrxlrZDx9bXW74f0aKYcfETRbE
AWgVtwB3oLnicOmh6/48u9vyOXAkKdWlM8hBKqxhGoK9GHMnbQ8QbcgBbyYN9H+S7ZxmGPGmJ9nZ
+I4J/YwqSsXIje7N4zUs3EQsGN3y6fSkZJA+/ACZ7iNOfM9wCbYWG8I4hnoS6D0Bkw5xPJFqU0fD
8wXWM5dbPYh8Xtsu4gehadOCjHZw2rIOQcwujhk5roMsxAXGsWyHG47LLny5ovuWCx0f59a8K9tX
r8ywJeIS6V9f46omdm96487+rMkKSuhnulX5zeYXa9Ck8cI5Wcda5d809IJHwhUo9tPjOjUndvd1
9AO+TxUwnk6DNqs4rOcDBPBE/uN+Wb2WKiC+3YdlTPmvmyEdvR7Mndjm6XziLI7lV78rX8TJaeeg
k/uWkGOnw3J/I4sJe5WVWwj/DDLKG2UFuKM36D96N7j4tWTPWMhuLnlLQ/o7gOtjqw6CHRuhvJnX
UzhWcVosnlc6t5huuHbKnIWzv2apsMb4whPQnORHdAe73zWmG6cNSPbElGXQnyPBrvqlzyiDkKfr
gsUmHmHYNgkb98kOOlLcyp4wp92Wi5N9BQD9RXW4MgxVg8QiY2lx+VMtUGpFWHQEwkYQq8KE68EG
lr0e+Nva4Ni4bhYGOOkeBRLi56stiAtgiD+zT4XEUAFWIcrWAYhK4/1YMid2GHXNeUXBQTVnwcmg
ApntsLqS7VQISHR4MwfdGtDgtygigsItN2aIUfcmCrAsLsOtX+YPaqVJicjXnqQ45X9Jbk7j6O5U
T6X4/ObbCuBniXLTHCxmLt8C4QyGhsMWr0H6CTlnbdOtwr6nXU/GlDdfO1QV8K23aOr5jkF84nWe
kTl5GgvmL/4Uauz7caaXJHPn6gLWS+gGykAzxLpj5pQSipzBN57q4NYg+z9gqssFeeGeGyK2O4nT
sjmhoPf7KqK/UkJ8A8DUuIJrlSCSB7J+5wRU2HXK8GXn0FE6gsFXRVNDBIwxK7cxyOU3MqssCyBq
BdddM2tSZbJ1Sg/DFiFKmvndjaCDFdCGXenDgysCuhvexHHHjEu75HFvLn+j6x0+qtIRxzKRolM8
Vetx65TQRrPJdn68n7iEEEKS8yRU1YBbm8+ZALEko2Wy/0ASgBYVZut+bXg87kMLNaVB4RZv2ZNl
GsXOchz2v3NlnV9HY1I+RW8bV+KTzgyHSpa4ujqIqW9GyitIqjMFM8f1C5a3OB4nO2+GIAOznbiT
5haaU76GVMILEgUvBDXXV76UeYi4HLao4EX7ARYSV74vqGf7ok/qzbakVNpfLj5hCnmD9QX5I2/m
UWkkgnAeuvQNso3+XIT6rBNS/T/KboJdq4r6b9nI9OnbfqYDU/oQjGqfLcWaZOIgtgM4u1CoDFKd
wRKa1l3Bs5QaXreRCLGmxOF2jII69UXxUFu6D0RDTJZHLwT1PerWV6ONJYZfsSjoLuudb94YtN0l
uZ1XXoR37y42L1Y4cjcfmL2lpxvuAwlO1Ryc1e0WrJNfxk5EJVJtbsaSeAUqMCvTFxbbtuca5s9+
n8JpCFeGalKOw2U5MhwrTdE2UIgIsIvHVPR5vBkQmUTePCGPM+GU9PCaXBqlwgm4EPuOU2nHGxc6
0gb2oBPSBOZKeKfcswGN0EySjBEGiNCAUrLTDYZ5KDR2Prbj9Y57Us2ZaHSm28RdcgpoDLSbFerk
9yGgKml6tCazbWazsAH/Q2hBehOiARllAFHm4P79ohpbO9/5+qvak5b0CIRSgNGNYxE/H7FTyMWu
EFmwLV4j3vaArD3efT8qxGv+Ya7YU0T8wugaPeoPyn3OPeSasSP+JL8DVkFo3Km6jyGhMiiHrgsc
9Jf9CbiyumOM8OE2RUC5huOl2F7OplFoCkJks2ISEKXKQjGbZ4kVrtqX6z2OKMoic4vNm61DiWCL
t0EvIsVihhzQJbO2Iy9TqVNgcM2UvwYHDGJ9I3nM+2NWQutENGIWZlqR3WywVoEZPLhuWg3mMpXC
wlxH8KxkIpbMAtXz6HHDTgcyChbe67ExW+b5NaxUV53qhmOJbzxxxQ4xkkn95EHfIaP8pU+23EBn
EFa+cLDSPpxz8sE/KcwcO1C2kXL2yOTXrIcXTkaG8IPmvQQvH5HSulL0pETkkp4ec2ujMmVv7BGG
hGBuchhhDLSeWs1u0uWFkx4z+oy9BCN/RYbJiXV4ouWKwDx9Lu4+NDaaJFPvuBWmvUB0VHAg5Vy4
2nyjG2keZIT5k4+5bu6JTr9zA3T76ivNH+O3SQ9Vqw6DDr1CVObkLv4gDSy71qVpIkCL0/Ap4an+
vIpy8K3Ot//w5qJEf9LkRoCPgoar5gW+rD6NHkA9YgXBnLMYAECHabBTvyc2dcaHFKfv3YLg8Ao7
k4QZT0DXnaiN1bKIeKBy5q/yjnLXcH7H8XaDT81YXX28hQlN/f9PEzTm9QVkMWLrCGnCc8MAG8At
xmuwKCMUFdffJ2kU9upujJmd5HVW//Qsf4RYqvgjbjJrsf2lMcJRLitG3DKPU+VBx/c0njDUVmTX
gVJJOCS1MNMWX/t26JdsOqbR378Fe/D4FfsgEA9w3zeU8tp/dmV06dyvwv/zovWE0GRnEw7+Ou54
SUNDZHBr4WryxRUb1Q/tIY6LI1gukpY6d0RsWQLImWKhlfCKPF9S2IMdXWu+1ErEm/O6frfJn1uC
Gnw6yAtvPOhbPyREGVX5jacyzjQWvqOHb/SqAIL5eEPw0C/1U50SnECK0i8zyobhzfmmozeovIXV
rmz0mjBvMjtxgRihF6+BzgU60se+pH+1nYPfZAKD2QBfFOqyGH5Klt2qSLUXEULPuesQsHivFOfE
cvQiQOKkui2VZecEJbkf26bge5cHlx04b7e7c/Zn18VpI4lNL5v6bYrQxkptSTewphssPyexOU92
5D2dOV8zvo4i5rD2RtWuR3tCOwoyCo/h1FJWpOLHI1LUZa5ATPt2AJgmiugmH4pEVHRpBRaWRQmI
GddeAg+XMLvR4PEHk99PAiMRz7yP32y+RDn/OwHIGer6uMGf9q+tG67KN5/kFqlVQ23jEPfDMTMs
M3ln0eUfvwduGVNmRqNO+Ca0elDuDgCbt3FCseDV88Z6YOj9N/sqiCXnsS0ZuWn69bfueVrktetb
77exfoZGAGp+Rzl67i8jVriVss9Xg8bO2gvgdFjgOniAXu7tRyTfqYG26OvRe3JqG5Vn9Y6D4p/q
6KbXyZ6quVLsnNDTEPUU0hiKRZ63c3tydtgc/wS14FlYZ6b+EZ5aNPeqdLNneYIB9v2vastkV6g8
OOI/oRXbumirwYkdmpf1ZdtyNbnuyVivy+1aM6MZKtb/c8ym/hoxPwK0JLZcYh6z0w1ovPD1dhqe
xClXMvxUVIMwukcFXOoayWpDbAmLjyvYmAY22sHO9g1nFdxmfoOejz97pza++JUfyVfcmFPb7SF5
fyOS88RnX0TMUTKFwAI8vGmP2HU8qeIU94a4B0nKL50OSRZdsFgKxgdHmZjbtHDBDOAiON/FSsRZ
O44H31tMUZwyK1Us3Z441czcAer+4fDAgy8B8dRcjmDxT027zbgYGbGX4kgNpv0hq7zAvqmE2hLP
qOU2YeidEAy+A4nQDdJdBDVUNDiQL2Y9L9XAaGdpcVbdz5s7OIlCbZthMBeTrNysrtOgQBsveTcJ
kEDeTRAhp/ud6q5jfCCSNYLAW67Jdgy1tbMNEk3woA7nq2Odbm9bbak28aLGb4Z/xIP3k3MplgwV
lg15IeehdYHPPY/koXivww1lsA8/91bYXPUS2x64hUky0aJpUiZdH6F+LFjzP2bLHOLvDiVYO9hC
mYWSOHxLC4zjkFSHkqzEq6jG8GsoCJ9KNyRsmQd2K9Mo55kl26rMAAnVTlN5bdhhTG9hf5SBcknt
oslmoPbeoOnclahsss5cvU4avqwCK6EX0NtYS4LxpRtV6mKlO0OLrWm5BiBsjst7TtoTTyHGAVq+
k3B5JCEUQovKLAMagU+49brs2rID/3vieWpouyA3VAz5bTouuL0XQ3uKIHIgkQUiOzJhxIH2yoGA
VZVm82BFw3nhfB0086UrKtc/p1uvMDcZ+vNQ3bw2Ksl/DmK8hqZG8YwjNOy3yGJRWyiBlR7zX1CT
HAPVrzesolk9dXI3RZ6hTBKeoX1/8fuj+5ozNhuF3BXo4Hlss0AejHT1tcnrNO8HgBErFocVFTZH
kb5ta5Py/bnUGjJItJ/GXKcEfXGwUPf0nnfcPZjwS5QfGlpBM1NdJoFeUpNyezFIpUw4TyhBzxUT
NipN7tjICnJTBSxj2wr05EHjkiNCR2xH7xJezmHnCo9PuVvsjWfRBHj6HSVjNidle8RrlKmna9f7
Byqe7UC5hoKQKsr5xZ4sDTHc4jSvOIVS45btFk7JWd9p5U1rqppyKBfKCzlC1jHQvzk1Lpd7oQci
y5u+xYPijkBDvbfre+OHtYLZ920EQiArK2ct3vRZXxPdbTuE3Ck4JQ6x5k29l4cUwS3cZLw1FTCq
7VUq/A6iE/YyNb0lgWiuIzOFxQCoZqimQ3F8dz8/La8NMV1IsqQ+Q0AxS6eBehegvHEBPqYzWUmm
35oWPLk2H5WCPPSpWa8CHvpMN7c/B7nbgB5U2zuNqkbaUeDW5z+/BjkKAcLfsQf5gEJrGZPuv+Vs
vx14dk+HThDqTzy8LzznhNeujjZ36OgrizdBWrJ92oQ/T3uwHjkAWpyTmyAOlyDz4+1cwGH9Ulcr
P+fO+Q0k0TTKRDppCjqUMm8jByYhqqkxZ9y5EgVMeG5Hbjf2NBBUVf39DF9Jn5fxfenrQdezIE4W
dOWFMIpEQZAma5/+NpqvNJKSUdrF916lS9uu9oItQQv1LsqaSAnDEXCERBMDMqjdnFL0Tv0vPVjE
33Ppd95QqRBOPoQyJW3Ndk8oKKMl4VLi1oP/VkY/p1Vd2EuXalQFMInxPLBKDrvD5xE/V7gauOBc
zVm4IfN9yxWsJtUuwgRI6LnAE0d5vHDNF8g78btFAxmRXsv5zHiE20HE0ogSLkAa+m0UQaYVaMeE
aASESw60Vhrdv3QIE4SHY6aH5/M+a4OWBEVgGZl1/ZNqwRP8ZqE3cWtzRRuu0n8PROSCJzKoFq9q
Upjj4YKSXnreoNGDI7PSCjJIUPQT8915DqgwzJb1uz2U5Rvp7ZESXjGFliMT/rJbb+36wOGPhfud
+k2ih6DZjbNdPSdqjXMxoHla/jnPSNvikOg7vw8b4gYcYLZ0WbdKFOjXHBOdhwIEQBvYgb5DVsBL
boGSdhsitMoaP2rrUiiqD7EwS6uBGVkWwMhiVUUy097MmcMQMq/M2Cso771im8j3SOgEYheX6mQg
aPVpfDqfOgLtj3vGym8rPTkD1QQ1HatUNbmw66lJMUEDz6NrBUxDalZtZmfkD3oDU8kuGnBAiAJX
BJYk5XAPoI+jepFy9VpyKP7njyylE56gsnBpyKtpm0diCpLGevZGUWhJg3r0jE3kv2i52jAcRMVB
AUswUjaJEcjuXx6187ywlIs9+T2IXLCm0evPWEIAwLHcbiMDn0LqWdZ5TqxMH0W6doOJZPG+8wxf
p7Ljt0caMmM36DHt4qg0PHRajWRweRrz+SAdLm8wZjvPLozy0/T25kcYsL8M79vbhmXAoMfIPTcr
pKgh5FHBprCpfJ4VBHM13xOglpKpB905zCl9GpQJzABd1tIDbmzVDX1feXq+aE8x51F7CtFXScXJ
7TA/16OVdwWIkB2/RztulddgudOObiROnVUjfjJMVFfYoVW9bdMju34cbUiYOsHoUF0Kre1FJtfh
IgBpKTe3LrjcmznKIml/jNnfu18P0Z6u6W0cLdgjjx+CQpUZng9i6dFNpysMDlSU5iFVsHM09M52
YvCuQvLk4jGekqEvN5n5mzDGHMxUGrG8WP6yNXs82xfGuT7A2w6PQXOn/Gc2WRpX6cOsqNuqCW/S
6iQW2A40wojMweEDukMoL/O+yqLf4qfixXUfSapX13I4jPr9yHAgu/ZSfrMzqNXdI4QkzDc7wqa4
sE7kMhanb2J+7zUqYsZQyLlOd6AaXy/cXfjEdubWwxvJt9cHhE7QdUYLcIIOT1iE+ugWXFg/pk9P
b9+x340iUREfnhVxE9gpHbND4hxBaWDWN2/7Xwf4ATq9C5kYhLSOK9eUmnG4MA6lT5YmhDShQWu6
eBrwTeV8PZl6Kfc11Xy+MwnfVHORy9Wauj3Yj+/kOheAWmZ33VojIIoPct7SSS044PMI/L9iZWHu
kL7zlpd3FKllkVMFnzylCyQzyd1delHRrtW400+Guzopzhny8BTTWAqIkAPpA+e9I6Nwd+D+ZrcF
D8/ZBpQea3ppHdrzuWu7tA7aLSKf6sh1BsiujsoISsBV2e1KmEPD3fvH3pvYc+jkpH6KBLzS6WFE
jKFpy6zEtMTGaUhDM8IpEaAuJ1JzccvORAuau5NZbYtC57L9cm4Ecgqg/l0MDGeAF1oBXr//y8qC
3iDdQJL2ropSOFAz59RwJioxR95DtkuWXEebPalVsrfcXrCE+P40TZR62IKZh42rxeinL48meQ2p
GfH5S7vRggVEKjBLagfk8buRmupt6TCb4Opr1uK2WuvWbjliplZV+OeImAk+sxNOBLGb+3vfd1l4
vSitm5NXLL9aDc1kW0JJ1IqC+R7o0XHbMX2lgNKGsq7TCYCXqFcHDk18Vld64h126z9Zd8FB1+Yl
YjyNL1REfZRL+sihssLohpBh/xdo/54pYqh2SqFNp/4ADEWeBdzNVDLLfmeo/5rwVIU4SmiM+6Uu
OT+88QpOLAsghbCSu6Oca5cXlAlNlhWEum+lqqwArCsp5uDm+tU+pYIDrX9Iyy5FvAuf0vHvdccB
ZjYq7ZkpUngBH/dIrs//cKzBS9nxE8B2PgKU+d2Squ9+D3jZpkfyQA1nSrEb5ze5dGmZLKBP/ZLy
rqzOSrUKxtlNt64OaFBx5QD2FtW8odTDQv4GAsJihbzrB9X57KL7R6xznAbvsP6CJHSsputolS1Z
bo83f2EnIaXEkO0s5mxM/JEwSAklO7EIXudCFSNvuzkdIV36AUypQS+X8/NC9t5MrfRs5IRMrsOt
feXlw86DaxnwWfBvoLnIbtKK2dZElqi2sML9A1AHHjJoSfmcWs6MUiqzg+oMelfKnjTWFNthfpNQ
Zgy5cAiw/m7gPQYpdrtgUUZeDSkse2ydygsANZOgybXhKLGDafrLA4n5SIFVmk6yv8qYDi06BGlH
idjqQmRskiHaIirqvvQJuz8lz7KYgKR3W/X+FmCzm7fJLbSDbxeDJEEdrHHPZABzj6QP9MycLh8P
GPD5kIvIbSO6/9B5qTIhilL0QBxZPa41NGOvrB4G0NbbJWRKc1AOjW4qXedmfrONBuMLnk51qOY9
jGR8Bj4hmHFXCotXUxNJ5Jia0XG2N4nYO/85/lwvbK2h3MNGMCYNnATupqkmUbqLWqZc+tGwpVhh
0SYGaePbrA9qAXTaX7Lck4M6xHzNDPDjLylXy96O2vw50vEPk7VQdzDyjD68yXcIbofIWr7UR4oF
ZZJLuOqL0Qf9nAdkjBGOl7+vCV9lDYkgqyGZYhSMj4KXQ1enf+NyvsCuVeoitCUNR6lZEtg5L7b+
ZbpfNO0Gdu+vashv6rY8rZ6Oepp0u4gc7JNoKLd1/qkaahwVlaRx0vg8/OgWuVTWk/qK3J1pJUKH
NbI8u61h/P4iHt55uN3WuvYTOF7smGlGB4p/yCUyetZaITGRPWViFJrOTuq6yzTILne724u97Vcs
/s/H+8euKsUGJlEedyaXgbZ74KcaHpuMmtmxYwMXQA75gxv9XuOwu06SYawizjS6GM9tOxzjlhvY
01UFwUcbDlmfXuLFbnRKuJLfGeU0B4TjbfSZyIwxNhoiJVPAzHS3Atg1wHPCOBUK7h0VwxMl+dmr
klqb/YNVOLnZqo4BFoIkVbtFAbZh01F2BlRxML2PlTgoJeZlhZ3qppQ+2spSbIMPIzq9j29VEPu2
DZWTFVp2SqBHBpaqVPs1quOZZQGQkxcUA9xRbmjuH6tn6iKygIPmUr1H09R38HsgTKq7wa/nT/R9
0WVZ8N61Uz9N6QqHEyaV1ShF0RHP4QRx7GfJDdRHxXFYt2Bm9DZPQePJpauIAi35H/gvbgosq3D8
V2hWK8VC80JCVjlg9M5QXbKEHswR/1nR5zJRHhRRN39Q+BA+L1M0IU1wK9mAhjBeEvFfbqapRVhS
kcTbz4gOKI9ZfrgoDsAtLvK8uEc7kbpSzZ/qm8gbXL8J/UB+8+XLfc9tVlAQD18VGXlVEg5We9N+
nnLPkTFARgjbwNhtFMlKMYDOU6OKmNoNIhm1QYfpHuAEun6/+SnfUbDkjgVbQyzX966ABTD/EKGj
fYGXMdNKPJQnt/dZOFMC5l/QA3deHh7ZCUVU02RMOwdw/45eUEoE/6jhO5+tWfvQxLgz6ew/l2PE
9kwlNMDDI5mu80ihIfn2HHbWE4ZrU6TQ06+XdhatIfMxZDyJqo2UuwGSRRBK6bNVnSaHPCgBTLZl
uXIMJ4jrrio59Bsn/bTjB2NuBVHXqWXSBdHcL5vgJf+4K2RXbCEaM99bXJIm1Vk41Iv2hnKnzKNU
FPQkoptoF8UdeJA7WHb8Nqii6bbm1lZiC301qfKCCvgP/3gG1SCaCMXSc+KXNVKhYX17tSQRTJDH
iGZc26U/SIxMW8Nm8hdL5W+0mQC7PApP3iU+N/yFEcSzayQedpxpItnZx3vrv7p3Xplp5L4iP5aN
2I0JGKT94Ok6vFUe/lnkPIsuTciaKFK2AHjt4RseEKIPrFcCJHrGnEVtIs/SbCgZY5gfTg7bQtUB
H+DKMZRuPu2MNbldr98/Fwpl9P/cLNR4GqTy/iZWvzFVSI0ysBaPzmXon9jdtr1j3vzahpr+XJxe
J6eW8Vm8Vl2frxTfM0eXj6OShcz0+U5aIbkvHIy35E2JNv6pCEshxIfqqowDQset8NcED6inKe3U
vnSjCjEHgkWpzK26QFjZxG+aEtDBCJV3IATchRk3z+STIOiSUZrivMcMnZ3UnJ/psQ9NKVkj287C
JaFIjEK+dTEaJ+QLoGUmZ0A2RA22znfz+hvNrD4VMozpKCt+FwrPOtY7ssUtL0useDGz0+TEh3wg
YESLYQPjdbmlLPpYiJZHaTPlxfYEHZaiWg8peS5U7lD022xCc8zPMqmfHl0fQ6E7oFQyhEe0vr7c
bnd21EtSMkR1cKazGhtgzV6Zcr1pP6SbZJ+TRWJCYS+b7pMGBKnShJ9PSTqSat451vYBxIOHS5l2
lkowL413YSDpr3OtyTWz01XxSRFNpAdZ2rTpuFltavqvTEk7aPstGKPcoeT1k1qInwTAjGQZBFhL
exxrZyqsXyfPqIS16tMscQrBI6AAIK8DQNnxRGHIDExTouyRSVa7T82H/Vqw1AJA6BaIYRoby0gf
fR3BLUZpm9W4Ux4N+ambxXydPtOKgcVvhgFjZYxz7Y6rOSIjAM9HT9KTDsr+1g6kZN8lbdAKB9zf
o3Hpv6iAJY3iLn3KXvVK3fWePt8LnfbCtwejtLXMfCDGl5jXjmbPIngQyl3JWxiSJOt3Q4Ij1X5h
xtTubMo0a7EFlgH+5DwgS1tc7AIdzOhOerA8L8uJ9HLfLhboJOp+5MRYOIsrOmcrB53huEQWsgNb
ZdZ+USEad12IA0WVUSE9P/cw6OuUC8UuY1lZ8dHzk2JaqtGBoUgxynCcnRF68qA2DWi1M3rNFGt+
d0b7yhaO3mPeJpBbGEBNkO/ziu2bG5i2QqOvM+U9i4zQh6bfC1VITPj4fKagPGWYfJ7ng8a/p4Zj
O8bW8WDpNbWfbpVg8abTSakB6s+RcogURGOvDg/It1EbUj4C6CFS2cCziYt2Bo6Ct7FqKpv1KDNa
uReDhjfuVuaywDshYggJk5irSIh9UIq1/D6c3zClGOsZziDAqExqhHlKYDcZomAB9GZ2u17BOCwG
R2zr+akCyYcC088kyENDc6nXg5Y7z0s5Ao2XHyzSqQdnVbNw/WO1cSgQnLsane0tJE5l9xIAaB39
M40cYjAKI9s+iimPwBMQQXJ8WICLjxl4MSbG5Pm6Kn//vwnqw2qVGs4Z9j+9DWdVDZqjlNFJLPer
n+6Yww0JXcKtQCP3izPXL97p2C3xJRXEVl8Gju9MxnRkgaF/W2/YWsy1bQAerO81jhgiMEH3O4rE
6GwdRvSz1Yu6XdUWyLe9W9VP/6mcnkwMdZCm2PolewL5LHaR8Lk4+F3k6vzakzjnVD2WaFTulICt
zerJxk4oScqCi6LC1wf4L6taObM2wLbfVymwyJ82YlUN5W55oYCGARijQKvJCNRNJCIUVf1BsjKM
yRmXHIp3QUwSyDurJTaiQwlCWqK7lZ85Xq0CaCFrIi3dp4P+TxGx1OWksV5ewxeOPlaZVOGpsS71
bZRvylp57nrEIlCOoqd0IpRE7bmVck/8TjEdSNsVkGUQU2dhh04gio+jgervKOYPJL9TWpqM5/Zv
0yqU9xMZDPuUhhRe4gOounspkaFx8UOB4lEbkc3X8oeMyIguyZhWnE6X1gJvZsXZSZZ2vfw4bvWS
rcIsU5QCo1mmhFGuJ8Jcueongq2GDxOT03yr2Uzn0lWf/bF14KNsHKnK4pmhtwhI2RoSPiO2Rejl
p9fGm1EONmCbwbzuf0lObDsgVpLSCek0ovwOnRb6pSepcpMbIHRMhqQcYVez0WefJs1x+nfqYoVk
dMOLcjmNsWC09ggMzeMYbVBCj68AFJD3sS6/n9sQ7XkDzmcRhTrc9n9vWuQ1b+vB2m+bVfh4OsjV
oUZ0nlEWcv92oQfqYmHj1vBa9DLVO9i1U+eXx5KUbz0n8sxDnrRc0lqOAiiwekXLw09wrd4ugD5J
przpqug+8/g6855HMf1Blu1h7qbRWWUGbCgVnI+QtNc6JHqEF90rsJYn0dsk+ggThkYi++CySjbW
jduA0XxPYtcgU8vI5MAJv0GsZAEVa528JVwwRo4x4/tKoZ62L/fWugv/pwCP+e7fOawVl6kmexbN
Grww+bzrk6BE1Z+7Rk08RUH4ZtDen/Ci695ygOvcVgsR51rI4zzcck91invtFbRc0ialng9fCdEa
biT4oy0/SRY6pSRG9QMrsSs5LGC4I6DQjCEWIS74pEPxAhmhDtXMlnR9T7Hi/pCV0b8KBjJS4a8V
7kig01PDwhOWaJ1S8brCAj9e/25sc6hnzxjhxXEnsgCqpIury1tPZlzIGRmaJINrWPwaWbmPBJMF
tE/tY+eM8czHsx7OJlvz6NXvxc02MWhqqALwnNGZEPkG/1P9zucYcqS2SUleukc9sy+zWOvxzYY4
GvGRL4Q9V22Biw5xNxBWJqel73ZOZchip55QVbnU4xy5Eus7WLtGPmOIKbnZCizksipqm5nNpj94
vM0iq2fTd03idFtJroFUzvK066wPHIeCBZBRTtqCLh+qvh5olsjC0zIED0LYeTL37v1j0Oj4xZaZ
2zASLpluxwXpCrU7LFDStFxfXvp35i7bY5Z1dKqA0Jmg/SORaOq3+W6PKig+lDiPZ5ms6deYUCpK
kzowB62+2JqgHl4rLYmVGOjOXctYYnmCth1KATklX7W233GDvX1PJRHK7l2F4RAxgk77G0H9Cs+f
Ba+D/zbwTvQpnX8HrZou9HpIrlL8Ns0eCMzpespu8YlewxXgco0+dsoR6lThIUSSnhAaASEiVC1r
NOKHzTB3socf9UHCr6RUAJL9QcGXR5ocbJ+PBVQhOGhBVxbBoP5tm6Icbqxv7fmvpvqd2D5WiFvL
Qzejk//XNjMjxHXT4DIrHZbh8OJ3FTbuk/kFIPKooLvyr6fmTalz7POb9pDesurH/t3I3v9PWwqp
YiQpHZiLzZo0fRlWSc2j/8mijiknhPDF0VQ0wbTb/u+jnN5E7Khht3ZMoGBy+H5xK803haJpoMMJ
Qp9748F4dj5Phq7fGI44ShD1CMICb/uBMAsXz1GWxp3HNd7oUR6vzSvat6Gu0V/7F+sbfFHEp5Ai
6UfT54wTioZq9rg8COA4fpqrnpH/Bhz99YwsNfY4XDpOQlV5NMsvX5oUNHDvs1MHFsN5UflGOtNm
G+VGHMnSBjdWWrOtAlW/PK5u3uxhJggtOD2ZBsUFKprBxQiBZmUqIJrvSr0z2VtamutfsVViou5P
51/vBXN69I7fYT2s3rSx4ed5ydVd06LjmMqaPUT0BpYSzZ+EGZoivN0tcyhLwJSJry+alWf209YL
8DEXwPruBdzSLV3/1nV8mNzNgO6J//g0RchPwjwGSgTWx3xGTFCcS4b+R640CCWr1P4Vf2EZxa1l
uSzS/YJk8LUBzP1JQPq8bV3pYjUI739QyP0KZbPqeXfQcLHmvr0GUyMS7fguQtR4vKwusRNOpXwl
JgF6wA2FDBOQWkNuSXO5MmaH2l8UfUy7pLlAvA56uTuiO2Hn9sGcaeUalu8j+6/pHuHZ9SqsvibW
109ZnbTAXaoLepeFsGvRi8lUs6eAmlhmagIo9dUVemZ0usdo+3BVegsswaVNRQf7NyVEyxPxzc+Q
fRDjUxVkUg0zmJSyMaoYeiK0DwoJTpy5J8g+FeOgJLDD9ydCMPqxteALHXzyEk/iQoRBMlpzmQFB
FB4iPZKh4kjQzZqZf0t2J4eyCMS+mNiugfYnzhZUeYEbomv3+uuL/BU7oiLHL032urouk9CYf6UX
AJxUeKUd9aayFOA/og24PU9sbtpT9gsr5l4x2edLLEDTvPYa6clsr7EDdTHNf+cTOLqF4V6/h1nU
YWCKHpm27BPVeYOtkOrQn4kbjls32JwqqNfSQD0+lPZ06tl3IWu77r8eqnpClbmxgfKP2XpGWGm0
g0qnInl3bJ3YQ4fBfyjjCaORzPYLV8COz8/L0TwD0DK7mYaJpjiLKGADKYPYVZ1+ww0r6R5Jmkhp
4LfMPTlOuF66KQxOdqLMa1kU1/6RY0GF/FVTXmQfFPrX3frUsStRvHJumk8jhIcimAOxwU5+0Btf
XVAxnSASRdVN+MPwgy3MaeTtfqK/eOpmwI7QDm7sAIz6fNF22ecqxTXCnzbfT53DUJQN+JenZbvs
ONNQe27cAPK1fZuJyDaQfS8zTm9Ckp1Dj81DuiAPuBAj/PwLDXzqg4L3HmDk+P0Um1Bu0m6sOJex
WGlOPAMDbwgUoCfug+p9OXZ6DRN+eX+/P3pfsq1WNDQX7aUyOVx4Eas4b9kmaRQOUniwJQko2GRn
4JCQZo7De/A4yLrC+0drTXSs3UrWkmIKdOR/vbZ0f3cRN6IoG3mdArk53mP2qO/EVwgfTqEMGq+7
jAAefjxkS1IcRdpUVBCJ0znwaGBqLJalNTcLGaCj5YWYpmkniSE95T1PN8H1Hw7kb/7GHPUuQpNE
jjnvvrq9KruaY2JlC9SuvD7CseXa2Ltmn8DKtNlLMV1g4zVNVQwUU0Z+O5TLhS4mA2CYOhnXEzhk
h/7VIoJxk5WJa0fKAnI+m9Ns9qBehzmKmwZRb9jqojGmugxd/91HDz0pAonG+63aGO/Scr8F7mnp
+gbB6LdwRf7964HIaNXnaGUNPDozSq14qSbZQhPthgEbkKz3XKpfxseprGwEp1hOCU3gQ7tBX4lV
Z9RjuAUGCiTgwlavw90piapExGzjfIJnTY9orqAPox4uTerAG39AjhRJGaaQWVlmagvEYGl/K93y
ogK2+bYLH4AD2mIdEAIAIH+UrYOxqHNCj2Qok8xK54FeXdaNbFymuzmlpdX1S7cq/AY8CFaP/AM+
ZJq0gTeC5f2prHRGjKOWPdKL2dt/Xn6vO5ByMekyXtwT+CzFpobiYX8WmlBI4yhQ2ANF2QkKTLts
xcN3nPQo16HV3GidNbQbWcFm0K8iejujAFUr2V6vuEgvV4phFypzw6D1jAlWbB+vYKehlb2Kbhvg
7GwnJJM7SvAfYklSFOI2Kqn74RYadmt8uwzUeb7Bx9bLfTJniEn52vbOz/cqHfORwx5tMj78P+Bw
Sy3Z6wflkKGRJ6LWNFRMcjJM2Yu4tjZZdmFn0NavEB6UvPU+EzIMUYzkdaagkOb5Vg89/L5XuSys
Arq913zPOzScJnVTCFBPVevhxYJlu7Gl2QDxwjbvzUDfdOK/GsajWL/dizn8QVh0B3rJzFcMnV+c
nyz57afWT+kcBxMnEz23ePioNBOXWTtte4vYRNR8Hrzh8GW8SEGumglHgLgT9hvx1u5HXCN0ZFch
q6pxF7Ao053s2CV4fOcHCKATsapJiByoUojs+U6yYZWMXd9QWYV1KzIlKVJJVpuHS1HCFEVeX0fs
tsU3xFdNO+LB9Gjf48qpy3VW4vJu4zmqUvqkGBm30OU4WAx2cpv0a7K81MZMXpPUUFJ+zelz16ja
YdRx+82BGU4LpMZAwxEBKDgFZg2xl/MVzqHgb04HWUGHK5SJUcdaN2W4pe+lEDgoOA/3OAdxRLHY
CSF4k51KUdJYgE/LFC3UH789+gw0lwiDvaIng1NwUPu5qrHoG0LwB4AEJTsFgjBOIQmxzsxgXLtH
rO5Y9WNggC9gYRj6SVZri6hLEf73rbFTn7G7HDK/7UmxKDdcrFNspB9MATcT7np58GuuQHDNhYEW
Gn9LQb09j7DWJ1tU2IcMri4NMXyzG5k8DM00b3KtdFGW0mTxmkBbRGP8xCyI3h/sthCiv1q6cUao
LMAtb8HpC+EmGDdVGfH3M3b9GnTTmo03uiJbl1oi+UPLu5dcpZmpOMTDymORhIReElMNe9E/Mp+Q
U08ML/FdsUeMtLM2Yxiqcb3m1bJE/7Pw1Olo0rb9dQFVbK6/V8292OqVLh0ordi4AMMtqDFd/vSW
bYfLsi92Tm0Bx2GoImoNF/5TZvuCzphNICnbqTeYZVu6N2C2mRqmudCUfd+9XGNARKxHkJptbCNO
rcdsdXCA87COUR9HOQ2xchRExpwMhLJ2Xeb9Z8BXQDQ0KWuZgnlsfQUXcx6a8r5VdVU0OoBJCm/I
7mtIYsyy12GnTdwD2Bkuu4xglEaK9V5HiEy/rXZwrZK5sYwZpY+KNdNRyYuTxV+tldkmbq+vpV2B
0Fe4BemSelQZVSZFEAvmtI169o1Gfw91e/xsLvLEC48TJVzFCG1tdRdCq9frR6OkktS9oo1ZdDP2
RhWH+szSNFcRqO/VI1C978k77zaYn8ypd0Qf4aF0J1j7XwgEM8Y+BHgk7dFpKpSin/sral0JHEJ8
nTarfrG05Jr5aVeLByxz9I2lw1ZgSPJXEJitFOPpooQ+dcEeUbMkn8p7Wz1djnFaq62VZVqkmz+H
RdmTxHH0+/yIbFP01jyJByLAIPFVitSR90CfeeDuSKXPnbY6zbNrShhX3ny9hMRXnwlwZ7EI7KuK
eo/I5HREoPCFYu3u8nRdCusV1RQDXBLg1QWLXJafLxncr/1uTy83gEnXk4RI2Wx8xB2DwRzMKtKV
+BAFA5VtyVwIVoODPU6qNLpGMWhosfKD169Epp0Ln0JKG+5CQdc8wLONn9ngffBdHw+RlEHvbK7e
pIzefHIZx8RBieovhYgy5jZZmj9L2X36MG0fQX9cDRbpYTRcQJSkuvQDI4dXWf6ccrvAXHIPJXh4
R8DwcrsmmI7UXJizj36zd7mDIVNngsSFUBHat+466JLYGIx6xxD+ucUnDFlQX//Au0tBoLGFzZ72
UbNGeHnn7Pf1+y/Rxc38T5pFM1WEMYPzdgQUvuoQNCqdvjmywhlL8Lt/r0+qwE2W8rIvshmdJSCi
/ZyMvzxut38WNzxcVZ0f30qkGtjYRQD4cShMgkgY4cfvfjpCGe9g8WZsu5og76Okw7dy9GGdiWUE
4JWhWElsDfIDZpoa0tbQzeNerEnVUuT0OncJwlY8aKjWE34dsGlXgLEx0txch0DfodtfoPG4A53P
IEN4eL+awsJVsDJRjyfuiGNd0AKzpoRRqoh1HRtzggNnm50gRoOsWGqPZa6g81nVGZiM1kqZvYrv
5pL6S2Cs4gOIIRbgonOfBLaCqDb+BQ3jjR13NiGBA4Rpp1JWDfMu9uN/d9ixQYdOOAPGGd0/afaF
IipCAjSWUizWwEmmortClF4C14nMd6zyK6DWPAB5WV2OJWGGkuzDnpERyUhwUkWmQ02EkHn787Yy
84zDILp01UDZ+OPxE9EggpvytfFACABbjodxaSvSCFJJi+XqQEN2QPdQxcGvEhkhldFgNSxO/zdr
n3gEw76O/dEW3ZNOob7KND8zpEtBDeUP4vDjersQnmULow0zIPevrExJlXYziQ/xWwbGgC2dH1o0
aBqlb/LJHdDtkDGx6D4Z1bm9ymWYUoTFdmOnKdlb1sAfo2dP2zWuFZyaiqR6aX9g/lMvCnKM6PlG
ULWqHFmbSV0pLBYEvqynfMYGTny8LXfLpz9/0uQWYu5XRnnTNGRHZaQuVYdKEPIF9pHxAVvfugfj
7KS+YgInA5lkZzzFmG3UZpvnivHVUen59t0bESlluwY9z6JWdwUuOB3DdLjZ9ILh4sCNh1MV/Iw1
3zWOEBameX5lsOVXyOXqkSmef950o6zg1JXm5NmHoh31DXbEcs/bPwp1PaJX6AoRpyy/Jjq3h+55
mcVSR82qdUWt0Q36GQN41CH4qo26AOteZegS4Pifr/DG9hnhcGo9Kmqp+NTeKMo/DJdJDc+yorz1
V0+gsupi6dGbFMW/PHoeh3jqe9EgKNZCx+C5r8Rgei0RyL/byp2/ozaCMxaB3vv37/Ew1s4Mxdd4
M/k38in8nQOROmKNuNeZpybcE/qXMJuerQjSYqFsGRZZmHAFR+fA+jVDEmSl+pr4Z6J8xJxBZ8Fw
rJGzTQBsfJBKaLj4cnqfl48HqrI41sjrgaxac4x+p53ylT3R1PWbUFF+OWk8qSxExZ5hxo3/VwhA
U+6ILL3zk0OlTOUhGAF1UnIQthfpleOQEVXnlgv7KwIn5cFKoB/gC7rrj1vaweuSAS9QkugdT/Kw
9ePssE5yaqF1byiWAZHqdhD/IfxRLkIv1HfNy8qzsEDKcnkm/2/FgBt9pS+FvGOzHntr2zTwEPls
vrCa97xfTHH1CxwSUGiHwr5qprLrKHSjmumUt4/JjYCNL66upeTDVwKoljJEg2n90V0/pLXO2b9L
mMgYFO4CdQpkgP9kIzKziR4YP4ceXiMnHYEzTZg/gayTziE0aHlhDuyge5Ua8h+FPw55auXL7PcU
Cq68ejBMrxrByHKaRRMLZqyGxBnvTG4EAkly665CJqP4z6Q78DPwO0K2yGyTDio6P9Db1FDk6Zyo
GT9uw0HA1Jh5zak0CKqNDIdCNXxAm/zfWzW4OUQg+j0CJgKyQcfOgTw8K22tBLgDm8uIhLqZwi7q
Nrokbiyxpj9r5aEY1uGCtrxxUBCbm9g61uvuCs5yyZ8hmt/t96KbbA9yJVxBQJj4iYw5WYtCtjuO
aKNxnYnXIQhiCRIPeZGOsqKGPdL3Fbvcv2JmU2QPFpCNnSAQV9fhpMSMQi+3D5sxLQeIvmNwGYE6
lw630BWJKzNApjchblHHEaT1jp2EaorqVuttsRkiZ7s3gzuYL0P0Pud8QsoL170NVbipaXqpbbQ2
bJV5pGvHSyP2Bwz1InLVfic+hyCGdYZd+1BH8Ir37J+P8GukS6Dj8DpmDWLBL6AxT+bY2pSHogI6
gf8EOVmALMCcB0GXtprgzzje2gsWUPV6B1ehM+wHDytmNfI37WsHJFRKShoBKO02VziOTCAH4iXx
lPlRjg1OCzSTjnpBLuYHp3TaKyZot2llcUEnzoNWyED6T/vaD1S8uaWcwzaRw5kmdTp8w8uFeWno
jg4qUJAbz+fjHmr2vY61y+BOW0X4+K5kcGKpEzFGUhMc0aWU3MiYGh4lJxX7YsASyUtbFxkLETcW
5CaU9gVdVhJBsUASxW87ADFWCycbcAYHmwtxfWFo08QniAE9L3JZai+svEBmgaEGRnFnDH0mtCoU
AuzaFRmmeXNukrwDeo12Cs2eGnqXO3w+WDu6OrFHbO/PYCsK5wyPdlx+wy50XarE3zCDnG+tPmSi
GK/aw7ZS/Fz9o11Z0Fv1mH/6kIiTX9/o28K1UERbpvd0cuaIgYmWpi0TloTueemhy4OvlbJtZTAR
HOAoURzFUQyiFw4gdP9iVG0y6B34eVWRGu68DH29J2+q+gd1tfdo7Q7tJ7iSZ/RgiLRYpFhcvhFA
30Ua0oaKg1EJtI/ynQl99V6c8YTRzX4i1gcZiP8ATTafGeOv2JL3MAdsZvvcgXmiDn/Fc3UTam65
KmpyWCDZ7PtirJUAzhpSf1aW5MoXlzUgq87zp9CNJbygOE6z0ZtsLskoFyzFXXK3t4L6IJksQkF5
KDCA+Wt36wBP5W05MJ9WH9UMxHHcjN++gIORXOXaBQns8pj0kNqHB8d+/yARZieryCobdkO7HGNr
l742QnyzE1TQ27jn6uzyGhDkKcb8ss6TtmqV7X8n5J3X4ZR+oKO53nOnQkTvsp9QEtUgskIIotup
anGDgH7oSkiGWCCXGc1sYJrvD21aUjv0wIXpkfhKbeD7xTPCJcwehxxPPv0/nCFlZrv80vlMuXEu
QWx7y+Hj0g33aFp9lJJIrpmo5jLSmsh46Effo7ePzRa5uh9USCXuHhGXzMNdrseUCvzPcUKwRGSD
fRyFvZI7Zst3G274PW4378mUQRFXevtTvlj6Fwf5HyTNhAUgROmhwbv5WmM8+H/3F5WT3TSRFlHb
N7ayIZuffwUcW73AX9S3GPIBInsIpJXj6yXAto5upLBcUdxdYHSr/GIq1gAeTeW9/rZpuuTX4lMi
2onEaOT595YfV/DEueHBczWwqIK9h7sU/gGMoz3+57M83ihb3xV+VhyHLKxkN0NZYZBsYPLv1uft
fCHa74OZucA4bKnB6yAxo5746H5/jlYH8eECvSt3o71bG9j9VNs84pN4QFFA3lMxgEE0ABJrLdaH
x7jaQ6cT5OIpxrVg4huMaw1gOkWpLQc5vBqEK2++VSFUjVr4KQ1WzB/1DsVKjOTQ6LONdkkGMMWo
Kn4iDoJmx25S7NZIiRuJ5+RqeIy3TwS5gzfM0ucCuOb+kCNVSe+c8WmsJjjXoKSyMOM4q3PN83Je
sjPLziYvcrQXjGBFjqBqsZvw4pKFSMWaFL9v0s2IH5xYHjnmh9p69e88wxAaSCNH1dCnw/ku3FuJ
PeX2c60GdCwuoCLXz+IxcWAo2hkekJEnPwQqcQ7P93uOLd49L6o+BVeBIvNfi56LiuGYzZygCPSs
D16GPRY1z26XRLLfpn/ZwtkyuaMbUEyx7tapxxxQQ6lzIJeMVZraI6bKIpNZlDoVDKhKvEmlUJeD
3NGfoek+vJr0g6UzKomJs4c9dPnwZEyuZL22vT5gfZWJziPQDoTnOFNW7Z9Vc1aGWL9nGteBAiwH
eIkClYMn6geDoEyAKDGSXZlWSHbQwskzk20fe1hpog7DIQY1icV/+176zin+tNMS+5jC0MDxA4DQ
YGZ2hOwdR7BSs42GsgO4Vv6T+Jg4IxGDYixS4DuZNDt4XPpbHKaoqBh7sbXzvsxnjut6Cbf2eZgg
KOABdBDsXI5OH4381UJfzu67MlbQiNu0wDzMo+ublybg1Drf0gle7GBc/im+3T5ZB1Q8KJVdeAEe
IhG9VjBYQ8CdUIrr7VonUU6Rim8B5PYq2KplL5IaQov7BmYW5hHmHUCZH9l1qBpASUtgLsqyJbTN
o2sl38xenDG+6dwyK/rEIADXFwDeNXXzL3tr5JiwJ7z6Z7+13aH8GiSdSfg0+0GCOk+y68+wGZBP
lG7QNbY38SGxYIXpOispwx5QMlXZt0svO1E7K21dDZOP3TaeLghEc29rdH6CetxIeg9GCWvO6CB8
hr1Iv6bI6yYtcYHMVvRw3gAHKPrGnmkFT94XK0kGS1B8QTM2jRdgz5/0iLjLCvO2CxksozemYS6e
0XOrFHafOWB2ENjOMPCGeNHAcW8WhrSh2cSjmElclYhXhar7bYjRS2PxfHmTXrwrheqUGGYYhxWr
cjpgauGuD7RKgKRzbOIQII5Bw0sa/yR6DcOK7rXm9/FaR5VlXkTgvyaryc1EilTw1vZgw+urBYz+
T9Q9W0ULOKuaPKx4uOKaufZfNmhuI8zcQ3XYNBQARMBpFJ0vlBjSNjFuGr+U4GS6H4bS7ico2/rv
d9CDoJ6RC1DYhF07N4kniN/+/u7QWnySSJJaSoKn8onGJ7GQN6jYOwfwtF1oUmH3f9HqBUigNHGV
AuQGhZkcSDJopeHWU11pGa1s6fL1NhgVhm3w1gaCFFNIjbqmdGDjQpq2XXq1mI8M4qx4lSvg7Xzs
q/TojLPgfYkO34NExDC0WAYuVC6NdNieXPmrwP8k+7ru1URP+0TebkglnqdOsO3FXwPOI3bRMMG8
Vofozqqtyf8qwe7fv0Dwaxc0PpRkQTSxKoiYNhrq8VJMpGhr/lCRHKkWqWB1Jlr7dSBQ8jTiSTxz
2I7pCKsPcnVmlmCSU9LyCpy90UdTqT8J68mUmvbxjQ18fbhrHmM6Z8j3qMbW3be8RcHQyv06BAU1
zWkUDcIR/LKuDiEWKASk71rdwGlN0xH+g/5ykNOymuKZbHRGZ4I6biNb8qE1eFNpGRWtRqUuRlIv
E/DjHzmQXNPIkKN83Mpi5ay9n8MMLXON4YCJe8+DbS/zY3uk9lQRLBeGRp740mTqLw94+vi8PHuW
51hNpiXvQzOAFLPLW3L+PCIUmBGJsf11a+6h2v6+HsbE6OXJN5yQk7srjyryUQvhiZYr+9wJ1E1K
k1MsINc0BWyx98JKq82eRzuDLy66fivElBsqBT9ugeAG41zvR6x3Aim/+e4vmApkwIuS6wk60ATT
+bo4StT1hkDvgli3gc5Ri8jYMKS3EYBtG/99bdhP+6u0wAIj3pVpYQ6Yobn0/lAHmlNelBuYVGjr
hZu4QU2H5XjzVv8ll8GKPBscnQfSLUqWAHVR5j2Sdwnejigns+04dV2vvM9HBMyHazFdvgcitgEq
Defmg+ucnZB2vkH425DFXTg2K2n/Fj8fkEN0j55kTRa9m7Bz/grNOM0ECei4M8ULMVUK6NMXrFMS
d2Si0FEC4V88HktXYXlhkd/rMvgNoOhn2fMYNysBN6g2WBvves+bwxUNe4JLAlC/Nc+q3sbZbpE7
+Xt6ls16IFeJCrFMl2VPXw2C2RKMKFpy32z6WJc5Et1lIvnJQZYvtuMk7uCzmQ23P13Dlq8/CA2W
NXBKEa1Xz6AInml8foDMcvsmmq+6hRzhiaFrsSFiLr5MRSMsa8z2y+/DzTaZC1hilqBtqEiutNXw
0EAwMCxHeP5dWs51MQhe1Ye4XwSxkAa0P31pmOuQ7bCZn8a+tCn7ogsptgbZr12LnZ0cid3X7wvy
bocnXVs2Wa9p9aTs2z1YYFDDTPqTJ5fIRPB7tzeIFaN7aEaXNpyAJysVvt6XliUlAXMf517CXUzS
lIRHm2VoljntpYPMb/3tuazk6q4TP2HCAYPFaCjysARdYAx5X8AXZtnYDKaa6vlzMLScDzPqBJQM
xsW06v6jYFZsMGbj3hzDrsOUGhu0lgX1+AsizHdVHyh6Nc1gqmib6O5uCNVOPs6EjXxWxzb3r497
NF3lGHNGri0lJ1IeFpOecdhATXIEqUO6KhORJXrlb1iW5Eo4w6LXxb/dgB6xPfJm8Yj2FYRWEWgI
fFOcaiwb48uPgW/qSABY2o0cVhrVdl+KK0+cnuwcwiAGvBAtNhELc1L1AXCd2iPSIn2Uet/eNvq+
IbKZ98IovTtKSOHQwBQUwPNnEf5vKioSHwMP5lrbrmuZjjvUobTdg4h14olcygwDdjAgv5hC6t6N
mwt1MZROtlHkiFRSTlRmlgD5AHGa1fn0UqANN4HISOxFjGQNVaGY7UPmF+8vKAeweDmZRWZNuW5j
dkhQFRDNeaPIbkjQyT7+9ctiQ8QXJzu60LvUqpc9iGPAlbfZ0of0osE+TwY4aVCHhkSsrhj2xyKT
0FPNfMUKRWYkMq6x027QhJfwZd5jliwLV30pahFz7gmCZYWQJKyBrXcCceH357iT0hhUafz1OC/Q
KyuUksdjchA/efHgmvavYhUBlpO/pes+1GcQgjPwdpKlBO3dn/sR8q/clYy/ja6sgcn9ro1kA3/9
ik/ANRIu8U+Kgg9JYIuNUACmVUmOj5ebzezUXkeCWPaUgNrr4B1CYwkHTW062SyPRv6dhLkcZSDB
YWcniLJgfrol7+g6wE0tR/Z0vur40KcFECaBWxYRB+itCUw8qYaCSiC8S8rM3HIVu1H8LU1cof0g
nkDFYkzJOn2W8jdBTj+/OdAZOQ9GqRiSYy8HU61MLmTvjixntCpVkhzQozRH2Lh2H3o8o7JBd6VY
RGvvFGsZBGw1invslvZs+X3bK7evct3UJoASAPQ4wvKFLwf0ZZcD87KcofmXQXduDcddZkS1QdJx
6VzxeP2qZRCqKueiVLZ5JyP0ApA3sSDF05l4UghbDn1C5a95xNCyRIIl7VkjSZP5iSpL39W6/b6H
l0GEbj08cNzR05FlEuXRFBdxokQzmn3Wat0z1pEjP+BVgkWrq0/GhL9BMEyapTCJpsTIzd7PvTh7
Fo4/e56YY1rylFx5/Eu2fquBSORJE+a+vQXzINbKARQOUvZN6rhx9tnJle+ufH7qD+b7uc72pTW8
97EHWrFkVIJr7Rky0opc1AbM4+nmpJietija5jhtyR51NVHsaOzlvvMEYnKdvTjIGGP75Lwvz7nF
8+PpK0pEgppo++v1FrKVMGg0VXJgWBmYKTbbWMfx6d9jm0H5daCJ9HG4PjQxC/U7CeELF/7hgKS8
/JrC9suWIw2lPcaCmsy2168xTmlZpsTCHZwzbQmg0nePYLzt2RcVXH8F8G/xt2O9grwPaBYjtOBF
7TU1UAGbHtp1pUfpoXyqRye59BNs7xtrIWAHVHm+tEDmc3TsktYEzDmUeLA1jNO1Gq6iJKYgZvMf
+UMDjXKxwtCZ04mRRhLxtCZedZ+i8BVEbsd5xWWDBj9ubcH6evjF420/g/YXe3PQ4rqQvPlXYloh
Mk7uh7zYoy9ipKhiPEzAZ+4tXmD3lcNr6RQBtDClgM9Jbl56WZvv9UUcU9cSxXUtFJi9HHmIVRng
t6huPOPMlWTd4px88FU3+CXVOg3Bs5i8ssYFO50WMx2+YQtghDhODlS8/za+HnLqRXa1YbRhaj8u
m044SNUQlPzfGeXN52NWkDY96kZgKtId9maTA6QSbMxtDArBjOiEM0mAJUS33Y9FwiAnPT8FkJzV
Q9pdN6/Fe8zhur58q6n4Mx5vVCEsee740VH7bUMbZnDlN7mYNWnkopJrqUCb1F/M2Ph3BYmO21iX
eCNqWn/ASyGSrKePIP9AlwyVyNDcMiIuCX4LMt7Ab2AIbp8nSjybblOGcNVMa5EBOD9IkYrc9a5D
IdfFf9ZClB4f5H90tl2nhexLq4m0Bc6d2jeB9QnUpivDxCO60H5M0kRD2xNaa41KGrhH2cOzg0aR
A034PaqkXZ0gDsdDfMOr/txwj9zS8P+vCRBHCDouNd62ahH3MVk8+JaCAX/mSKfK1DjdqnBLK1BC
2nXNb95R12enF7WZXl09ByhnKOF7PFVIXU/C9ZsZV9ELIyC36dF+VYtqQfwOfTREZuCPhjLbuAk9
vHsNcVsc2mKIgFrukiA6FvsbODqbp2G+tSib6Ma4Yx9dnVpteEVp2whXGYG7o2B//uiL9brKKVQH
4NgCmYiUQ0apV+sxPGpLL8gnde9JbTFeLbYCGBr43bvQ5g9qkTMt6rtjpwYAa+oMZaad3sYqpR5b
v5sPY0yXHVDxfptvoBdH36qN5YdRtkhXjGVmifC/TxN06IU5l5tsntQxmmvWRnHlQ318WJ7fg5PM
egr/NPythIR5XJShBPSBjLm3iO2emJ3Bin5kwE0w+fBs+yLkDBom6DcQhI6sVu4v/wsycJ/FgXTy
5eT+Ka1mMg220+MT/Ywnugf/SGAhOg8vdk+oExW5x71a334vqsvr6MR5UgAD+amVhUjUQQZyFauv
7xf8cbXbxY5lVCIUZhCGutIaWQzWDgZwrfhoRXIOdJsEzYkS1/szA4OUGFSap8RG4p5eNtxc+5Ub
kr216j8EABQqkRzwBscUtZt7fCSAXx2ytB80WqX2CRMwlgkohsYjOCT473qpBvMKodcLU2uCLLox
iaQPFXvIAVaovJ+qvBqI/SDNaYKxytQim+FWWE4v1CUo0trUZStFUoYs8cfcaZkqGHAdJmNn+2Ha
9izgAdPqhzjrJq/ejssbTzTuSqnQgZRMUHyUuHbZiA/ff+6Y17WRezB1tsjRxmzhjAVmWZlEy4mO
SIoqaZHP9tNDYsY0GL+SMp16HvwFB6cB/ST6mDeoWP3foKGsQDpjSuZna2PLN34+q8In320mFOr9
YR53PQbZlFxbJJDJjK7ROFErqcqwT9svSPukDSkqnXCOvGXemYNDlauiF4endwxZlcFSSPodBXBC
dB45CuA0UCoehuOvv5iOIeZNZp1ZEXMn9Qb8XDgvIB5CDy1h2ZLiSEzWj6QX1fP2ZeihonP8tBNM
cIF2K7fAHZvyXHiJ8rYcmFkHEWdPIdG5G7uEBC9HgHiaA7N8AYeijPuXioCZ2ss84U/nSKX6s8MW
KIpsWqqBQ7RgYx6p8FbDQ47BKB/HoHbrK4utgMA7WpbpBrBiZwrHzxbxZ/n8wfJTV7ryASScAEMI
Ulcsd10N//DYfb3wo+D091yCUmR4gmwpERaVc3fp/cToBC1YDMTvd5lUzYu1Nban3ggmpcsceCo9
NTbAeMCffyFLYohUWV+9To300/RbSGK3ibdAe8ZgGRW3BCZIXjCVQIx3UoEtPxfg9bYXttukcp79
zD692VlejoigbhlcwhXf3Iuz5V4tYWauQu5/6KJJD4Q9L7sApagOoJIo9ZuGM+2ceZkZ0WIUzv7n
Cbl7YW7Fd5BI2BNe3irdJUuprQVOZ3eDsddUbLhpr5u85tqR+g8NnalIEC003pRmZz3/4Osyn1G4
BZihy+wcUa3JL9qvsHthq3PO9ZTxfLyQN3hoVDjGZHhwR5rPOD8uu7LOMfSey84ZVrVvj2Nbm0KQ
wuyiwBWju9YdajwDRWQaeT7Y4xaMJemBLtJybAoJMBmP6CbTLUhTXiQ/SbT0EpYsx7yTX3FXFUjO
IP7KQeinrguCAg35zesiO2pSNLZQNlrbVM9+ZF1klRbXBsxF1pF5p1dGfifbe4qZJ6YyKcUPAaWv
yhJsrpxjjfhZh0sgx3IJlM2VOtquw28xuhcgEEZZ+loozrKoJBw1BM1oqAcyKQIhg1hMsiiasjkH
dYDwm+EhBLZ0sjDKORAfPOT+l+nfWjRIF5iYyuEDtW6axNHKRwHBNIVzBboryaoDOTpA2o7jYhOO
IoeMTQzx2lJ2sgGZCGG07JvctDuQkT4Y317uQ7bV4T/Pr4EqDz1/vpz/eszEb8X1R3VHOd2DiNLG
iNLMTvyyhMojHgTaVhzmP5JyLBcl94fBkLcYb/ZS7bNccv1KlmccYKsgMahVTi1JBV8+vvCOVVNy
fd8qtashjXp4+37g7xygbH1nRazJIOGlPUHud9fOsSWOOUtTn5t9u4fyooC7ibuZ4e+C13TAy60N
6mvDzBVbbValcoFkRWzZWFxNwmjJEZpqGeQk+MoU4GJLM8bd89kDkywOncHxq7tYQUDG+wkaPHQP
zBaJ/dHnJ9dct+16boStwtB//s6KU6ViWoxGEz5PtyHC23D315aoxPEc5GV5ATb5tPE6c/R1eUsk
k6G78D/g5uASEb006/PnBuRI47XQ4YmQoBNS4DSHk73UJaD2OHbDJIMZL5kn6BWrVMTZnvi557Tk
vFpeE9x5qfjihQmDMLy7A65f5CWAIX1apxvqLWZux4Pnx9uqT4nusR6qwFCeSA7Oi+88jG7jse/8
IuO46Sfg9SlGTFuXB1yFvSNobEdNYJtO1myTqBjchyhGsSQbX8VE1ZDQwc0wEDRhwVCj/poIZPP2
I8UVxOORPjGpV1iDiP82gslqTghVHhg0K86oX9BKZlYaHz34VxNq4qZuhxEgpDkCPeqQs+5IgEry
rlIhINe8m75o1pITAIQRSjargECGSTdDvjlSQZd3IYW1AhgA5qyE8PNrzPn7TYhUtQG08cjGqP0k
qNPmYNGMYlVpWVpNZ/If/myDZZCq9HQ2YGKVEG/JieLZk/Acbwj7GVFwCgknhzZLKt2vnFXZwzIF
+JjSuWGgqX7l1zHgvQ7CNoLmoipmv0/7YXy85dF4/0nwA9RK1M9HTaoJFeWfI5Bld7ltf7RjYm0M
82Ykgn4tcvGxwizEaF8nDmSBJl/fg69sf3vn723RkRMyQ+7lhS/06+J/46ehko+Viq3nvVhkjM52
4mS0IXv8hIZNOoTokaRxEwSIb5E+kvQ7uoAoshyXpmaGqlRCU3nyHY3qN80BjhMTyd9Lv6Lk7tcw
V9Yn88qmEutuyx64Mp6jfsO9Ubq+XSAp1W1nAwiJJXWoZJncev+D+jjqves+JC3RPtQ7nlHPImhB
jjrXX6lc+04oQIcVZusxBgPmr1vWQakbG2U9MPHunNBjx0v7GYLrkhL+5FWRGuV3VG1vgMiJx06C
eA9jgiXVwYk382Syf55gO0rlbhgaanGzDDHTNI2/9dTwIRl0zEg1n6B1cZu+9Lnei0P3+G9Uur4d
+EZAjZFdj+XdcnjMqnxg0OYSwXFtBbOTuz/bJ1rUjXwVB1GhVgsAEFBFXJpZvGLn1//tFOqrQ23D
DPa221k8rI8x0A95hdThzdzDTwU6B5kyPJoVp3mr/Cs4KNx6ieEc0gdlxJ3BWdFfmBgbUXyfe64F
+CxTZIU8yJ58XYQ4Ymc7iAgSwP6XeWaNvKYorHsKXHCBAzk4msBTzAZpOSNImkuNMdV6cjBru4Jr
QwhACOzgFrL6fMmpVaxQRVLRebRxKcIb3PpPXhYhE/GjkbWWIalSetXVbdtlf93HRNbgIXPbYGFq
QrG3F/EOkiiomJxzD+q9u0n/9WmLvFd5RKghPsP+Tm0dPvVbyhtLASsMOoNLyqZbRUyB0fOMm9Lo
9f79zDRwkz7kjxfQJyC1tLRW5a5JXtX2O/du8yOnaeNoHMoTv1nmSuYT+Ysg5Gb8nJDupvWD/1R7
m+IxyQnaFNjyuJ9zyrHCL5WXuQ2Q6sphLpxDN6zHn5LtFSRX7Bn6kaVS4+cBo+tUAmwpvKG3PeSv
pFcFWEio96H9pF0M1S4FsloLU7pqO/RVR6D39GAeVtzDYYvbTJH5NFT335wI7o+8IppvRn7vKyTp
Jz4zKGRy+o0YdDe+BWoCcaw1aLC39zVODI4SssYFzeYhwwirMt5v2/P/CYfV8SddK5yqFjrYzBO3
xgKvP9yw5nIGtZb4wPQ5NaT8ccX33qbCZ1PEQTEsFWZyI9g7JAOzqWVRdk8gwUjsMj/034cxcOSJ
QnMWh0uCVbwAwjJZ0gl86HZPlla+wQxQcOT2tHakN+yEmjpeilx4Wo/zIEFc6d/rKHECJj7OIE6I
olwJZ7873CF5piEE6VTqBC/U23zfW3WdePpUZjVzXT2m0elmDPNtJIrIEkC7b5QCXN+RAPnaNgOx
VXjNEKch57h6+Fd870Ybsdd6sp84SQAdRLQQCdY83dhV4BjquoImHLifgJ6RKs3ynSegZOR7IvmS
t8yEQqLHhpun05JOFWBJ+qF7wGSajMpG7jZ6oD0rzyw5f7Ue6JIkQw0fQod8t4QNSriXoO8w6KSn
Nj/2eLJ6HzejqRHWgSeN+jayhun4W7yKoMyJ+5WeI2LLDNnqaN9QFJgTSp0WBe4pjZI4oGspBw9f
bmpjzXIV7sO5lViRlKnQvkJSrvg5TwFdYaLisrXTtxXF1A7DF+CzovsLmH7kO5mvyf38YbfG9fLB
CNVu/umf55QylczgeEP7DcTwEoJZVzqugbaQMMbW6n3VlzBq2KuKxGSsQpZGPQ7tnIVgzQDvMCVr
TIPshj72dfwgY8S/0WzqpJYROfxSVu+nXrCwvxbf3yIrDMpqhUC8bqYpxnm53g5/jbHn01XDZjQj
SQrGriAGbRR4gw6QmeQNRtOcxDyzRYKBQHb+iUh0oj8WzoxBS+6fn+u3R0/7YLwvzaFYRd0akf/j
+dz0tXnVkgH83qh3WgPHSnhW3TSBWH8CbMhbWIgLq/9xBN94j0ziwXcX+7JILqwccNpkon5bAcJR
4N2oPOFYPrloeSTJSN3QhvifUji73ehjPcfJSblGNCUR9QIe18zP4Es/ChEc2JgPExhqS/XHzY3B
ugbY3I382NwEcoV2VPcdUuJ+bpxdv8MooUlfULLSdaKuJj0EmZBtEAtg6wma4Lz89+w8meH163aN
uRW7msxYcMO9mO+NnOIV9gex7vH781vZ6tF2r1FSqEzKSEERsa2Jzf/Hk2LOl7aPPEIpP33QgWkw
ULJjRoweMz8GqukPmsYAMugd8Vhrp2lNZdiXgXdwY+aeBJ0LysrY53KlGbRtyH6DfDvl/jgF6HUS
q3rltAZ2SXtCgNf/8C4bm6+3bmznUOQkGRQH/bRJkJJP6suGchhlgFCrEZ6AMM8+i5C9CDuxjVDg
sw2PI9xuLykHLhORILTpKJCUP+3kUn+pMZoHyun9yKbu1WVYYEbwFJxWYPgzaMHVSDVQ/pP90yfy
qNEnNrh63ST9xWG/9CgPVxN84dqSGlTZX5hkiUHbfin4uiA7tXxb1cY50DIyq0ob/0Zy/ZaYkuHI
KGgaA9Z/jzURNftuMGYC6vuGl8bl1aJ69L9ETSd1hCzTdfdUcldaHVAAaoRp43I4FGMVVFzZ31qe
Fv2FwpRgjiJ6YgoExEm44W+PH6k9Qw/03u6uvIsxtP9SY47QWXBD7ga/h0vE0iZ19qu2DFJldBW7
ZpUNhrYv+NLXE1bg6y6ycQZsAdI5CBE+lcvkIWVBu6euk6mydnvq5tTwGn0m+FbYFPko8RXxmsVO
CrSvkeA2bMhizVIsoAxmqx59+53MsJj58O7ZhoufdtNK7igBLHuFoGLZe1HgjNN1oUwQHsZ/WSF5
9EiNgS3tWbvs+e/H4t0ru4MdzEBk4pb+C348JiyCitv1C9KVQI+hc472KvtbybwtLUkVx4eCeOtR
UWCMdq+pGiTWNPnz2vDv6KdbxlUJwhCBW75Ix7CyH7zkwoRt47xGgpl/jbYAcaeB/XDtZvrhddYA
6ozdm78tvRTHDo4Gi+kfzQWwMsvXGRQl3OcFdGdiniUAJQjiP5FejEVom2zn/7m1cMSI/TKiVKXI
70Ae38UAMLe9Iqj3n9SoYPggQC+/hqfRA2UJrOuuJib6bCFkG0jwQQPvk/nXuC6JUgX2Gpyuo3HG
73diemzMEmjQ79yUE0/Adq37P5daAMNucUGloKvRrmRYcV/DUcVrWOyU1lPdrtacpIf4G1kyypog
Z6XzctRi74CaAEnJUjM65cfEq4vTweanH4zFQnYCSP2dWSlBJmVQgzm7gChlWGoXd6b88BsmnLCR
z9wH8yZJJ9V2EZV0iSJdxF6fP7i2d3vj16iiGmk8cPWZ8c4YC5004PvxrP1MNG0pwBydR1pjM3BE
+zRwV4h1sV3jBypWyzXXPKFDnPnkU25WpwkpQhVu0s0qxuWOmsUSafHTGNJdN+0TzubrLsDaJfHa
6USFPnjGkNFiK1TzTFOU94aZT+NYbUYmEc2aUz4HYgC03jyVpfeHTiqxojh0aDAp1oV1krAej8Q6
nFuAWVi9fVABD+kOWp8axdGXg7SsVx+VsEXDAA2fARVIwjSNSuye4ySN3BmJCKLZYNT64IovPp9i
oY7dR2DeCBsUe/JeDLsyRnQHhqSpWbAC/aVroy7Ay1qMgM5g8AmII325He4pFtZRMFFSmIw3r33Y
VFG/nhjm5GBkmb3UvnqaG39Fw8aLZ6NP0Eem1PnU6a935NERSHY/4JOilY8jmwwFCvHo6Dr1lrwU
b4/OCJcfFiC6jZgVUhGrtnqUWR/0yTB7p3nRQSsnFcujNAsGdoxB62KYtd5BVBkcTkUY8BfkM2Aj
y44QWB5HywoHg7sVoxARYAYzP4frc8zvwdBUBgctQKmsKq8cJmBUElXMnr+OiQl8UsUy1olJzBrD
mGIzeGC3ckX754fvwqi4rnHqX2v+bS+Ains/z/T2ERf3ciGAmE8DjTgHzjKov7xzFLpmoAmpw2j+
Oet9Ou04K3DzPDdIVAMaios7ehfb6TfkcESSaR7mK8P6JbdLU1wTlpqaNll52eAZ/WaCNao+lHAQ
ewgVdshwG4m6hA54E6mmeOyxuBKIaADQF6+QbJqhTC23biT+Vk7qIKCgfod66EH5HMeb5Rgw7f7/
6ldofKsHoZv+OBxyRKOwRBkqVxuG+ae5a4hdJJD2HIE3pJ+KPWu8SWQqo10Zz0w8desMtfWjHTr1
SMhWPh4zdPMcIWP4ANPYcPfVveCyS5AuQKExLqGOgDithGYyBu8TnXpx/FGgvjlVGqwydAvTxSGA
OzvlOts/c0f3blVDNpZry8GPUouvYzMV5SjMPzu9dhLdmQXkUWc+fhAAdC3SX8emJkSE2AizJaCN
WxdycLdkz+1lXQSSYM906QfagJg+HrExIn0xXFS9IB4jqFSOmUWjXEpyTh/LIll8Ib3vQ/vYrRCp
CDUlhS+DY9djiYEQMHDgD0YjYdZ395QzpanxCe3gH/YREezGlFbiywhvGPyoNMpj18VfxOlsKng7
MWfxkhil+w16eyplEp/UkgkJZHjvW/Rw19+XUWB7ykI7bcQ6ZKYmQf4WICCT4JIPSs27ra7/tllB
ZhaNM5d4ERcvEnxhTF2UWV9wx6TaZ2fVsNzEvgsAUzuIBYUr+0/qAofE/uwsIyj/II9WoQ72yvvn
NBzuXzCvZ0OnmRgoqKc4B2dcnZwuzarRFmH3xgji5yEASvX0OHD/6HvkOWn/9l8ZYKm619sy+vgq
P6fAfo7UiwDKvOwMHJ02kcNmmENOPmLB7js+RAV73hn9lyQol0ykY/YXTO+FC69jS73DTIPYWORi
8wAWQ5USXqw35hrufMNDxzJ1otJDhOTYdDMtx4VBNhXhMSodK2v6tTjJm3ArXKLKqvi7Lo7dwM7g
fO9Q/VhoySGaWR07dvqWfxQ0fdC6RMN+AL/T3Hyt4bJhIZgL9QBwVO7uUrUrxb4I87m+gqw6lX6f
ds2dpFTz/YZdNEBWyzLfbExnRIhis6CFzIkphdS7ol3Wj3LzevUDo7xtv/M/q2UVNQ/CHY09BCbk
62Y+jVL4sbLyQJGmSse89UorM8d04blcbuC7YZxwyx3fRWJTUq3QpicM9QMSLxL57jvcUfpHLv2G
yQlbmE53JQ8BiEychwqmWYFDqncFG55w5sSPdQfDN95IyGe8ca51JWfODkgRNZu58facAvgWVgwZ
yPYMa+W7Yyw/abeYJ12favrYXRj1ofQlygR1dmSIwEBJPLD3IfUK22W0e0j9hW7XuHn5BXC/z+tL
XhoBF9bE7Az3AVY+lMDSJxMsyy4LAqTZFaqsTURxnzHBKF0f0Z/WITLOxwMOJ8/Gs4fhM2h3zUiB
cnpIMuyBB4Enx23+xRu1kzji6LScgLvL6FBXMFl+gX44EebjQYz8FubVW5K0v8I4KSno82cLYMwm
C/6YzMqoubLbxfk6iu9hjgpb6p4+ozvbVmKpI58BGIocK9qR9FipdKzZ+iTW8CZsld6r4LjSM0up
9+9gU/eXfJ6Di6e6BvYFC5hprO7B6aEW2QZbxzSV9CDfaOJWBQFBFUZ0WzPEJ4OH1qVQoO/SVCh1
yf3nvUThPxaloUfVCNwcUPxET5aHQM4AJRXhJ3woDk3LUa0ThK9DMMJDun3nIuvDPpa6kv8Jq4VH
5Un7tQShZsWuf6Thmj7h0Id2XVGaIYjTUXFHhVXY+wXBJHafBysGnAuqtHf1GAPNdl1Ud5u9nGeR
FtDP3lxtuhXOnmWjHNl/9dQpD6W38PBnB8SRB0w3W24iUQVwMUwIgr7ocwzyTFXzUkbmqhC9T11/
B8j9xBQu+01Q+F6BN9BHvOd+z1yP54kh9orX/FmzyenGqFkQKYg8nlAeS+vBvqTNMV0W7XKqOCkY
xE/0v0jNP0fS5VTFQDnZGFKeaP6qy9gdOGZjrIzQbY5oXsi3o4LPydUhEmUmshitiFJSgFGELIXG
EEkF68g1Vsje1eKVZb8ZVOa5fk7c5rSzm9G8orbF4jBTQD+mWrOFjWrtBP9so/qMFVuQxilR7tG1
397PGkvloqqcxwxAXZ3X0xLnpKRLrxJEcoOqhnRUipDd8UqCW04UOCUMRtfKE3FhMv2GyisbqR5S
5Wb4KubBGvttk//g/fqg2RTaminM131VlH5MgwYMllIJ3c50ZlLMtFYFjH5PFPHqx7+OcqzIH/cO
UrBNOsUQM+7EQ+ciXCLjGc7i3giFQ1W+9LU2eFUAprbpeXXuJBe2joSw+FaMOCqPlg/2OYjo8af7
q38Yiqd8JgRJY4NtSD8gvklbrnR6+Em4vuNc6kAsOsray/MTglWnL6x9+ynpTgT0zk7zyMlbIQuB
qfxoI4ITbZ9gAQ2k2g0TvtK8gfkPAeqU4qHYw19s+MJhcS30E3DViZ4CseLejBxMOmLRaPVAK1dD
n3dzteRc5g65r1zhR+GcP+GYA5yFK/WmctdUa3FEdFfqdqaMopdlpRtguI/ONKE7mfFzt4bdLytw
KanNGslF9kLq+mBj6Qeycoapy0ox7qR+fpm258lFX+ch82Akm59JWyjUPsTjxB9A+PJTn1bjGbqQ
Ld7ZchPBfoTMB/pJdwWcjLtvQZ4PWKdwK8zgYJHQf3sswAQTrX2pRc8WPl636rSCpoh6z2e6XLd9
kG6YZINRdyzFhHPKyO85o2f8lofBpvDiQFpsp5DX/kbAgtWyU6a8WZNV1pjGdwL3RykiFxMnYEHj
dYoMeUU1ZAIyzYb/BpuIBV846K8kjVvkCNHRZNq2MtXoVtF0kxqSOKGE89mDTPi1CQMBWEN36qRd
RZKLQtQlOVCVW6XsZMoliTr9qVCan2Q2KgCu4UfH3A2b/mwGT46K95LqcvTioTaCrHLETsuK5XBK
puJnoXMrDXx9iW78/X3X407ThvvNLiacnynsSnBd1ypAwkKyyWLZ0WXhEWVtyv26d9ZR3Z4HaW82
qu5KbSmhUKpIC5CLk6qgL6eL0Ow5TBaq+PUhK0SLYmXleUnFLbDLUSzErc6yQD7WW4sqKJan5qaV
Zn2vTGkMvTk/Twu0bHc3YWbLMHLUcZOfsMPr4hASJFQRKxJb2V5EoUFABuasynwQhBWOIdbCsUNS
u7gHLFjAl+i/LNMrEI8NsJI17GmDyjGaS2WF+fRG47tLgyXq+lABO958Dt5mY6dtmn00flPTi3JB
Xth3OkRL36/Ce9RQP7W41l4YxjmJvxve1nb/L5lgK/JEu11wM1l13mLi/gPJLqkOort2mdvHNVXm
Fgsx62u9SmOeFNTDjSH4YZbs0WKfDeZJApNs0ooHlc0AMMY4FWEt2X33gy7uY13Q0oiZ12BAZuIg
1TfbRJKzEeipZtA8n7z65RlJPd88DNl9Ro42GfW/L0wSFa3Kal4d3e/CXET3rzAFd1nhNbzNe49g
5icD0hX1A3AayayskunI1gNSDmEnACJjnXVBBx9YF2knHR6A5lOErbRkR2xg/zhuuhOuxwE8Xt+K
dHKHNsHKUwsOPj0C84BcOkkAngLd9nwzU/kMapfjpWtaLnV1q4MEQ1nN+KYvGV81IQFkXAHHvvMt
YQ8vuCOmby9J903B0W+qqjuB3ZGyAOLNbkJudpTiEN14A0eaooTdPccdVWGn+mMCQkxXp5csRHQN
lhjVIN6b4jc0lhTOJSA99dFwyxfSJdvKFTkMQ7KCCH/NWam3+J64BtKWhBOW0MsflzDHRcTSfB6F
yvrKqnzEss6eY771ofFWpRKoSOKy/7uCFyyKN+Ekz3GZppjfovgW/WWx6DMNoc4mmVFC0uiwh0Vm
4nU64dFy7EfZngyiwQ+PEd+8ANd8TSV2GwvuxHcv/ztoeto1g6lxbF65M9nIK6v9v11mvk0/r3Cm
CynAaXDeixHMbragt1ddowCDlKNiwUt6v+x2Afdht7Fz6FuEHMSePPCr7u1FT674XVQWGYCV76N/
WIg0e0RnTrZwmyHXIYGOz40WkzNXEj5hhutNn3O222jjTxiL9bgFhYqzzBzYI6qAKWeQGaTI1GPN
4t8vjTE9HIm/eFKAuMLpubCFsb/zj/TDOLoTOX/wWauqiM5gUtI9ajbt8Dj2LykecOVxcU+2l6/V
ZUjYSnWCAVV8jQzNmoVl5uhj6+9CUUrsZQY1VfpXo5hd7qDqCXOTm+6TFxq5LOYv1XveJvzpdDwy
kf16GEo2zCrLr0liWY8KU23kSr0Pw/t55nrEHFLX9XGp4MqwNWRGFVv2juUBDbofnaR5aG72orPU
dYtLMXpJewGeAzSWz6kPL/Rw2MY/IAIaLuAYESf9HwRSean43lINd/38OXwo6Pyc9R6MvDfaWIZu
a47BI9S0Ap0eyz1+15x+eNpLSZx/6Vv4VLtQs8F1gT8vl9MCpU58aL3I9oCkBMyF2+rsfqCNQ25D
lzfr/Tidb/Tr/CedI4QDxEmm6oDdfDcIicw6UjYdpjWvHTUIdhz7r+ltp2zGmVOJHND86CPeuhKB
fY0uPA2gWEIRFxnXjjCExsrxquiQQb72fQpCvM0vkF7JjBen8roLgbAUgbyeZwWKa2YXDU3TT7D8
ZWjauD0Az5Jmdp4rBMPqPMqKrCzu6qOUsphxRZmLX6jPwp4nKETJzv5xnTPW2MBeaZo+PvBMJWcC
yc9mxV74Tag14EHCLmafBiAiSWpvAcsOSzek4vgEN2UzTnw7JRvALJuvefvvWG10WcZI/ZCcQbby
kYhQVC9FRauoE2vMzrfRnL2pKIWSFSoeIOGRm611kIExIa/O2sOJYRTg1cJQvMLANLEBMuEAK/qv
xx0GJzrw6hnoCyZoE+eZ3kKm03A4JJMewj1hVuEzNU7HIGhlW3oy6se4tsCM+QR6/5lDMqjS+Zdg
aUXLeUcBqCrb4pHNzy9F2+g5b4++vYoFPZXCTX8J2PWWJQIQqaMYAX96joZ5IKazxJZhJ/IVJJRT
qXkEYJprQeRlBhh++RpoeFk97Vdz5R2XKnqS8HOUrKl/k45UoglRfGiHtX81Xpf/fZnvw3ywJzJN
+e60abm83U7NcTcujXa9P4qYgo0yp/KUaxMUR+I9OWs9iaGAZrbS47HZCVOPhmh4mNvDOesIUbVS
Jl3G172YIwXNmhIurPNFAqAC8iWR2U5od2ymzAFwfvyfrWvvLG7Wx1F48Ywc5iUPignv1fAN02Nb
ilYY/NFNZR3+d8cUs2Bw04nzdM42/IY5PvacRbISE48cmvuorrrYUjzS8wI7+2Z5eN2yOfhWXfgx
uaf7Lg7qCV7CvSkJY3YnUrr2m9+dZhlNQ60b586e51/JDeAhud5OWwa1569JKe2iRB7B5YPKTEX6
JxeRylYAXSxxnUr7OJy79lOJ/6kXOWiFl/78bWhQY67+0uTxLn072rRJfI/vB6Ylaf8R/cewISex
uHjUteVODI9mgddzsrZQGyjofy9ynACak/0ihoLjlPgsK3TCQgucelPiOZfD9dmd9SdH1Tj73IU9
E/F42HTR6tDMUqiwUlGSWlzC9z5MbrMOmObhz2AYBl/t7G/nKPQ5eDd9Y0ndZhO1JnxekklHh+U9
nURlvgDjWVgNKrcJXOjRE9CqADHM8LmT3iJFZtR5pt9qiiLTk140Gin4OOjOY5/cHmpMbVVr8Bg5
kC0dRCEXv+cml8eB9n5LDXoWcedVY5vwojxXi4WKuHITfurxh3Lv0o2fsjbanZjoq4Xlo8IzhoOA
5/wm3OAbiDQJOT0qaaE3zZ/n6qZN+kft1Je0OIJ8qHVEloHhvGnJFTye6cWkrxQWQNMuu195tZPk
EOX7F5nzBhS5YkDThsJn8LMtFpinPzogCCjTdysCmwMNg4IUnnLxm8URZL6UphCnycOhcBO5AupR
qhznSmWP5hoDNRsxtuxEUw5Z4F69uX/ToWKdnzuLG+XHhcv30ahjmJnota4qr1m2/fFCTGtnK7ud
FvgNuca3Ust5aS3v7jLELy9ExeHkvtIjOTyctllocYoA0JHvH0K4kZXZBxVLbIly8H0LTO1DZcsB
Zkjkaj7JB6OzGjkurbi6QA+scJuir+yMv/Euf+zvwTK3BP0OlbwC4EPZi1GQUQqCHkWIJkWnSmCo
i/kPqs1Z9juw1CRlj53cNxIETaDIMilJ1mvLRIUKpJf+mN8DV3TTRjLNqV2qtfA3mJrHI39nBbhe
ncGqjDp7K8UPFBabmQvdCbjB09qJ/SXiFjDMS4orvVVPri4rEYMFkJY8SjHSrLvcDYKegJEocQtC
sfMO3FEDsU6NWoqKN7PicEQf70B23rRVC8bYaSRcTPM6OfDDY/Hw6QkHnkYXIuk+wK2ak2stl6LV
1eSesPqQRgtfgv/RPQuN1ESyS9phCScO2lpcsvW3YKvBuonwN9dFkKkyTaTNygaBSW0EnVad0r1i
h2ysrasKi32Y3UlU/1tQElZR3ZImXd15MypJOuOAOSvpHCAbb7joG2gx2sSl4HAVyHqlilJt+mAZ
RV8dfHRP98YLgOLpPDZao1AubaKGJi53mjEAu1ymk+qukjCyA+oyGCwvsIsPtSBypCuavRGYs9FN
+zL/88SNhLviisYS0KIFVlVm/d8IAEIAW/5I3sSt4Lvl98yABSfYprUAMI1M0+MdqmMNMDCKObju
7Tb7RLPYgOEr+SaBov6Ofw0oCmrX/GSnEm7yZpC3c5hwngYWyyzvdXwkKq06xDZhCUEOGtyCG752
HZy1IWSMDOkwaGHujPv1aw9HXSpd7cNYtrgux1T44d36cOD6gP9YkYFbam+ddXDO07Ck8dL5YSyv
EeI7wLXg5QLpJ+gBeTMvc2ncmU1GjHjvinxDi9Us3j3C7wK6ApcphxlWECGMdr4ICNktkAdUWrBf
yoYnaNxJu9bfJPSyaiMPxxRx7AMi4PZTpfrIb+ZyLVCJnO/Pp0vYnrB+5cOm3t/3NOaxe3qltBe9
1nIHqIEACCvcEjam18fJEbD37D+a5j5wnvFFWpvp2wCYHpIv8lLPz1PTbTZuoAMBoGsAn0h06pOF
cWAPAJEspnZWlXrWuT02cVPWkG7k0x4vg+YjsmCmWPd2q33Wn8b2k83OS9vzRUtMv2GG6HkQFBQR
NH1OdI3lEWBAr8LSTQV3f8Wo+w8Sainx0utJ4I7adndBVisjBr2JUwu++/GZ1cfTCoJTHsk7UXJC
FTAGob07yMb0EDCKBTnWRB6yfb7bSVZqgpux82x/jz3eAaHYpzv8SmAcep7iVwJskqloF99ekTQu
EbOpiqp+mL70yMrcZXpIWI8xh67SBU3BB+GucAW/fNnC0AQicVkl/EUfPVA2uNTVVDJcdlTOG2Y8
28uSfSY3ebo5x7wTSzMVGJq6jQ3PkmH4RyrEAFioKPBCIawLDErQDC0z5GU5MpvtK6SoYgOMkcbD
Yx/ubCx7jxQW0u3mRighTf+y71X3qbNCdLEISSP6yT+qacGyhsfB7G1zairOL8UvOFsjfDwsAz7M
M6oJ++0s5pZ6pQXzOBiTbuIbiJOs+9NNaTRXijzrbmGJ84CeaMnJAIMdr7qLUw6jZTC/4ThxYSgg
bjIuz3B7n6DwJEF19JQzQh1Xh5ci5tKkHhe/C3qzrpl2b/0DKBkGIFgp7YFwcly1n0pXeaPqC8qY
N9eOI7w5nzbuH/f8H9gCnGUixb84bgjRF6uTmL34ga8DcS3YtBm6k/eKgslgP1rv27Z/Kn+JMGfl
Dr7Coy0pJYuPPz/Sbfzf4N1z77UfuemaoQOkPlUHCwjmwdHjow6MHwfvUr5p0YUQnLXh3fiS5Ewc
kXu/V4HRBYyEr18uc4+CxLkSJimbEAPS70zAwYQtIAr1RgKbgJ9QzZ49eumSfC3Z2B0CVWp0FkwT
8SFvicrubu+BJpCCMIP3c/GcKjTlKJW6qnbFj2wHub70qtJI3AUGFDXP/pqD9Sx/rER0Ef8heRpI
K0unb2CQVAdMhavZr7yXXLBWvtPxcUXLvMgU2pVchx25RLFnxUVOORI98rv7sFQF03d281Dm5fKS
RAsd7fKYiAfpT5wZhWDNQcq1sTxu55NPM9ZzhedfMoudVq97XNW/qmSiJOf9t8SKIgqu4jcSRu04
0RN1HXMbLCh5TP3sGe1ZVr9/1oH7pO3hQDqsXBWcDggdbUqdFWfS6MfaBB0s4XSRIVgoSSugj2gP
m6E0EkqzkwhakN4BoSwgd2s36YDwbO6m9sLhIWxzF0uC0XFFkGnDKc25a/juKhozu2BPPmz4fXqT
pdO8dVWg8go/gs0soe7mg/4esIAaV0a/Ek/BffkQMHOI92BrnTubF1JiU39h/Yu61S7o0pM0ASE5
MTRdx9M/SUcygIQYFH4eTo/GQvxACse0VJoiNRtScQrGrHO21cYKmFq1EyWYPNgVCSkQrvOcxUAn
85SXJVxq4nm9g2wxTDQPdECrkPAryY8hlSn0jFoDsX1jIVzlyaqEDh/W9xr/VqudvwV8Q8MuHmDZ
AZE4Tomhy1eJYFRDVQpekDX0pgy+n4gNALkMBo66mq4y3KaCGi522DnVAcd/B9xBg9i6ecXsCjZK
IQE0wg3ZyOETrfMo3Y1wzNZKSRc/yDxvTOxgTU++JZunNDxfqgo+FUgYXFnBpBn2xahtGA3wZXqK
ZVwdC6d5N0ksuEE5O11m19m05cG5sYuE5eJRWFqer9naj6zl5NrZpJN+zFM+pa6+05f6geCS9mXq
tJKAdCj8UQk21eu3H8cUYfQk5RiaLQuobs54zIGK/zXTOD1rJgcBxf5hxYVhfFaSIroOPu8b9Iy7
C3yhQXL0SdJBi9KgsQUnqDwgKCo+9jvc0rginwXnI2vlqPW9da33UbzyRtaICpApvkJAJs7h9SPb
pPnU0Ms3C2GpFxCBn+IG7ytB6aQaiIM8SRn0OkdqsdpqJXevjFlNyY4Nph9/DoNLLA0AQsFijQD3
Et1WyoU3foZ8rcQujkIWK9l9ZB6t49cVa6Q3FkpoGyHwZYnDfKYoCEGuV+C0rFhuepwpWaj7n1AJ
WEbEFvexDZZ8yqzl/13e/La4YIKgq9kiEBeCRW6iqWrqwvoOXhbzackFmMWOdgsL5MZD5sJi8hWz
JECnGOYl3Kf0cf6UPqT5CHhMp7MKR6ftpUsunjKRJ37lS5cqHNKoQBlPCf1OeYXh8VwJQ4Tw+9Gb
uNQ0R/4+eiWVL6Rps9W/RlYN+oK5NKstLMXhMnOGhlhGgTEpmbmpBzXh6JDRT6mE3lprc9sficZV
Rl1o8ts1SpDzA8bW6pASr3lwwyOj3sYiqLgpQTbIRwW4GrJ0AnuWQzKZoD6N+9eR0E4Uk3T/oGee
AkXE7dVPxoGGmxfc18wPcuWUJ7+iDnwJ1X9yt/riep9tSTSHBXMfSdDCd/0JeNG8sK9x+8GBhjqq
3KwxOkYh4yQnEUzZKoha4YsA7dB7VFkZLbycdtyOO2Osdud3wFXhZKAFPn2HcV/Ej/dDF+4jepVG
es+M4vAzAi1P83aCrxGMwNH0rf30oSdFWpYrhsiVjx2k/XDRLYJOM0iu4y+mVMIAT1eH5dkRqBrc
H34WQSHq9Y1pFysngt8ErRvvP1lvvKYYaAkYyoxesGEE4ryFsHKDBHkmDy30mjkQLj9QVZHF2qgJ
eXInmGnOaHle7I4NH2KfTdt6kofVAqfVTnUX8aSSxZYZ+RZM140t0hftOxH86x89P9XHwVKGoktW
15QUv76LeI6orF/XShRWPeyI1GXmRaGQz67wnfckx5OpkVnDiIpogMWg5hz1ddlImxuNBtU3KMVw
wvkD8cPG8heelOQUhKxcttX2+szvOnPWALNEi39WnAdky5h8cbQce1RvSFy4l7t1+mDt4VEQEaVB
RvVEUhiInFfIjn1Y1auFp09eA3vJEQ+VcsUKGTLxHEeh6x4cJXdg88mD6nfpC/F0zsRYbZdb4qlx
EojgZU/R+4FAhHxwT/xJx0PYR18kq8sa22vWWVDz6vToMIX8yDkH4d25eDFJlVIxDMyK8UT4jeHB
O8dCsGspJbpRupTHI1EIAC6Q6epmCCY92PbSF/5dFt+RJ/qIn9Ak6KlHhA/ahjavWxaWlG01NxGk
NEZBH95lu8SxRyRHAyEz953xGeFJpy3HQTqqb/xdKMOszxEKFda5uNRPTp9/ToIFDq2cPM/7OYiq
lPFvlRQ2I7g/zjZ0sSn1iiv3OgpPY80P/Yiv5JkxO2e/+00SAyGoTX7EGkWdIKDXdduITHolrzsJ
xr71N3GcCc3j9/d7EzTd/iRybk6h0g9naYTQTqLBJcgXRDQOuSPATnBhqE/Pj38d/hjFo/8y9l9T
sQk1Ah5LAOZbTeJt7unZlteaG1tGH/oopugfHJkucc5ly6vZCk0hC+G/xjJAbYgmudP9EeywF3R3
5g2dnqpWCpx1Die5txl2Su8o8IgTUcSPPfqj3U6bd+NUhFVQpfqpkMnoy6uc+fbSt2FiWxWlXbg/
VqmjA75+ihzvmUOJH1mC+kIoUzHLDmd9dLJZkUBM/Ioa6a82NSg2T/Xqn8bhmT9nUL2u8u0tZ9Y2
MvfP8nmzxG3MduEb6vU3DMTxiatb1BSoRPVAjGnQdNFIHpt34251qJ3EEJqLkDolDgsdJqEt0PUM
Bs6LUUaDlNd4vuNaCUOi4Ut/78xEhZ1iPKrc9apkZ8QPC0ZMNL3T3aqoI7+6oB8zKweAE+hOpiFz
9LfCy5zfPy0mvQ2NLDh6gIBhKFj1ajwqH4TlJw1kQpnsfIvOgzUW3lqa6Nu2GRyUU0BoK5rGmjyc
s6dxHyujCu6PT1Gk1nZcuoRxuaKpdwPnzRue8TWdwTPJK5YgyMztQ4wSiZHPH8Qfx9TGkyajmvBs
fVPE70s+fx2RZksrE+8g5wtPARAMrjgeRzyr13XFrtDnvQsRFJELzzPyg1eKva289OSGayNF8Nwt
x/RtA7/zzJyFmrgDE3+Rwyiz6/ulllvLtg4wBH2HH1lGej2MYL1AkhMbEk7+9k0cEyedtlsPzldv
Nptk5+3DeezbVGA6/LWAt1EvRwATug/n97e6SKmwLahWCsYkIpIPY57AZDTyC6xJHdp3cmxPH/Ww
C37hehocx60aaz/HzZAUTlF/+xwkAmr9zGjWH+YnDeCtLkh/9InRFqbFcULsRgsiz8ynvW/n2f79
8daAg0cEjK8z6NujOHEacGFyhcaL8eeaE1VxSM3HqGycX19eLOsKbYomUd+30ITnEkTe+oyCKkTx
2UMilseL4zpgqN3iP5Mr+QgwoSx93pASm15TouDd1ovAvWPCzSGW+W7BZdPF62504XHD8MyMA+YH
TI4k/HJwTzMe7iclLCQ/8Y883cHXdjDV1M5dCt8Fdm92J8X1SKBCx9ur9Zft5VdGeOEovnr48f+g
Cn5Ld2/W929TJKGO9G6sp4ZPKIyy6AxGKTknPYuCRr6uL/TPTJbOxUITZBR2wfxyv0KlwUjtpKk7
Bpr+dattyoUGTsh5d2eks/NQTDtvRQG6cI83D+1lpDnUcYrfnUDVCgUnVtHHBYoAkFDGPnjHx/jZ
tRH+gJoAuGW69NgIwGe8LLH7AlHvLrw6E2gDTSNpxdYsYkS82t80S4Rt1tNm3A4RpRciW2pu4efh
aIfMbS9nX+R2DF1hgTh4xjoF88LucwxDxPAjfF6DMr8/T9uwWm3LaoFbEqwnwq/fCzNlTBKeWBSH
6C0izUotMYWWaU5vs22e6ZXTcntXbAyeL7dpJyk259yI04p3ULLFnDiKAgbeTJVoQYgn4GKN8x7J
NNVKro3ozRg9tnouV/sGh0/7daa8EyxJfQ0Uy6FK7SrBNx5DiS07p+m1vueKFcDpCHXaPRyQiXws
bAjIVJtebcG6On4wqoTxSmU9Pf7cMOXxAXikho17n9AmOM0nBO2R+/iO2M0v1vmjyMHKkXmCK2DT
ipGkMbS8PQdRoB4hp9aljnqeDgMwTn/X4k7f4sM3CpLHmwPjvzYAQzR6I2VoqSgDP0AYjUp20biI
EC8fIqwilzSqAfAM981PmOWfBr+YE8woE/7AsN9chEbdMKKVTIGRu5nM2Tt2R/NMiHDQzfXprbOQ
fZ2br8iHWVRnIi02nRr9oaHncPw9xLssdmkZ/8fr8FrzeJHFUoLy+FYyJDF2gB0ITKrWxYd9YSTf
JeWCbYTc2yduTO8akyfuNekit4Ul9L6+6coU5cAUMiUwUjjVb0zsrhahqHPb+kEFELkWgvvaI7pZ
Mh5z49+kdiTiUcc3uZPpB094xnJOqaR+ghUl9houTeBlUQRBftITybHtl3bcXQmx4hA69j1wZaWi
T+6wHrt68Idmwsa6/PP6FIhjoMl6+noR2YaRIZbHAFkPmv8A0iMHuWfRYr7lQdjLtFNUB3yq5Bgs
ulhmSGCfCca/YX56raXcXnzmsFR+Hrfgpa41NTgGcgg3nlSpzd6wX+W5cFt+kp83gd/sW60AkzLm
5Y2h9lBNLpIb+55tEfuc0g+7P9bhLTq/rIml0ERWkOubqLO9ikGPAihlmw0VUOVOk366O/+qH4Yk
hi2E7ENAUif18bCs0lnGmEvv2nQ4Yy+CkRBbsGgLPXzB8oqzcVYCCDHURY/a+GKE88CC9YrI6KGg
I8h+22v8Mt02sPVncRWmCU3ApKnsJcw2grFzcA7BVbtYHDNVT8DbzpzUptLzZH9qCBO1zDSdh642
GGgseapmsRFkpj3Q0aKbmebY9yJRhAnxTwX2EkUnLktDaCH0PqF36mMif2dloaD7zf54U2kKLvG6
FX3eDJC4qoEsqGPR1PllTAQdg9zkPsjIkS2FfVKBNYqA53NPI/fHeMWR3UAdI2PhWiKwRVIJo1Rm
nWGW+6yRAzgCgAnMIOD/HcBvram3n4xE+RX3AuGDcDBmKF+Slz/17yr8phKgjjQ/r9WeZmw0XevR
aHTr/1Lj6K8BW6E4eyf0mr5LoO1riC8bKswHKlrCbsMTMPHBHvIUoRWEp7ySq78LNI1ESrtbN8aF
2TKaUCK1aMX0OJ36y4wbBE4GQFAoGmwAjo+YMKw22u7BHUb9nslhnra0AaQigbM1QnihPw7xoqfl
Llwx8PatF3GEX77oGJjPWTggzFMcOzKgHybwx/R00mIyR1c3Zy8svLyEgR/F/vZ4yfpwFKnbD8B+
N3QYybjDF+m74K1xl4/NkqpU0g1Wguu1lcLnKCK7Ou5qger1pO6up7jZXkbWSTjdN/DXoWAs/Rwz
3br6I4Umwys4PKJnPDPWy7mY5A8ka16i8aUclqhkI0pHh4zZOsgLTN+JozPNbgMdOkVzTDu0f/E2
zzlfpQQSuZpsaHF6NfhxWxzgJXK/NJtdoKjnByDGCqwI/Jci4Z6t4HBIWjXOw0EabtDJ58G5vECG
/y5q1r41rUOy8EeNdJif+7n1w6aTiRIiN54j9t6AwiVidCZDxG1lqPoVd9qsPzcghVDaYre+DS0u
AdiR+CsikVfdjPfCpnflhimjUcCXuE3BtuSvPXYn3nS1D1i6Pjr9qAJCNURLkH2/ESso4OpWw5pO
ZGJQnuvqrQ/GCKXbGEHjXArDXRKed6/6Gbv9uynnHaARnlKUDFmfl7KWh6BkKX0+fVIDumlpqaob
IWZr6DPho3zUmRRaLPz8COfkPOuFmmc916KMTMUehTerdgys3uqtQ/pi1ZClUU7GPVjr7v9ovPty
q6geM5+8fRCFaPt53k96TIyMf52X0NqS/b/0xzd4BC2V0u+8dSblwoAjo3ZhdLcVskirrWyB8lMc
m/qILNaxsg7bc+CKOsBVY0g+gA9tSg9AYLptwExGdvKMh6xX10l0i2gY0RZR+4OsTmFf/tiFYDnx
yxL0c8kXLJqtTbDvVagW4xwYmzlJV1GhODKNoYrjD93KbSjT8RRA5BWPngCK5b+hZv2n1vR++m5V
xHbp3QHif+Q0hFGbkUoiMV9f47Dl3QAoIvVe1hGHOGOMI6f568WbTvSB8ele/SAzAB6mpArXSVRP
d6TOkXRkKXIOyScMgFIOjkPsMFVljD/XUnumUgvq9FtG0ZkUapMs7hzAOm8JMdW7NLA1V+B4E/W7
lJSIsV6dVAbIyEmu7Yf8NbEvY7nTS7yNinj3WKn6tiFDHk6T7SNykYRGAkmbZIMsCWdKypNWHuQB
8YtNjHwH38pCHDOA+8JGZz6Sbk8NR1etGUq/EoBrTvNbHCbFbEIUnEO7q53jcPxChpRUNxbr1uJk
AKEs8mKrt4IbcOOMSklLvKkWE/SlP4sJvGO/ZtCE19m4R/fd+vDDAboo+z8gO3mrXhHAYDoX5i1W
fHF81icBG3C3Y77/qxsG7+vW20dFo8Cxa2E1XloM4x5uQKtuTxXgBYQ4qHR3eRXwMEGQXiOB6wYo
QUybBuLax3lH2owXkHPx0qnm1xlKQ+pzmMLKRzbZLpYNfDHQ6aZZYdDCB1NVeMonflIcYorqoOld
0h8EDO8kyHW0OpQ3A9W3elrh/bYmJ6IOHI19i/4pzpXAtLykUlJcd8skildBYeQ/MK5Zh/xFNzOS
QJTr4gC22ADekGS4b0px5gY0FNHVCEg3YUUxexK/KYQcWw2b8yk0lS7/rXu3p+f6JkchOyh/AQ94
4teNiZP2YnLzEdMIPOWySILN1XAakeUciXzhhtaPAEGIXHIZNGnvSz6yMUZk+d85r5hqCMmvWLo+
/67aHLs4hc1VK/2xsWF/T2GJcXXQS9o/Le9wClUfS6+kfk0dlou3iY4jmYdDrTwwlJhJr+o5yNPX
N4EpdyI5140nOCVR6X4yHqTbC/V6cafJHOQGC1wk3yxWfo/BPiQhM+rfp2a/qt7wCxxg28LIeW0f
FKySayD8UMhCkdtFPI6ycIxA1izH1dofsqsoF7AGlH/XMu08HukjIEp/V2hYrfLFoIsdcZIt+lnU
RFbNFK3KaNg+5d9y2/1kmhrs/+7qitIOdYrJVtku1XesOlJbXiM/9X4OSQ38eWd2Fml1yv9Wc9/W
XZ0D+umyyPxGutz2BeJAHts3oYdg3SFxojqDQQHZuKaZPhJ9BDXBuA4qo/ugGwoe7C5LfACb7uie
McwQ8BIzLm5xJT7sHe2Dn9WmVQutRV3ZVHmWaBHPTb5CYzsbzA8oAGCcxoJCCaaKGtbVMAv2RzCb
nzPoIvchQtNkBY6nuzep+S1RxOkwGMNxWV+u+kQB49Y3v+h/i1PbDH/DSUtIqDZgnFnthKD4A3pT
M3f0nRvUEZbmV1LTH6GTrERqmnUJUEH2uNcn5w4rQZAWS9Najwh+UJu4ntDMq+n/JkP2nVVF3H2E
yZogS4pDeHGB/u63XV/LP7EfEZIwVt9IZwQvVUut9S3llI/hlBtxiUtjuvesCVzXt4RgU1Vz1wnV
sI1zs080PndLcF7mdIm5Ri7LTY+pLS2LLj6VLZ4Eo81R5dfTliil82E7vIVBANDoYpsagLMGbMn3
WMVAR+8MRqILIxVFyf+EGnlag+W+9wBHHEFIpoXsr68mjDWFra2OulqL65s/uF7MrnxWclHKAyEB
U7NJFDyk+DQ2yeDCSstDGmQxTGzcdmdwBRj9g0iVgUGYazPyU3RLyIsQ9d6WAIpugrKvA7FzerFD
xZoKc039QwW13eAt30QhRH9KDz4aZOk7isDOMXL5zMwjsuNSkAnxWaYoqBu4LpMgDPGTpxUwcz7z
F1rtibHGp+xaGPg/9RewYM39fbIeJXBfQ89u29GUmI5kVrKc50yn+eb9idvR8pEA3M2Y7KBjxLcZ
4XW8pGjPcJV5RVyCsy1Q1O6bck8NJKy7PnTN2lJQ2n7rXHbKIErBpEqwIKAVPOAxjO0VrwO25pwA
NqXSWBgUmMLjV0h+TYoG/QOv6DxeCLUhbkxSaZdcvutfdjA7mfdxTYpktcpNVbVhQOLPimP9uVcw
3v9b8YgQNdfN5L2OC57HblrPlvFpgyp3iWvdVakzuTP+H90bmwqzJ+gJWEzMvc0pEGrF4V8iCeAI
bck5ZaWWWFlgbIgWMMbW6jEmDg6zLCB8o7su1x2giMbcHwtaEGubuxn7Ij9/qV3tFl1yOdTXAo2h
DF1Vik/4qSlnF7fLdpB/GzCU5bKRYtfSYRnIpVL17zvLYVnQuNqL9MaiormCQYb3tUtV9p8wDzOh
tuHU1qjf10cPsm899Mjw6/JDKJCARNXXhJs77R5quNHrAoWZHWjtf/D8WLy9WJRr3uY8040YO1lp
V3HtWO1t7fPQGeOHscjNIDzs5OMYukxERlfotj/GbBBTAB/687/jyu+1Ob0ytLtrSiC4nrnZeLc2
rw6fZVqe5JC1W4SP9i2N6LuIJv4GlRgIqN8fjHuZ2xtzASRXr7t612PtdwcUGBbCwHe5ANxo2fq8
HapYrFSnViYSXvlet5HnIgJBBGfM3Vdoe6lzxtM0ukDmlempOq6puZgga4bWqPTdpWDNFLjkp4m+
3iHtkz4hwAf/Is1J2YpIduV+yzgPeocHlkVuTcNTVYKJri6h2djSQIqfp2KKNAxNdi8UXADF/P68
8L8DHIVjUYPkO+RZHhpI0wRJIZmJ3uXEmEaaR8v1g2RbwZIzsU42wNLGNUWkTct62ixAk7qt8ZV0
LDfmh58SNf7eOz4K4gIZLqcbHBdB55o/FZETvlfgA4se/uCJ5ljMSc2VHThsNKZIho9o6VbXhRiQ
XkyR6+pp2huiHfk7q++SsyRts+l6/bpuFDtGIAgJFYFVM2cIXJkYUGT4aeqC+XlEHvUiw0rKq0rj
4xJk/IvPcm2GQdymam06wjvwZBF2yXmc7z7pnJYvIrwc06VBeLrGQO8RkNSfoQYEse3BySyjpGbm
PkvIxCwcH/OUxvONKAVMircwmA4NW1Jl62zykdPF9GUiWu0U7u6s4cE/lsqmHFKMH4zb2eVIAgx4
1M85GR7bBDxtuvtjspU2d1Vp6jKrWdGVtoMX0ZRN9/Kd/NJssOobURDfp3hHsiFkLhtTd3XJNi0k
uzZr/Xaj75FtJbx67fIfn+Ii2ZEz4zGV8c/64Xw+F8zJDihvvROtIPOBS5kxALDmD50AShNl9/VC
IILatQkSyujtQBM1VcMVOzTj1XrPJx8xgKjVumNc20z+iryb6RCsXPOZSUZ4Gv+WcNi8EQgQvFWH
CQO6Bi8KOa8Tgtlapa4X9HuXKAcGS7GJuZAjzTjkD6UOGZnEzawnT9NQ7pZxNmKMS4iPSmwiHmZI
g3kC8MHFj0N8x+aNlomuS4SAHHw9R5lvhJvkx19kdm5PsYzWpBlxogATl2J9WPNX6mejV0jCcsBF
mzKGoOa6eOdbXSeM5GlEq75anxo8HR22IF9JPVz9pXJeSbS/gYgeHSKbSQOuGtKbJc0TuaVxwJT7
dwrJm27LzQ0hwG2pfHsB+EjiPoXN8u49rz3rFqQ/8ePk90PxkaNwMGBaCKRCCiDuqS6p3NPmAijQ
N91KtTNdheMT9lzWjAjA4hOXLreSz9mUPewGBscXo8CSIu7nnD6RTd4w7Zop3zDNhSnZG98RjaBM
2i29nvqar2KuSUGhCkmC39V9iIMdm/fqS4npsyYnJedl9k6hALQdo0c0/naVxNAJINao8tuT/jGd
3EXn9nW6o8+hilrMQcTSxfqFcxJqQa+T3kVTKbOZ0Uo20DOqszgegcu4HXrSJxQ5QcnJIM7W2dsY
VwdjR0LuQA22Lns7A4+88G5viHdiHKe+UZ0E6FOGNRWgvtL71Uk/3nmbRO0odOcIpCLpIXvZRBU9
MM9AY9IHaq6wND1V0QdP2ozW78vurQwXVILxIRI/pvbXFFEFysUOrImXCGZJKFGEGGY9QBW81x95
7k+HdV4wCBLqkDnI9eRGmvllToAPj9opcnp0zf3i+pbt/Uw35K10yBLMFpw+Vcguu0x5oxGU0Q4b
kTKAwRHt0avqYiVH2Ny70sSE2SorrBJurQIEz/kmHnwh3siwHA3xE46eCE+7fcvWWgApw7+kYnd7
9DmPB1sCimerLbgzUMK/V6vKLNBllWD4/bJaD5wd1WHDGA8RECtu7zVs6GHZDJAtb+rO6mHSZeSr
maW8HImRqBDha41fP5UbzpX12re//s8GEV3llAzeE3EX5U1ed1KyTHTyXwZXjCWJ3cEFdyEbJ+1E
dsjuEtxq+RsKFiSVcoaV5Td4n0JujQXPwUMQlENFEdlWpwgaud42C1V4dsp/NEkz3lGvs7CS/87r
AYJ3kOsGh1fpTH6yna1i/QR12SQF1mPUGf5CdNPRizspMjgHttspEInFthLRSR3dAqoaPwCi28X4
lMS0RdYqFSPCO+WR/WYYFvHyRxNvUHkTtAFhmCxoR9IJVwsc7Kz0+Bdmn5Q/txSlR2KEe6SWtm2n
JhzSZZ6eMDI1e4YL09CsjXcGRqIprPbAvZd8zNnm1RheBKMQwTCFvUwmRpfFPZ9577vM/aB/EZak
mZLZngGcMoCwBHX0OH7Kd+6G0qovQ3khBGXiTnFvGqJDOaN/k33z9ze48UmXb8uxrSuc3ju8OLQB
JIaYEjriMSA6xDlVaN5dAgkNqObMY7zMnTJzB+OYvae9syiYLcsHtC95y3C5HJF4dgtgLdk2+rUj
BYT8SQ5DXwRuhtZJ8Vxtqo9tYyBp1ZMWFl9LK4PNygpoCE+l/T8ZuZ/YRKxNktDjBbhu0Dlnkyo4
75goqUpbQo5ss9sl3e/PGllq2rRIhqYQzi6to2r24h6aWNB2naIT+ibR1pDF0RtyQBZF81MgyFnn
/fZNXXeuPpQulLWdhYIkGPKPHEjyLoWuAd2vz8ZJ8aXIdEDX4wmpAtU8JEw+IKlW+idmmgzPUL9m
4X8Lx3t/hvxSVDOovN7AXItKwDaUKkMFeaCWgvSqafrykVUk6EO71XO9BKKGcIfftEd+q9YcvMLK
t8iScqxnrkcwISDn78OjeHFIoaTrAUg2kQFcKKpWSOr/VfXOYIK1ulLdJN0CYla30Q+7ZcwmWo4C
Hu/8lEDYr+MtBN8X51bXg9/p9KFtajAq7jC36N8W+EcZy16WtIXsNtQWZ0zz/sN4+xeGrgQPPNop
Ltt9dzadduGm0rciiyPNIHqayeewvJsfUxdve6NR0gsYmwgHTozdMxBK3ewtOrL7Jh8TLfj3xita
nudYcSmqX8j75q0aDG+wXYi2D3tGvCI84GN1QrNgPR4Qix5QwVLD7ufTGxxmRHoO9hrsl0VEh3jA
JbDsqWRy0LPKzUZ5a4nAsZ50/KTuI9pAoW1THfDMi1bB5YVKrI551MpIfmiwwQDmwHgzh7396wvR
nAQqRwixQLv2xgA2VyQEaJq4WvhN/Pq82sYsA3vR21dVFRrECbdD8KMZA+I3u1OkSNOF1MDvaYqS
3Vmb+ZxdWANmWo+OZvz5U1xCtgCLj1ei+MoYNEZdKFLRAMQATKHvPPN12FHw5DuP83v3l4FZvdIW
xFrzRhCQ6aDRsr2NV58WBeZRI5a8y0kjRgrHi0SP3QlZJBae9nBgrs5HxUxLD3J2COCoCb6yj/rR
/Cc8teJRf5Cee/SKNZ9dXadmcHpwKeXL9rEM/X5lTC2cI/ZtPpNaUUe3lpDKNFGatRDzKXQwzPId
BffYcdFJ1M/rzKkRw132FLhEtyEHVS+UCBvMcagmyOGoudCrLe8vWHBmXlbtoRtKN47sUcclZC9z
+d/Ogaqpsp7oRHcPQOW6Yf7yaJKbcaz0B9YBzOLC1jWRGv4nYEJ9VLYhjUqA1p/QQsYW1UAwev7J
5blmmu8pgzOJHBoEHsXFNo6olY36I8IUSk1dev+C/TvKGKo9LRDeJ+Vpp8TikvmKpthY1+8ctFaj
S7Px/8edCAR9h2LBn6T0GKPLf/j/KQrUHQ8CEeabZCzBGXn+TdRccEtFvYaEfZnsHACay8r7G1b0
PcaZaHkzgoBhczCq0P5JQbptTp6nj0cKjOzC10HbLWLPXsU39wO7q5g4iqOidCYU7aJDEBYPXrvT
FOt8RDKzqDz5XAIZeLKivWLRYIJ0G2Yqz9KcADsKdveSXlMVDNmS/YkPj7X+uIQxVuBYJBMihB4+
U6ki423yiO9fZigZR6a+WLjs+ttiIr1aWzLUXca1iwsgnE+kFyboYlhjS4SQDj02+qhf23wJauh9
yJxOBjITOJS73wI4+szrp1EWHHeIkOfOrAlNEdi6sGH62nHcWwFlE/2B6WiuJPwSWFJx11O/qaI0
yHhzV8GdzeXBZLXjgPALG6iGzr4XESjr9wgkYigj/cSlQlTsSR8AayBE4Dyo9QUHrS0Icov48F87
8uK+LkwbpSE9X9qUR3p+UJovODs/enObrQ6xAkvY9XxrDH2QdAK0qV0nRa5dZ/j2hQva0ZTPlQVZ
UBMq/pvs7YWd+k4+xWGQSDVaFVQLBmx3FqpfjIA4y9VmW2ONTQ22xEXgvCULf1zWI1k0G16SHDIC
CjcW7lPyhzPRpzhrRw7MJ6r2Zk1j2v2L8or21Ys53lZMm1K2zQYUI3Km7hBomuxCGNhhOdbpcPNF
RRtuRzZQorEKI7PnABjND3U0W29ikuFgfCHXzhGj3V3/U/kfMYiUEGbet/V3/DhZwIBy5yQSEp9G
U++ZSpzg9Oq1u/hIFoVy9DCb0LTw5uIZYtPe5i8fPi9wiFryfFNz6daXxc+V1TioI3o+jhKRSp9I
wbB41tVT6Je1vjJ6x8go1Ip0JpeNcIBwJ/3Y4Ab5Eph0zHX7KFHDWCBD0OOB/5nCzuSL7ku6ujN6
0dIab1o8fIGOQuT8k8Rl4td5vW/f3u/TwN+ql5nahO/r3XWQwP5nP3l1DI9KDs8Wq1wteaVBQp2j
ARZdQEDEPwQanpqcPRpvzsmJzWGAvxM+9HxJC7/loxSpmsmA6ApBVVOAoJll8QjEnEfBuDChnQj1
hTKtQ8zLH61E1mlkTqzg9LelxViyJc20zDmodPFoNQ+6jyCJNGAAldOXQ4VldHlaet7exy7pCUyv
UNlgkYJ+ww47wVtNKPYCxNS3rZ1z09w4tuYmkzrW7mZ6sjsfMU0cU5TRVbv5Nvxl4qcasj248tiP
NWLgcnFLpQWGIKnBAW1XUAKwmdqlnE78VxyUow8cTZA4kDGmfT5rtjsDRBRl8oSnMhd850rYqC2y
JktRgjlGdFFCMqHH0f3WflKWYekWMpvJUS//glM61pLvb77h9A+pYjYtxAPB2XsRNrooaD6fA4Cw
KuxrXEp1b50n9tJKlUV97SS29ab9noMLnJP1gTJ/4p2OrnNilMOFHfsNJqOqn3dprhV3srxg2Bte
ADbUCqekDoyR0rmS6lS5w0/QTzMosdhFlSsn3aRAr/kvwUdOt7MpeEeHmdSVh1A6G0TITwVm62EV
cwRwfJ2W97lSs1gyFUorqmyakhrr5uo8RdUW0HiLndS/SK9B0PQ+S1GFNIxeWM2tegqrYu2x0AzO
ZgIl5jgs2eytLQTF9FuI50N4r3SdO6Nr6uZhphCQwBhCcCyINiIe8CNEU53xEQXjXWuZ4C/jVmNY
nzq5lT3GHac7Wc+HN0294pxiq4KQaF5NaXN81zszhtiEvfa+qvK8MD984dsreyNbNs797teUSshd
M7LcMMz9WSkzTIwXui0e9B6aziOVR8wHQ+3gO9zlArX1L5oNte7tVIw4WUcWKxSAf4tN6zrrK/9r
3Nj3QuILaCewHfHJ9F2ePzPF2VBgnVabUvNj9BJRjvqL2EiBYogoUd0SbFKRMaO4Nrasj3zvUK6u
8fKnt1l8OQhGKMz9c9m62qQ81zqC0jcmPtj1PcxL8XthHi+NNtoCh7cMix3CS2SbeFvYdLGnX53M
P1fmtFYs3A8Q7CY8gaagaZIpWhRLqxQYl4zR6kZLrXoKXNCDRi+4JzMcgMts5IdmBxg4egs7KfNU
XuQT/v7vT+8Yq1KsshfnvKWIVtiEOjhK9F/pLO66cQa7ZZriOzUeR/qdBA4T7zyJCWGfHZO1CZQ5
gG054XGFG8ybRzk0fhLxg6elApskfo5VaYmwZtB4h+8vTqXmOxC8n1tM8I8osfztYvmhPQd1djIe
OTLKE420057DRWQkDSFgd+We8IW/EApiBBfx0beQmWNR4HXLlTO25aCEzFDUfJC5qRBvJy5If9HW
8KuR1FRaR/p96BY880sysB6mjbeYjNWn7pM4miZXYJHlDaFJVN3Uq+KyzIC0J13iVhbnPL4=
`protect end_protected

