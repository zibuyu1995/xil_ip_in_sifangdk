

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DKaw2YF5X/sI0l9aLdTgbK/M5GUdtEMTnIFmxvSMohXCNpaRunL9ipaA59Dc71YrenIGtec5QT4M
zCoGKmFbyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QRHRuF+/6jbJdc98CuDuU1RSPkw4Mrd2rWInSv90clZq9I1OTAA5/xdv3Hk99Vg2prXDV3YjNqoB
pcpnTJxql+YZ6VAzN0qCk+oUeO1cCu3qiinofcBjVXCdgYxomUKUeE7FJeYz3Js2G/kJGoeHFW9U
+zAl6jadwyF9Jbvv+i4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lb7wQIOJLuT7MorOQ8eHbXO7nLYJ4w6DRb/CRc0KXgD29tV/pKu8nH2e+iVICJbGwJJtQ3k8P1j/
LscOU8Hk23tTbvsi/KP4jYIAhUNpSlUfm6H0KJ2yht05tm7/nGOSq+YwUD5ni46LH6TZmw9wRjLo
RAHSpBohLboc3y/hVTXta9kQmKPnqAmdZWZqkVyyS5o93+63/fdqbFaxxtwx1mXeZDQ2+2zbTCKf
tbrO065IQsNhLqpQ6GmWS0y4Yk762FiY/PW8xLoCZ1V1Fh8ocFk7LKyATUlQjo3T4vsNks0JLfh6
k4wW0gpjLf86zBHim396ye0D0jCoECOhPpGtaQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZXacKhqAwgw8zLrWO0Oej9oQ1uNqsfSW24Ju9AdSqiO9hJgeX3QSs/Auka01BXmxZF02hREfAK/G
6uXtwOuytUDW3C0vu69znjuzfKa65iqAvitXfuV2wV2SBDUohxstI576S9cHfGPfoJ7tVzjIg2t8
+fXxMYGWVW/hL5Dt3LeBc+ul5BEG9/vwugVmMP2uMG9nGEtDEQeLb7bWAsdsP6jyz5L4K49swiWc
6TrDCW/53r7o1y18s7qcumMrH+8e09lZWlV7gV/qSGCmNFjNoXkvbq7X5+RT29nF6kaEY/1Y1wcM
sqDv/0rI3Yh5PZatD+o2YnHnz7Es16C87EBZrw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pkb010SLYsAhKXcWm+QlAA9Be33Kx3pWG3KQ8c4OXZxiNI+ziOzdNGDZkUALVJhYeeODAczIsICK
xPobg5BZJdmnFjXMkYzJiVNc7H8OtQ+xwCOlZfGQy0nG30bs3aCt+0ciZZz0ed8EJ3QfOUNUrA8S
ACDctQvzk535zqal7JGqVOcbax0rksASegZXl9TYHMAWSFXsQNDtHG7HCq8QaEGySiiJnEz1Zygi
CXmAaOXrSZ/75eRU/jV0Zmfl2uX9M3RD4WyT2L0mtTPVI1Jo5riNKDciMqi09G5yCgGBizlVK0Le
ynsKW0Fvo5j+TrmGuES2+DcsvwzxQUmrQ9n9YA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
saU9xQVocYCNVhmm+/jaIKt7f7lGDiBCwD7GUeN8jk+fV3dDx7VH8BXnwqh3bO2UtgQTq4TYazR5
PsEJU9lk5Y+2uIztywixaUOcY0t6PGvi6DZ5S1UapcNaqz1GzVDJNMdFrGWeodfXgyVpIeng6Jtk
EKceFNW0p1SgbLjlCjU=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pbTosJ4LwLIDFDsIbDQWyryoCwFpua23V6z9HaJa95eQ/VgCaYwQRc0pJmp/UgRFI8GxRIcCfLjR
nDQiDTQUzYsgXuFi39wSqyum1ybk+zJc/c0tfa3zo7fAh7WEKBR6EfegxJoOfQ6umn8yMUOq35ku
5cQGVgAH0mV2j7kgcszzSTcMNu1shLKlPJejpCdXAsAct77F4/JiYgr35R62Nw5TiOPHxLGWKlD0
S4rOzGqDzYI4jb5eYbnrBMtpHWXse9ybFZPj47SvpsioKcFIHeUE7GrNOvNDQPdNPahScNll6gSb
fa6tuXH+3Q3DQNGg7RW23POGEp2w+WE6Kef4qQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
t9Sis5cp99vYxQK42Ey+0XFUhT2P9ZaNWUAXXt227i/7C1VUJn0rLZ38mR18Y3qSDVZIniCqCZaE
bFCkP/UM+LjG/biNqwKYKDJt6W821gqcAEl89+tpOBwXrHJ7gnW5p48qM5XuK3QqzOgnY9Fucgtq
VbkHQJ/+TM2ZYSRvAwIv/duTuhq9nKnQD7Yx4+GKaG3Lq5EsC+/oyMqiTPhEvjgRpwDMlyDZaKfb
1N76Zv+eQFK1b38nrrAYbe7WA+YuUcO4poZf9R6dEqmezOeGYgXg2U2EyTqgJpKDBqRpFP++hkmA
b6xYYsJP00yJJEsludMP4BYyR28zSmccpRKXNuAYLCP2SJQt9l3NgGstQ3+zlRYzKsC/cFd5Mjhf
f93AU5yxiVpCvCiZhlX4z0xhjvlK1HQJhB1OekLIYXKz+qjITkyva9FUzjMZzPf8H1hTLYqYmNJ2
4gNq8BCBBddDKe4uEpWQvJMZIGnqLjuzp/AvNyLfvpqdAD/fFdkBK4vPG7Kb4OdFmYvD70ZbnHE0
Ax8WQkBytmvyFMsj4KMiH1g26wTOfse/ClJIhT83d0wj+6yNWBwuXT5PZLQrXILkFYsQq8EEs1sW
e8SqXYZFR51AhxTG+5PY0VezxGr0AngorgQ7N3IrwssfEjdWHhd1igevycvmSzvYT/M4kdi+q1nQ
Mqtb8URM3lNPcqioOZCklotEexdn43kjQGB/O1qEYd9DwHhB6BDgcjIEdIIdyCvn+99VZRNWofFM
fiDV9yjAbLB5dD54xAJwur3+kXIdU7gjT80Pn5AEItcIZ69SwOCGCdF4qx/koyzBxA4tgSJwHa9Y
XqgBusocgwo1W224P+2RfO/u1TXkSsIY4qr1xxgKjMC7/qMg0U++byP5b6QzPQPr+9q9JFKqTSn8
deecJmc3O/P/MZ9wPuz0e0IioeewxaVGXX861lnmM16tEBSvkbFizYuXbV97EkKl0TyBluk/ZHrF
C4o7mqUmwHLbPT/CTHtKebkjyra0NkZzywWbCpeUjDPJDYPI581q8BbWtL84AgA1Q7TFSYJppz4J
nfyG0/XOquKLFAeHv+oPR/g6CnAzow+WoqqKpcVWY0EPFGRu3W1GeU1JOuUEj6zadbPX3u+zOoiE
vTJ9M9vKcFdFCBz79tme5HfkNhh6FqECXpREvELHU5Nr1OtcpDMfxkMwbFouSsTjmd57tOLnvvub
993Ly4efHtrpr7xWC/UkvhP498wpbBi3YhLNWAJSerZwKPQrs/buERF1mB8LoDNk3qxs32AYP5Wd
wLg8KKJ6O2DuNLjo2zMTa90w++TpunCgNCqRd5fMRh065PFUZcHeJvtb86l3rFf4sXzSfjJ9wvz9
jftKSsjGvUGmvpVUF9nrmo+92GLXVhMpznFzGAhGGnWUsvX8rOTWk5Fgc0W7G6qRPHZmvulO+ECd
l5rFoL2H5qopP9TusSafQBb8lmf3upGpD9IDsOTksXCXFjr2kgBWgLVtcPDjQjh6AVic5DnK06mm
glPnYwoMKhivkGGMSzRHVWcDNN1pKOyQCqLMkolVGrogKepIXNIDuBYX5dlgfddH/JweOlNh/gUt
LsZM3QI6u6l+e8L3F4xL94AYBKt7g70uHLPze4HVwlbtnmlb/7cyCKfeMesBscwrj+E5tFse1fQW
6XrzvMYGochPuznsJRJZBYb94qPDAHl0+hwAIjHB8UvnCwWBgw0TAQ/FSxEuKzbyRok4ZZwwShqG
/KhMMrG9z90Ot5TnBJaqwYaBTIRbVqovhXAyWJviFjVbvL/H4KtAXjQ9NYMQw2FzC+5+Lro9Quiy
CtkkCxNILAAnd5adbZzSFT4PLOrqT5nXio9WL/RPJsl4uXIp18Hf+OiWXpdBOVb4LtsoQM4mfHTf
Fpl6+0cxKiv+g7ElzqPvVxXrgsZNz8Jt+zOeL/TXNDaX6w31hbuzLFlCk81Dq5j0nsyHgL0CFVKN
Z1ivd6qpYle8K08bdK5goB2bxVKxzvACYZ1EZFPDNtxSx675cMl5U6A8CvO4ZYO2+S60Fn61k82Q
H7y7D591egHe8/2Jb+TaGMAKfi4cjVH4HjNqqPs9wtVeBMDkFwC05ACItauH2aJLHlMNh66jfSKz
9cCKCSiDRugAK06SjIFR7YQPLC0wnWKYzYOXAh0dVJt2a708nRX5hWd4PXFs5TU5RZyB3B5wo/0B
XqpoMaz6DNMAVd9CPj2v7SXAGNmDzpt/Td2siCDe6FsTyduCZd14+KEeSFBBKFgCjg67/o4N5UzZ
oTrxjgRy2O0kdn0C7c+r2V5SuouUZ3fcUIqcZ45zkDpYOLoMm9ccZKvFTssFI7uZbD0wAWEPXc4o
FZrc8citxRDXHr+4TxZmi8A3Qd8iUixK4r3bcHHuuzhvUhjDDIj+SGIbypBo+vQRtMd8kTEZVcmm
zPAk44e6536Lr2h7cU8MszBMWNQwZT2bMFsuShATP9+fs8Y6z4Njhk+xZoo4FOG5zZc2HG1BYrjK
6unyv39XJEo/xXyYCKc+cikJHR1AGhlZqzMuecvujyU+eo1hWnhTcE4C0jA9DgP0S/N7/viMIcPQ
C68ajDVI5D8zkO3OehjGy5tc4dZ7BAnvfPB0/0qwIqcHCRCntBIq00aI28/462X4lMli7l3osSN8
/oY9rd4pWF5gvyvd4G3+XG8pqtMUawUkcUj13lSmDOWDkT7evmaOYpHXwL1y8HILNIcGkcu2BR3d
nw4PIlkYdn+S5ow0WEPeoP3W3gKB2O6vdOjc2SslGQf6y39taTLIks1/Z+yiPOOJ/F8dzh0gl4xV
K6/OQJJcbrqOpD0KRefjcHby4ooQt7HRB8d19EeJ+fljHcyHSUZ3q3QsIA3Ei28q1cvgbq8rVeku
EvrL/HvA1K+t+O0RfiOJfjJMrV6AbD/GZKkSKyhsjLG/ZPT2rFhfxhz5y0FWNb9o4o9fmGXqjA0Q
ld7tSC87E73dHSldIPVZHj7ul/acI41mZPFqVlUH1MglBkUJpasOsXa0ErzMNhHd6pcLCnxitms/
yVxO+GgcviewjrnPuUnSeYd6wpntwpxzoLYByg10iVTEEuY8SVq67CU3jtFd8T4mLsfWCs7dtgNh
rn4ZEHhrYAsTYtwWzAyptz4avb/o2AvjkisAoVufDTnK13BRV9rUmz+bkD3BzBefaIaKj2ggTz1K
rVdszQIFfK0qknVFdtcy4uZkJXnGSLvoremkuMnuD6SykJbD1Iapaa/BByY98ICMmcUK+zIsGx2e
ww+e/LzbN3zA1Mlj5vZjDgQQwK5c9Or8gngKJhs1JlwNUML0vpjbmtv0gzUjpWPsLql/F0VyANAA
gBHCJA8El7msfGL4ebvJCp/GDc9jpG2j6TMVNOvvrU5yabqdtRgqZ1AWF/xthJdxy6o7sH4Ab5A9
wR6y24qmBz4vQB6ByqIx9rSH7xiJiaQia6iRzc1WQz8DLeWQy63tVoEtOZW00QZ/1Krt+XnAM8kw
buJn/NH1l2ePLAnPqJRR5ABN4bQZQ7NSZyZpa05RmhptFzViRSnzeId36tagW6cDV17SMkD75MnX
nhXX9swmQkjW+B1+xcb10ACLGafndqMCEvfy9pMtd0DAPtB4LGoy3+pi2QbXrSW9VPyBJQriGdcz
E3+1FXOSH4u3mcXx5DRJ4UeR3sxDVP2UaeVl9NA1RB3X6vEk6HKRt7tLGaradirr75ijkLL1P2Pl
DPm+AZWLPDO5VPPVtmLgvboAqXUS/ga68OZm0T+YOPV+N9rDIv2ZO6SR/ncdZUn34jBrgCfAvnBF
M6otTaTFwSTfvbmzNGYCIH0/Ob+pi7jWT6hnbWrHZPVV6SDPJ9oTwfHUzXFeH6RCi10ALX2kA/pk
aURJCptaQu5ZIvBkhNYhKYBwfE8TSzELpkhWH/kS8aw/78unfH4S9VnRzSInwIxJxIFUSpQOp1c2
PIdjdt+aIIZh0OYCwi1Ixv2WlE19HVSQtSbOIhfuw958lcoyQ6u+6tjtcoGneE0mMNO8XGVTWdrV
omaQX4TTHDO9ImVdPOLhp24t1Wy5KlDjHxUCXzFn560BQl01GWAJ9SCyATosvrzg7rbUmR1z3fhc
5T4I5nt4QIWutkyexWjiAy9C2VzwX+Bs8rsFbA+JbqjqQDYqkXnPwCdYpn2Px+gFzQk/J6TaKXC1
68dTiE/6vyEG/hG/lTYTX7O7Eo4W1Iglyn+++lI+zKdVCsgXnLQDYBqHa6jsFmsGqpNQMOQ2jlUm
Wt7sklFaW/78Qutc5jmkNyq7SaoulCzed+WPt/l/mC7PI9lNAJet3Lt3KVmLrcpL7ko53/scOUgr
Gg3jmhRNLBtr07utI4NgVRPec2m8gQCX2X7r+SyNzAnrzeQ7cgZYwBzNdcJQYF7bdLBAtICAZegL
7F2RHVpielRbDw0nvR/pDt/3aLAqpNq53Bf0X73wdzLP4KOcs6ZRn2Ns0Ow/igwWFmlDMbDLPH0p
TE89l81HzAkMZquBjkWC15x2UaV9agJPt09LqKXlAaPPHqchgp7qji9ml2lXnZESo4gotJPRcWfJ
XpAwEcYBY3Y6mmoYET2/FxWhkz4pEaVdPrFwuqd/J1HTbfOruXvxxd1Q4VSX3V5UfUIaZkeUpM9s
rJeStVRWUp7hq7MH7odRcpL5DzjxNgZSJY57thnEq1Pl0gjFG1HPTFdNcJ3Er/ONB362lWzvkVXE
2Net62NlbUPD/I7t2UVYW5JEy/dmK+WLGoXxHMCiZeopQ821rq217p//dMq2Xcou/t4V9KZg/TLN
w7NNwZTidQhSLawFpzVA3F8j8Di6MNybN7hjXPchAjT2ngOat5N62JqIBxs45h6M8CA0RJ7pIjdi
w3qXVUH6xwPHLEwqkVAdC+0Xu2e2/ES1vw7/pzgecgBDzYfbB49A5DhWN+yh0eESo9QmSWwm+5iY
Ih/UVtfetIqQs/5EQGohQG8/B5VaK6R3IwgpP+PvBkK4bWa6mKmFbuMlP8eBB+0hvF7A7kf/GinP
mE9o8xc11sQ1UOD7N+eNtJF8eQiUH9GTj7t2J2hXbZ+uGwJKqN5ZsKG622QnF7g3EHFeXnm08HOU
tUj/NOSujnXYdx01l7Gz0pbP9EQa9U/qY2cH9L8hNoyIKLT655MbbHauwysyuTTsO7KOJGRF8vxr
TamJ0zfk43xDOdcS8tANHf9ef5ITTWNLVz5tjrHioKbuZ881WNa8jLgh756bUSx8EFbCt7vV0M3w
fMGntIGvSr4Fqcnm2VoHDqGYF9bf2XP1aGuGvjPf9nRxDSvR2Na4Etzj61HzukZ8AXfEazOCQNdO
rM9TK6ibQAm5G8kcmtgNSQKlXCM5eFR6SbIsKfG6QrCG3zwnaYtSYhCSGInm0mS9ePEPupLkjPZs
Kh/EBM0V7sulZ2ZnMqbqTMWMkzhEUNz73h7rYsCLPIs6Hv59bsqlg5x5doaIKAxChosvoHSheq33
WzOiky3TwOuMq4zhGgVr/kXpCiDncpLshQQUqL4pC/9tK8z8cIkygJlCqajTCpLaqP5u1c5ktVD2
8i4/CIo5z+uN2oX2FzJ9L2gTN8FcAeSMAaJ0F2whnF60mgFHN/RJGWyNJWxJFKGAcHK4jTp3ET+C
7UoM73InH/5Lm8ns+pc6fhntsCwItqBKCLuKniZ59YDrtgLrOvV6QmwrQe6sB60urL0gxGIPEWrn
B2cut9nTlxUTOn0LOGWDHJ6GCh5iht5BkUbdzT9lb2ppWRzb8bGidCLfQ5jzE3jxzhUn69w+TgUk
16Eiv4xcEM7eDW3VdKM64wgd70M9AUw6/4DSbpU9auZc22B+qgzbNdMTkcCi6NtQoL06boFVNj77
dyEQ6dJbNfeX+q+QErYTVKpjN13uDjbbn9er9gYc50CfHCyOWHzRq8+0BXDei1sqiIqx6U9yeBKM
J8vZeop4kxFfZHK1aZ8pY1+BBVgBW15yV+kDhOQmmj+z3o2Sc63E2zMIuNj+LLArYj5weOtFK3oP
/0DJX23dL4gI8gb/yV7YryWncWcJEIbAhOkCUwPtMG2m+KsBF2xe9nGpz91Ph3IfTEHoO7j2b/wd
+P6P0NYMJnF7ngPk9cSHPDRUqERWnMSuIDhgu46U9txV4v0Z8w0MLhaqNOlv3qajT4xmLNq7vFd4
+9y5TcNuQGshOVP3EpErNOdRNf9h4L6lXiybC+B02EfPDr+yJgYFcQBS6yyrfeXyLubUU1A+d+FT
b6RkhcvXSYTq/WNxJ8abA8FDqg3AIl/vhz1AyJQhBw/OeDyx0+1N/yp6SGQuwJzofw9rlamrm3ax
JoKuNJM2KmeZrXF4n0aUDcH3vws+KBcqgqjxYyx0qnDtWRa8YgjDvynOmYQxhfatF9GqjUNgFCaT
vD3sSt0FJ3KefpGmS3JzMhXKEFw9dEJzuQXVZ8EHg2AlgNWFGFlB4bt7g/sDHy2mK4KdYpxQBqP2
hoeSw1ASQ+FoFFTd5r7/GuWuUYpezHSIUQcLAR4nvptszns/nB14XWCndH3c4e4e18T1eTHvGpuH
P8cLCcQu3k7cwYZ5F0bmW6Eq3r/0rfr2rPGeCIjhr/xB03MAbmI/xIe2H9WqG0nxATFVovXpdJax
JqTIHA8qOhTkS8WORAxIkuRVR5JWuvNQXnUAnbHsIYwnRG6R7sxVTPuL14iSaR54C0Keer4zDeTj
R1LUecA14IYAZ/QnavmtR6NmYLuENPJEj7mRhEeAPGO0IRU/x/CtvyNrAehJhVMtRS18hygttJfD
ebPWomxUYpm4awluIsKeZczVfl6LHNA3gvPQCAcH75Hgt+RO39ic9EoXTxFuWQ1Hr9dZ0YkNqfxh
SdVAvidNmykEcSQvLYZvD2Tgup6608WGp7ScsS1wENY3xCuOL3JUYqw/oio1nmGgJdSZUoAtCTIW
qoQAvS9eBl/RQKkCJUWB7JaD5PLvQX1hcbH2aVX7mwBFqmvoO0wriR0nnWocaeObWmtcF6tFUzgl
46i3S0NhqTXKj5zixT6J5HR/0VaeqriSbf9315RkglQ7ESvyDxtblfrM7uNOvzrFIMohQZqtIZZY
jgRAGs8S4q6G00YKtXXSSLWi18BYde1Vps7HTg7InvBnj65xRmRulUfZgRBcGuvbcfkIzKB+2AZQ
nGMVPNdRHCKv2Yiq0T/hTKUcVfk1hYC04qQZyWhxPyZU9YuWx6hOMgWjCXNmJPNXF2pfbRhydpl/
7VW979eGeCyFS9nfi6WqL49hVTcYWV0igkhjWVL6gg5MiLsACtMjpLuGf8iWygvzXMS/JTdWRK2w
tzuT+qeBvFY0TYR84+wfXc386FsjL66RpwBu/hg49uxOVjY2jAgqfNV2Xhl7xkKXoDLQOH56QVhe
nMH5WgtUo7EIhHl+Iqoa+s+t/z3n2CGtLdDeHZw+JY/yKQdzMLywb51MStvUhqq2yWoZv2tNvD3W
KUwrctDlTn8FR3QH4VJNAQSyjHK/9WHq+q1aXowx6d2kntHwK8+i8vj4o+KpSvREbxTitbCzysOY
BKuolDiU+QQBPmNREFVxE63ez3Ljw/+WwIGqxtNO532Ax68uqx/vWXf/ytgi7G9UxXuACWaVxy2r
l/ZiC167pfRqqT5v49G9h1JoXDm/6OFudyYOyQ91sf8SI2UW1SuRIh6j+WaqmIU9edKVHvdy7qgv
amn4DYFB8DWa5Y0w1oBJBOe6BlMwpkK2qicJFV634xEp451W0k8YYdkyra/tLOBrDAzpA5pyjuTp
1noxiCGbkf/fELN0VDJKDYAcM1z1Dd5bTaodhKKTvRo/Osh93TDSVNrVOvtn2j/mucRt1MJRPeT4
7B7EDczbSUf9M5VIfZG5e+vvQE3FAvwCoF5USGTyrZabLJaVlFFYiNgPSM3lFbwfOeyABimVjkQZ
Nd24JX2+rsSuMl3DFgO/6FhnVOOwst5QLBccz4ZcTar85fLfHFFBdNvSIabFk49osbtAeo0hNjKT
afmy53asZ95T6/dyUAfPc8UUiqqC+5p1ctYU0mqdRNV2HHtit9NpbmrdroEJIX8OOo8kImsySDrt
jKcn8RNe2qrTzD/W0oKeKa7+HzmRg7/qTK9feNeck359HuDekv0hWmjI9dFkwfrpD1w+qrRQQqKi
cv5E5NzANvsCPdgqnzho3AdsbsAmWjRbzLLHxbBzeb9gI4WdQE/GFjYm2h7MugsEzl6c4R4cUf99
8+kH5sZ6rK7Fsej1KDgYIqWMuBeFK6BR0Vi5EeNBi4ilEz9OQ5OudmN8qY6k5RFA0zIfua33eUkO
qYFmbc5LzsSoDT2B65N1yl2U/zIhYTDGOgPU/PTXet7hGOHe/k/apso9JcUVflVoW8x4vLiIxM1/
nlgdQEGGclG3EbUE787epRnmezZkdV0aq6TPrVOI3RfpfJ3sG8QLwivVesLx+zjf1P2HWVXgKwRN
py8orWMZVfVSCJPtv7AF7WoF9HhVIZe62pt1r6sJijjlhHrUy1t1bbCTrM3168uBIl4FtLQLMU5b
nRyvdlA5r45Y9bPXZuufPeq5a8kzHJ4vC+QmQTZlfk9Thuqia3TapzUW83kLXTEkgmr9i5UCTqt0
VGTAfEzURmm+nkczRi9dRyWumPDBctNhNvGuhg4Uf+OxfEeBnW/LpvS7LLzO9nyexkH9rFLNsN7h
+GebXlWxDG/K1BiqsHsG8UWuDuupPDnp2WRVarnyHPmGkOkjZdo9nK9rDk9Oqc5xt3/DTIe3uYIh
TB5jU1aDOSrcdw/acmsioDoOjoR9qSyw2DxvYtaR5stZrim1fr5M/xf/5gPnEjTeOfT1hcUR83ID
bEZz8bBtHEaycl/IP8wQbdvKhSm9xDZUR7IwxihPdUod9AXUmhgTqfEmz8/r96nshaHON0XWWRfI
B9aYbzqIGAGheFapLO8gsquoaciaJOF+4BD7KkO05P/YrAv5+81mBV29u6PLVtWDt1JbUmKCy26Y
UWh8rbMh2udGd/UoRaVuDzBzZncHCK4CUTBW5UF+9p3XDaI1mcEffL+S034wTOP5FkuYuacS0KG4
WUnXgt1wJfdElNTn9VeDCrnMN5lsykoMP7e3kpMW1ktpOOOHhgu3jGEwXVXztOv9i/c68b/qlmwK
Yj7Uqd2S1FBKvRC4pQYxF5fb0UUJEW9iCVO3m7+0nh/B4L7pSt5dZqlJciqBpMXWQziJ5DqXjmDg
pC0DF81J26R84yKf3DkldLcJru7nmdpKytdxIdZsFuv9AlnO5eMtgYwnWTthhmKBgkVjaE0A9VmL
eQJ4eYn1vsIOufsp+VsIqJ2V0gqrkTrlbSlWdnv9pii2BaNOR4Cp3Pu+YYCbI8+iRfWoVhYGXgeo
JXtOAbRIQ0RXjdZ3QmKCR/BE8vtjA+rjoTJLabXWzxMaa4qwGeXkO1EMd9/pPf7UEVqQPfloK0YT
QLm6oq+buloVHI0FeOezQGEgoqjq5ipEzQHUbdUBysLSqkDOW21aQx/3yIHclFn6iTNJ4NSQU9vz
Taycp1+RZSp0B4253dJRf+GAs5or5wxKgwQjCqtaPwjxX8Ts+VN1NphCh+m8EnONoYMn2cqu/UMp
3G+8Oa5DpVs0ANEWh6lWyCEj1EvXKxmfI5uai/dEJywxvS5iTImnVGRtV37mWCQw60JkXbTOr7qu
7YyU882p8fJEObE7cA2sSDjwmmYr1l4xz8EswKkbAY5RmwqHgL7dULGjfw7hfduFbF9k3DRF8BpX
JXmdF0mIvFLTzMi/u9n4BK6VE69D5MguUvgwtgc7LuT4Hq3Py8Z+Kx6LzlNQGhgaSMfSkGB5+HO6
hpxa4fQvxot+52UxeU92OCsX08zYkw+CEAiMpaYJ0F/gpWNV/289iN0Qid2zFdjlCb8URIHpZ/nH
BTmAL5Y7zpNDf5XkejP2b2LBgwVFiEA6W9ftsVj4x/EE5WPA9m0TiHhnfciCsTs2mm8fTSI8D3mi
jW1ff0y3Wq3nTrmb42IrapTWWNGz+BJQlgFmURh7gHAZAECH7SWPFJVBa594i8OBulMtjBDB6KEo
uEclUX6f1Z5Zo8gJDMdXDz+pPLZdqijM1Y9g2WCogNoy45+nPLWno6oP1k0+aCVlyRmSP23q13I6
GIvPr+m5yjFHiKg92c28Erb9AHVPiaqfzYJnMtLHuYbaxAiOLCZnAIwMLl4gQVBPy8oG6hR8Xv2u
13PbiMSuJv0Dc6gG6oJvGcWBcyO3ea1zhKavKD5jy6xXYXUi37127kJOfsiCjlCjwCjFC1y1kCbq
ecfitxFwYaGzhg/KlR7+mrYUH42yHmrJunjxR2CruyFVkTxhrse5gC68dm83xSpc1kK9ghBWtuzt
gkFLb5ZL6qxXax7Z4+uq1cX40AyuCKNDkveK/SMro/0JMXUPmjieBYvmBjn4eRmtLweB90QWUxYp
WQpHE6l0EOwMarn4Hm1XRURXoHR7FipomAcJ04LlEcDSXlmWBsl8dGv44aBS7nX4vS8Jzs+7xdT+
cC7035iCVyI/0PDdyatmepW26CUAA/w/W2akDGy8PA0eYs3JoC0/IZ8vy2w2l0ftF82L8d6nrbrA
yKJc5PaLKEfKAbLz5wmU/izsz+uAU5xCYo9M0W5b4mo4jrwrkDYazbGBKn/1kry4u6CmgIlvz15V
dh0pERar8L79EpPMEut8N+XFpsRTjXFmkG7cUA/A0ElaKS+STCf6tUDUQY/crFjwgKiJJuNB060a
gmmaf9Q7JT6RTl7tp+JPhJMN9d596Zk631L3s48EZuEpeZsCk2c9zQeBZJiTiYpGDJ3sLNOOHcTT
9VlC87+Wb1v5YRDzrETtwMZHrWfjP1VHPdIm9abHp5xVIUM3UrbziQILDC3qXNTsm0qutsLnIaKD
iNRVEXTwTGtIzw9HyrMCJpp21yu2HncN5tdlwq6wZ742yizWmrLRyZHDZOEOC0LRFMP1x8NDcRhb
lczNmAVjo6gMf6n5ONW1oEmHglXyaUX+6qRDOMgl9HJHbofjP6ukUxiUfM4F0MvE2cPGarnPWUGM
KcUnwcERRwR8e9nu5OLw+0ojXtxs2wQ3gJ+v+jXmRdcuyKr4zUdz+lfyct/MzxVjPBKhWLe0PQpj
YVi7VIn2XKwXAVMqYFUw8tGm7gA/sWac51n7JSUybuDZ4p793iTeSEO/ZWcsfbecRfRsULC2ERJx
07MGCVDuVWs+PnBx7rv752Y82Q4jgm2ctRT9SfwhOWhT83hHufqMQd44W+KQEO3PmNcTHQtfHeZO
vYOrPs+rizcN06LJQyDuITArqfb4kRRi8IdgcibZpiElNQ1lQtZMUR8xWDyYztV87N7DSsrZkm3V
2DxMA1t1egAyowDWiHxNNUQFnTaBujQ5qCHjIg1BoEjRvydc+sAd1Tb29K6uDtRKh82If6Uwwy0l
kkPiaZ2fYc5dvzQDj0ggO6zRVZERf9kw3JjpavTp6r2kAqGnnH5VEZdck1FH2VR+hGKVUCfCK0PH
Ff6+XfaWPljDZnK2EmRfagKref2HzAbv1rNJOwheD5ux7uq/f3LS/nka4LvIwH1I7iGi58XT+trn
JitbbeDO28FZQdpHNsfLzH7mArrtd+Kbo4IWzfUP73u63XeN/aX1RFy5bXm7LYQ5I9aOOCyUJhx9
Lo8ZMPy9s1h80/df0wQMIYmLbthRvhmSeu7zdD5A93v1mxuol2KpSgKNBlHczFcO3eBIajD9Mkj1
U8mMrlF695JDgjyLSuqXayPXIbibnZQqL1aN861Uomj/JIQvUA0FmzIusXTUT0o1ymG9+jnmpjRk
+xWYDk1NWT7/i3JKw5ZNNDAw1aqUI5M6oYP4a7FKdKNBKQEaPMQdz7uLJ2hDxp6OwSC8NXRp3Ufh
ybl3Ad9vkesI0kVNUbTQFzAERHgu0ctf5RXt8gdK55wFF12a0IY8Wxg7iSZhAeEq+ag9RMp/FbjZ
kg0igPPlBn4aQZdwbjhyucD8d4OgemKuwdPWuFW8mb5uh2OTgyqNUXtS9htizI/IWP4d9nzy5T08
scmp+MN0hLlU3ccjAIli7FpyMnAfa7qG1zwvMnS1tNAzgqy4kfkIRYkLL5p1r/BwYP2kVi7v6StW
wfFECXsdyXdHuRyDl/oBkSBc9ehwubzIwjQIPe+2jpeuiHE9sXvZeGfB5yCdzUoz+ZJEy8pQMWSN
0QPWPDE7IP81vYxX/GbHpQMU0WXuhujj5H3taZ/5kBkMEfxekZ7ySmp1h6WYnk2jtqXkj/6ZBaUP
Etl2P/MNOuNNx0qlifPuzAbbjzU5TkE6hbRwbCwCcyx43kwKOrEZJCZll94ijXZe0q1IM+72qAZh
tJXJpj6LLkrcNn4Ly15JLt1g2NZEDPInYbF4MKElIsYQL5SPbbnJ0qQq9N/RBRx7Lq9zLbudQg/J
RHY0C2hBTomlE1+86RWtjffNujnNVsFCp/ALy0+V1ZyeBOKnM3zw7TaSEoviHZJp6NsYODyBilKp
gQzRvh7RElP+rnGIL2rj3aYkB82pMzC8Htv+g9bfjWiEB4/r0EU+oCRUSlFX18MILPCAH0QABNbE
VeuAnsIuu6PMcKQhDEiKQBNLJk4tKrDF/Fce2BqWWbIfeCIODvkYNXx/pAKdzxSEdifWcnOsToI0
TcdOr1stlSGk7sXOoOXYZa9y+GsDiEK8a/EGoCZaewzX6rLx1RCWlSOAZ3OnY3GJUpBBDG9hzUjk
/CpeWp2CXFpoew6eZlejc+g0YHJCW8AKIgB+K6exi8RetjptuLdcaWNPsyWMohWICu4mEJyNWnDb
PdBWgKT8pHEEamTlL4AzvhcER5vnnzZSp30JJzchEIHitGcSl9XI49fWXZ870C/Or7VB4I86asVZ
2dTS/tHLuBvglNXg/z/3Lv8jnHxyJQkAWIyt4oUW0CWb8jvkTzR59hwOienqTp4Izry5ssVVb7x7
BBhox1ZQYHxEZMux/Miwq7BG/ervZqOt60iF9EeFs+/Nr8JrxiVlfpeNPceSYRmTsBD0kta175y9
Nya97pzMa5+Sc3w3OoWhDPGSa9SusSAry1TrUPV3KFA6cx5io9ODr0Vt0UkcqBFmzhP7vBp12NQ+
QFGI6QFMyDvrNB5+Aj96TYDXyfE2hkBtn1JsjCsf3hKSqbAPYuQxF6LlXHwDSOLrZxkpIKvFApfz
eBA99TNeNDSCUpaQkYEyWkEiDMF48xfjKMj9rZFYOOf7qObOdqdJ0iE8x6nc9e4CelFA7AdHdsR3
iz8U/3MQN4VI9i7BzOfmLN4eHkD6vgDju+eOc3uSGM38QOcH93gvndkKqDD+uT4tMaWkPxoQccqp
W9NYIpzogLSGSkQZDrt4TXsoGt6DCsr+ldIZGLgi8tSk1V25PgOAe3mZAvO8C8wA7tSZ5LsdKQkc
Fi3J/Q2o8MtLsiCV/XpcxbpzasVdqinp0iQVqGwOO7GkBdEERVxdwEONCsKhuGAKpCF48TSMhKQ9
5DpLB+AysK2y+QYHcLK6wqO5JoFarkNBZsP8SktVTdoZKLGpiSJrn1QVGDdVsXEbHj5GTiBsQaLg
cgZ+tUE/ySS8zEWRRGPfiu4B5MlYAn1sb7IFehsAt9S9QkT0M03EtCKIqiVnsoOKGhbSNpclrZvT
2mmjs1acAc0qnKwTc8GhYOON2E0VxI5ZKhwajEb+gVN2Jy5J1nL5PwyEvFFC1zgECqnBVXvtDGIa
id8RTrZGhyqkOktc4BB/T8WU3zqMLuas6IMzPeyqAju2Tls7Tgr80jB4p5KsIPjbYmdpH45ZLw7c
nzBwIQQWHb4KWimt+CZ1dSbhUIVgUVYmC2nfiFYgJZEluqnbAHkxEtID//Mq3cEtCEXDyxsMiSDB
i5HdkHuP/rDzStJdF4YqjT0+JR7/iK6JnY6NqpxnnpKsxSI2HTCnoGFhZ1r7MvYiq2L7KEVnMZwK
6APNJ+T22MNAMpiI/FZTofZ+NEuAtRQqQeta/D18J3xpMEAIgYY8abJzi/nUvfXzLPD9pYl0Ao2H
fqnrhXR08tz6hAky2ZP+/zNzDjAicmVxfd/POduT/wb7dYX7mM6zv9kzR3WztnAvNam5j+LrBED8
AyHO9whLIqriuh0HCxNFImLL6tyY5bTFCPD7PfeMcIizGnS3yZqFE0E1QZiabBxducVzAEdlSPVG
v4x5bUJyUARAgAJWMHGIZAQXDrQCW3Z0WiShOfmabrMXgqK+78cULxRhNQuDx3BZqQR1kM3edJXd
7gVqGkhKmH+FUUKrO0jEx7mD8qtSk8Ra9Nhp//E47PaVLvUw3dTQmqXP/dHfU5LTcU9wlLWHfkMj
ki1EXMtOyOikpxzxANv+bb6wPBIlCjo7IN8fIa3ECA2q5OOcRWqGI0zceRHjw5kcHVhpH+s9KcZr
XteIoZcBQEcoXydMvsxw/Vcro6sN81XA1oetkkrD7WESlO+WH10dENDTOYIITmRwFZD4Zf3SuTjE
WDmU++DJI64WhWYp15ahODBgZYw4PXRkAV3h9hNOEC3bSNE+NnPaOvOG/YInm7+dSxNC/Yz6nb5Y
LOAbvSVjLZiid/PZNc8ycOXGbjiBUv+BE73rc1UUUn+HewnDxvF2rQlI/QuZxC3GllSC+GWTTtad
Fbb8/skBETZ/n4QaUe3XyDhVlBT8/zYp1teNFaHXKAjMuEbngIumoAyWlr+TMgNbUjqIJKoXUdGC
CgNwu76puFaUqC2GPvUtXbi8B1cIOHuvpW876rFOHWuFRg2zVrWN089alwhbO7/NagzTbqP5rJ4W
GZbEV+s5hOC6zROUg4eL+fd2lEeOHrb70Hvpm8vNB9eUoYnYLyAClZmhPa6CGMwMkPdkezDs5JQV
iVipLhcANoXWC6ILevep2kWZN4blJ9l9ALOMlowB1ykYqqUdrb0arTOcBAEs7y7YzRjFY1uwi2ID
el+jOtFsISEcyIjWUBsnKC4Gv2kiGuaOomLbU35qSM5mIHJMuIxHm9lzkOZiNV4Ds3/GLJlKmyVy
0+QOqgX0H7KJV9Vr/I44FFrci7JJykr24TYyiTallsdTi/UCjPW838Tj8zInG39kdxqk7fr39Pyy
bfuKbCJHrBiQZz+m8GYtNx975eV0OBGzlLLOhHdUfzGV7PyL+QKT66fk6OtzvnUYAnrns30Ytc1v
PNd/6Jasz7jAXzn4UE1jB4GY6EEtkd+HVOPurRtXsbrfP8nE7KARetcABMZsWo6BIHdOPYNuEQUc
bvztNQMdy/5NSoA0rL5TXzqHLtBbJ0eHjY+DlQ2A0AtL5vmJVaMxC0h+g6G916Mzmyvqar3wOS+d
gvHhGRAcqf/w87egKFCgPyhTGWuNzXAOV/GRAZxIx35LpsMOGDTTq2l1L71GYJVeGdmrhvMqO5ZN
6IY/C45ZIzDT6Q8ghzqZYdeRiOBnyN7j/rZr4ozx2uqfkjo+P9M7beq/qbTyCLXj5/bayvJPx9V/
xKTAAJKx3Y6AgK++SqeX88EWg+d6BtXr0A00sJKeYfJ0VutO6XK+moY4Ba30iZpQxc3pTQkLHSl5
ZNZREEJHy6/sO9ss5vPon65wA2pyLfGM7bK5DSujgyV+4E+dz/w49N4EQJQ2wd0TPzMD+J+Ofu6o
gZYPjjfOsCR5N20nWeK5ujPFGc0rZDgovrgJ8FhIP6z+EE+gdgiIAh8MiyYRl5sNLSJDUspKYHl6
v31pxhqqyG2dI8YA0vMlVH+wCsGNRMxfTJtcY457uaN7YRvocmgrDLihDE0hGLiHT9ybv7qAFcEt
KBYAY25kN0RFlRB5lVRMNR2apa6ChMYD1PKwCVWrb/U5OH9zlaTh0NdwV2Fn2wUgPmF99sm8s1cO
1H1dDAx9ADt38vKwehrcYAQEqh8XIgUbkyqHLfL+RUgp9WUCIhFtTcGKsbXcm3yWqdTOy89JHePo
ZZm8giMqY6GW043xR97btHK2d74tjtE14L6JAoHOgR3X0E2KtdwVz3h3YBygSNZ2XwRnhKKqoHHJ
tGb4rCthT8gVqi5+zTz2LrhK8C3KTkwtJdaoZT7pCCVUnza+bHjxaK+EgLwi6cntKNG1v1j6FtLc
5hmZzoH8X+uk2ouFwXi81dGZroHXWFH1IbWSkiBKSLUg+TAapjK4XJTcfYHFhZ2IvZLO1pNT0ciS
A2tls79d8uxIxm7JNShKONJdYQg34leAQ/60nXL+V8nuVa15qAj8j0eUjlufpRFbBTlOIeKrOWGw
Jm6VS1IxDkk0v/dGBNGziPAS2mqMBXXuVpar+74dnCpqxpyvl4cx9/hekj9gjS+h5wCWkc3FTn39
0QGkz9oCFq+AtNSEVpmgG/B+0eSOOVEcoCS1iegOif8fp0GGmKI68Wi+wTbrfagDMXdtCN7zsTOC
hcKTmPmKlgtTK+AVBdZs9gEE2QrKv6Cfr6LxT8v3a4xVfJn4Pwiw1g6u0PYMbAG9uF9UmHA2WAoG
7+eAtaBfn/aGoPJFh+LayhBbjVzKl3erQBQGzuGAjYAbubKHGrt+kE4qS+O7dyK/bK3nfiydAKKM
jk4XQcnic8U7I/9kJhn2mSyH6iQkWX0l8MvRU/uuP18o6VH4wU6nwFddPVj3jQ1t/ctyk3Ytozn2
E2DaaYI/Sx6v7HWW/OvoMWTim8bJ0CDmzbjOdo8cP35vdVdhuEoUeSPXHLmJgJmQEJuIBETDny0x
dQqFIZ2X7kO3rrKMv4EGYLOcsgEQBQp2oGxq3wnNSV9W/4MpCJ90KMwIKi9U/Z8DqMC0yfrDYngO
FtI2O0OLf3zig45q5KF3paJngA4HkkmFouJV+sK/MkAYCn6YubTm9t87WjVTvuoFfh6YgFMnqqSb
Gryh1YpE0JRUuawsfzhc8Qyeayx7xRasXgBZhp3XxPv0CqOOAFv76p/V2VjeF7J2iOXm9B+iPPMf
d8x3tB72nrdQNObLR6GhZldS2ja2vRJtvE+vI33bnT9vkbg5tWom5Y4F9htQRIcH89GMBDApcq5y
fGUUDXlGQbGO1NJBRv4IMZnoP3sabkPlV6pbXBBwOvtFLtx5HTOq3cFdkKsBLVS/RwQaHx+zqU2u
gTHULvGXYPyOKIYB8RDWV+P+Pdz2lmWqv7Ctt5xuxfIF+BlxJHHpl13pIOfKRqgLkA0IsBFCAaaO
snapRQn2bCNFwHgrzkE0YRlEt02uS9jSG/XHHDV1iWKJRizTTfzfi5OVJiUr48RBpniI++QkSCbO
E7koS+4xeyTbXez9syU/f1F3HlWw/pC/e6QHuCa7aCcdSOuOwkW+Y81C8bqU0fRRV+Q6kUmrvrSp
N20MQ3faAcsbJ7niZMGIkKrRFTDL2IJf7N2Nj4BObZg9yKMsqW16NPz3O6//XU7RSx0Qt3y7Gj8d
asgyp01aRo4z0w90Z6pHQFy632jWMYreJFYMxIZSNDEOzePR4SuVF8rZD2r3s9XPd0aGMVQCsbkr
RW5PHdUL1uXoSn0THG49I0b4vZERWdv/vPo//gEPCvzVcIpsMFcC1ZylmmDj4VXMpEua2EoQppel
3tqbwOJvHEZEl/WKUZdqEMaCcybzhqwWUC55x6XlzVN/EDgdKsI4q4jpJ8mZyO2dhZzyGG3b/6HN
Jfi9YOosBFJUM2emqzXn+RFVzbwxKSBEzdNHmNp8bqz4JsuWth4AOOXKOF/Wk2qhxUY4N8R8Zbyo
lKfE3vHCQoQ/HimrqHxxWHnrJQEm5ZAc/5waff8TjNjN9qO+JaLd+PLor9KlPCkxh7ut7I5s4XSh
A7691SX/AENsi4rg+4//GODIAx10CQZX946SQVRbWWSVhS1HAP05JowJSd9+KbdoIdGxWxDKjRC2
Oq28ddmko2hgefqBQv4qAsJ8cmsh3RfH+ni6Ki25GPc+mauuG2vUjlCjim5eue1EnF4cRiLdpPGQ
1hGNd/RWNz92wgqzDA3Vn20H3n1A5ByQMshDrCQ1DM46AAjhKGo04Gr7IwnmQBMGaUdX/GO7M+Yz
a/iXpu8CyJmut5xkYCTR1mVDCmRIeA+3IU0ElNNzAzZjOY/w6fh+7PqjIrFV4dae0nI2DR1/SdDo
7JGkdZ+aMXWA888oUmAKEfKKQx9DFizt3xfcQK+ITjfqYb34BagQydDTcOw2okL1Kyc2UKIn6soH
bA/z9T8SUbftwiRENNRM7vUbAIvlibVdb4JjMatlQb41isLDrJ9RWRPEIkC+V5RuTl6hqQ+2LFIG
xpYIJeeu04MDSmyBezxF45DeeCDL9epqFjMuEoRc37t9u8Yc9TXEKfKaR/gbmWM9w1GnqXOe2bH8
uWH0OUNfqBSBdah/Pgpzr4fD6bXXW2RghdmFpfp9VwH1PEEWeWYt+rVITW5QJ4jahN7zv6sSBcKu
5Tu6IoYQvY3/aBk9o+ArQhYj3jjRWI/HUiG3XxYT3ZGA1oeLp+JwUYBFXvZjGRWLs64qI2gPavYw
hferS+qPLd49Ec6a8sq3SfhjzUmxnuffIAFL+fYqjNNO5O5WEZGtC9vAp0L2irYpJf9DsUUTbVI7
5rUcLL8gPMrlNx+JxVepEsIIn10xsddwIcFzchxSjZa6+DiKpvC4lopKhxjZwTo/KKpPAgFV8VaP
O6mYqud6Wd+FBig4hCqydkUyJAm4DM7sLdHIYozVvPq5xf68pI6cRbc+Ee4KzgZG5+Ehd1ijQDKe
7pC38pgnks/uAjrJO7eJB33vZm72nCj06r6160kNDUJQLwWAEvulQjg5Ftv2DHLRKaQSdontEJNh
f5AvAW2O+yv8QwUTH0pAPuCvC360d4Cv2YF07P/b6B5XZ9aFRV1Dvv5OKA/QiJfJ9dgPnDOaCPN9
zqn4195nIYTP033ozOjHR1/MQY4gRisrTbuCuNwxMt1URPsTCxQw/DHKMerOvdgtCQeWXV46/p7h
TsB3l5ARKySrr2gdlSne6uc8xcSy78DTWMWN+EBiMwFYqCVXdH3doXV0y51ynG/g2XAFLFaflR7z
wyvHpIU7oH8J9KJdqVK/N5vPmJLc4NsmGZbDPboNexf2ZlACEuXvnSSjaKKmxaXkRGaAenz0K3pH
OT0bsyy7/OUs4PaDpeTDugn9mlOFjM7X0n3GUnjmuDJrb0F3N18Gd9sNgny7WXPX5Fr2CLv2n/0d
GoupIrvMY20T/a1QNL/IzwmSQQ4mCzjkehRYJQYLjcfBamXAn9HB0qoS+ZwDkCXjw4b6U5rh3/PD
tAvYZvgC8dlPYs+w+3F+GfBfb5X7hnuyHUy6/bZ4QzYJhFZGs+tWMTdiSxVig/wWKKfJzc9z8emt
J8UE9oPXGE3db6jon9yPZD5CWk1IzTW8n0xvZfXMunGIj086ctvYJL2spmxtgQH0qVxfj6F+/4OI
U6mfkKxbETq5IzoDxg7w8W9/ug0E0B2kls5jN7UvDhtK0HepEMsyAWfPdsS3J5VUByPwxdd56XD0
H4AN+mXAoTJEpsprPXcGtjmfCsTyTMpsYykErcSSJM9txmsqTa44ODMK+8X+/Bb6Hl57AmrHG6ig
VOXmGgErQPIu6P5/4VSczdnArJH8QznTvnyyhl9yBitkGNsII4pAD2fmQg3AJMNNcatAXJ0HhoSp
9vBjy11Bbvg89Qtt6fkeB8oEuGPPAIiRr6zH2vezUdESVuVctUnSygwqM+TWcbPt0KldaWTVm9rz
/sspqoHvYVopfviC/WSkmthyTC5JhJNf7JbQtZs66mDofzrEkCw+VWiAgzkfJFk1EcPhUb4KVK/D
RCyTqZGntNiHMPwe0vWamVNNs5G/mGQ3fuZxIZvkoLupVpO/KYs0KhUiDlGwLn2RiiLzE6L2KF2s
jnAk+JkAWNj//MR/y3EWux41yVnzcOR+YJwuWlX5bC02Yndd+qkFW5H6GZXnonf7lLRPp8hyNYih
UdgrRgcp9UTbQwKxBvfIFRko2D1p08Qontf+vA/mYqeGy3Zk2o8050c78v6OBwTYXL1/HTTKfF/h
r0ID04vpXkOuhf5vGqTLt/ZksXe2SX7CCD2oA4lNogxnh79aOCwtQA0/1U1LSHOY1tYmMxTSRD+j
ZbfBeIAb9B5NWsggACDny48+W2cPXWOOKIQHaS3uzp/zIE8vLgQI5Bkuw8EC4So2Yir7MaWL3f/C
nYsT7G06+1LKQR2xdsY5HHjDTj1tkpgJRzlQlLUw8UiHYPrRPepBt86UUxN3LieHTY2fhnphZ3A6
d1W1FEoX4NW85x8ZFbm2UUb+1YomOjOHbtohy9mBlU3Mhs+iuVDQlCpSJgjrCzl6eNobYb96aTPY
rRoYgF3jr0e7YG0xcdKuFhtuWMXpoWNPI/khOPRNYt3dQDBY0VeIZCZJc9MwnTSM0XggqHFD6T9J
dJ0QWT2BzMYSWb+1+twedrVG8mMT1poBtIQwlP9bEwIGq7ce1yzZRkyA8tLygyT2ff8MYghAnJWC
V2aQAWM5Mu2WSrj2IzVkvT1OI7RpXnJHLq46WSZLkHT7WCreme8QyT70hSnstVH5zITB6OYjp1On
d9M3rAHGQUJi0ArEn3j9bouEXWyYr9a3LA56c6yquYjlNMpo/YZ01sqY3u8B/46ShZyHMR6126lK
L3VAagVWaQ+9HSJpGkeKoKVIDWeBR2RuEpEeLBUD2+iqp75YdVDcqcwIwyLOwLhECxIAfZ9mehMe
GGZGkTtbz4g+vP/uAOolc7HpmSMyx9M5ayyGiS1r03qisCy2+xONbI3msdblvb8WrlJUKMG0XSsZ
qKzW769QtBBX40we0Gmg3nf4QjjmId7ILAtjbzVtBFyaCI1Xf3tvZDRhYbjBKZJI6CYxNhSo6f2X
mwt8/QD7Mj8YYSgUxi2Fo1jjzNHAsKaGjQEEsDBGxub6rm/NeX839TgRWBXZJ/ByvAn0V7vzniuW
JI3F2TqwWq0sJ1j9X2yfWEYvEJ+yEAcMA63hW+nZpeS/5uAOKyH7X6QWzeORkSc1SSvZyMZ8SSCt
n4lr74vDKKOwuqwCp9eT67lYD69V2+pcjA7WOam6pt3KPT3GphWC7IiHUp8LKko/RoNsro7Q5w6O
H03a7TZQyFqXaqEgfT3zuWFlUUK68+OZVo6h2UbABl9L368Jvkh8fPMBc2u6XzGhtnn4RdIUsyos
9109WW+ogspDVCyYNu2bKw4al8s8PSd9KrENZc30sylQ1HqEQ2OiuV6DpJie47R8k9vceOERa8+c
H8RJtHx4GzIwybCmrK19QYYFvW01QhRbGA1DuPJK9+amw72fbGdvh2NUiVmnKUjDLFHJK7SB+9ig
H16uaTOqDvfMqO2MSwJ4nv4yGZzsgwzQNWaiBZQA993hv8DAIo1Vilfn7C5I/L/+pGYFBScsS/Qc
q2dUwSPizjbX7A1dJJHf5d5b7cARGtip/pQ0R4y011uTj4G5zXTGDtCV+HN3/TVBX2DhYSAck6ab
MoLOvC5IQH7VjdpWIcKm3mD6wdbq/hUbhTobUUnGDXM89fE2PDmXilztmSocgk4CIF3s+EfVbHFF
ZlD8DqZltZNcihtD0i87pHVI479lDr+Pu2for/GerSqbf4wBVxNDERaeIw34Skk6tfwqT9nSFTFV
9jqhstOCmDAnBgw1ATe5cVmaDDe1bfjKD4fp0V8wsohgGKP4uW86fua7qwi4OKJanv8dMWSr0xMg
/9ZzGLLb454hS3SdTkdHdj0oAVRyOjJof0TwxRjMYJ1IDRkNjvj08V+u+u3IsJG0Q0BswtqauiXy
kYbY+XXpXye2mmCgQC3nDuO8QoWHwbiH1BQVOLcPYtw5AW33y5y15d8ZrY5VCEFMaVWxgtR+3J2Y
4D67YHg5IiAPop1lPQ5uyyOA/R2rWqFVlaxm6cNeOsQ92TQSc7MGh+MEOxFkQZRK0p+b3xXow3v/
2VAEVSy4RfEEDibwXv9jMDLIEIxa8XPlUaWUHfQoWnuUX5TW8938+QYXwSxS0gK3lKttzpYwIFEC
4Ae2cvCQ9DGWDiGfHE9Y7EBLMaOMD+LVN5LQeLITJjAAd/ReJHac5VnBWjqpuvpZ4B5v7KccjJAf
33ORDf7HrSXI0HMuUUMm6pqO8S7WNggiF+Jq3zOjxetUbLHF6WNgt9GPyFuAekpQMjYZLu1nu2A5
ugoK7pQhT3k3WTjGCVOK8dVJW7lUaK4KGhz0gYFN9ByxxTMBzKI4l9JInj8zWKvTuf6lYcCUnbJQ
N4enxaC4WZsRxqJmBm1onfXrj3qLIqIDgdK956osKxZ3pDP3qKLsF9vTXa56nARuid/vao909cSs
PuKX3Blv+nRGwA3zUqdo33WsT8MMaWR6FEzxtNvpn7h6NwzzV2bhapi6vUDlRuO8duYI8zlLHWfb
VJccyg4Ed5J56MI2RoW5vfhtAq05Ro9IIs30roUx3OwvA/CKZFaPEZ5NtLCBMyJhN/LsLitWyS/H
F3lB8LSwqAO1qKCWgOSS7vRjaaxKh63AgTnfWI2C7YiiLzevN8Y0gJdPtcJCUCfW6Qbq1LWdAnPX
2tJi4VW/+WvnPXUaswPCN9jQaH2QfeeMSEmK1fPBoo50QNuxk+vX397LPcGY7VGymY3bzozrvwNt
LHADavVmO2++8bTtgNZVJYCmPjJYxOxwczWUa2JlySHV5qid0Bgl69N0H1c5xAJjdKto3fgR3OKZ
6tTKcpj+YTp/NbE27tPLFvuhi7SbGtRYeZiM5tntfyyIV75v8e+62uh110cb4YLbSmepDtTrfl01
YMvBW/9yk2M+FNSFX51yWginJ3TOJoQmPCNAwxKh2RQ6fGiHEV/BCeCVLdJEa/qvenxW0sOzxuqM
86UQcd7BL2JvgYDLs2EnOmTZr2Wq1SngJhgbYrOoadAFs0e3FLvvDVwSQZ4oX/qbA+dTZC5sQuhL
n1YpJP0mYH0ap3mN+iM9YLUF2tbRtqV4slhYO5KoskgwQ29rSS7az29P5pLUTrjAG+D2N5xoiwPC
95PeUkl8N8Iflek51jt3swYQ9AHcJ3tzbBQd6r0Nfy31tk5Kz5cVKpRj503VWv5vMQXaRrkuUvzE
qRXHulJny7mr836pIitxyAbz0GGV7t9SC5NHbh1KedHU6gUbJWNB6mtql2ThGmT3WJjJFyx2kso0
/FRe5OOhGDuTFOuR1yhBAoGsSo4oGAD4skzZzZYEetq7UaVXYUNlcdy4UDzfn49TiM38X0pXSAnD
sjCo58tFjKSxAFr/q3AbRgekmx3ztEeGIWnRgYiqQ5fE5ok4JyVsIusFphH2KbQT0RAQ+IDa8NQh
AX0sHsubOd6pPOw0QNF1AtcfCbO5C6Q3/0+Ua8S4uWg1rypiB+XKEAbO4XDSdjMqYb8qTBFSoY9v
iIgHALkKh9xLOUf1gC3B7p8nslUeJyDVqGNdbUi0hOKVic5tQuu+FmhEP2dw9E8VKOuM0d+dSli/
IpQynVAX6jYJd54HECRNmpajrV5BuTivuOnJT8VFlqVJ+g8JSiyX9BbkVcEfqU6wGhHKA2DquKgx
4hbcm7ko3CMqB6GwH2OKggpEb6c1yYhtb1SuO4RQrefVpYwfRR+WWd28TRChdjolnw+Hnhy6kiCr
pMnpGA9tScc9mGBIViudC0BqRQmw+4Eh6LhktyurSFlnLASCVYOVfX+GdrTLcOHkpE8qPBpRibbo
Xz1Nbn0Mu5/NNeX5oAHUJGnGIfz9zU3GPSO/JWHLh+UlKIO0RLGVwCoxTua3XA4QHEQ0XDlVrHoU
lYbOSQpFSu88eAkhqnypLzF+w4ASY+M4ic+ffFPyVmvSs3+0bmOs780gt+Lyy/hqBByjWZqLIKRQ
oJUDbFzNpduXSGs+zqYo/F652w4NlegcXs0aewkiRV7KOlfAXmbAVPTP3E4mS7F4OtYXndf1rrvz
7B0SZQxrTunPE0naOt/2DtYFS7rK4rN9dyyfyEungMiVuV6rGwpf2dP1dO6Epk2+pmwORhvawBl6
kqHdu4pYxW+Tqg3qd9cQS9t5/Nb5naegUzKhipp5/Pgu0QAyhsIRuVePW7tpnt9NTIIMbrbGNmkX
2AuqfrvE30DyRYNvhWynOD/JHyhNCMuX5K7xQo04m9hZquYtG1vGrnE2GjSO7obdi9MdYC69w9wX
/HOVsClKr9UBmsy2ZbdzjwFO2wmpdThUeqnkuM1AcTZJ/YYI1GGQvcUkcYOHjNiiVAq3modwMDAF
Y53qYvZaswS4Kirh8zeygHuo6dHhucdbbTVqT/UDmroRER/Bnwik1bL0YTz9MlTcmRriCWUNpz1S
UKPeHd1LHFin3c0EljG+tHtacNMfustCQbtM5DdeGqBHlQlVeJbh1Pc/y4w7frm2X4I5X5OOT9vz
bACxk5KfmNPEYL/niCf8/ZCJEDM3GhBDh8/9MBvmsOzJmkBshVcq1q2OvJJAprtnrztZwvS4d7l3
WUlQfMgaK187hkmsQPezqj5oFJY7KXW4qAIfjHhzYhKvlg/zP0PxkscXbfz3P6ReflQfaRW950fv
bN6arHTq05K5Z6/6H1UCu7i3IWwulmfP2z38vxRLW8MaabnNbX4tIAqMDKYfD8IBdvxxbwofJShg
zzmXmy3k6bUiYYVBOOZbokUs2wrjH2195ZgMNVcgNUkwMSWDfHYdx8QaYTRboDq0ZnEMnzWWQ39p
76pdMLNdfPfN8L0yL9M7DO8p9Ez6up8P2Id0YPGeJTgkd+1EB/SzOQP9wuciNLxYrlNAxG78O87h
pISM2+yPG4OaURsZ3PwGJOX3D3N77u/d59PUxLlM94gYNJmbkFYnvvaOKk59O+CYtgZKm2J4rDNx
xp7VwaS5rZHjjCS5PtASj9huu1nku0MzqViEpoF9az2rwQkTKPG2ZcEMq71t5kSQnlPCshkkwERk
2TLp83nbqStbwb9flLVJ1uX3vKCA4oduvp4KK6jVejP850qeGaatW6VP/gF0VLOd4UoCgToO6+kO
kPSjk7MWS5mmK/U+6Bqitfv+Rot0cnX0dcVIXEEdsMEY403dh19brUv8a9WT9kjp7fBdMGLzkeVP
s9Eb87QYqoiGQFnkSUQk+hXPMcyohmhSVd9udy9Me6ctNpxp3Q6Bsm23tQBlWwKx40cmGWK6aSuC
XUNtboRdHRjuUaS6wqyFgleBSYEIKGBbyTg51pZpYSiYvEN1uap/WZezlFizibAGTdzeoQecRR+6
8mnWpMHAeUl1qHmXW3USEPTX8cmK568EZi0vtjILhKkPItU0DlXykjhDzHX2nrJ0d1kiCYvv2EsE
ofnfmEgUJ1mTNkYbn6+QvnrByvtKOL/NJzmwAWFBLWU1+QLOX3zzebtLCFndL761j/1SfVfKMnE0
TC9COxIL/rTiRwxxykiY+vYNn+RN2mD6ngeFk3nWxuep7yAIQZleN74r74esIowjmYlOaQbqkX/2
AVS6I/Yb/jQUifPIMGdCuTRe+TnTd4NiLJBkS1dFgXJFzlNPsZHTUWiFdKPKCf1fMEWYEhy2dckx
YJjC+p6InhbdYvC3CYb+HD8hV2aXMNR2nltzEqmq+LyJA38mhLSNsFhi+FmpXMuFZ1YACpJ4fJQd
/OnEEJIcTvKbTly8+yG2/Ho5u+1CSk6KTl0tpRasPOOkcMBcOg/buY18jt+sD6rHfHQ2+GMT0oSU
k6sX1vy6wesq9A8vZYtiCeN42oYoOWghi7z9yGr3mtEBtI8DW48JfTX4os53bzz/lrW8MUzYlUrO
Ej5MCej2sMHew5Szb9dwQhkCaPij8piZwrNBmEz2t5QJSuRG8/594MBqtnziQTprou5AH/wtjb6x
ilH42/ZHMjASOlRj63L7DATelDRId2tFTsQn3rl5sw3XMClAaD+46JGjf1g50dS/ONkaYAUsVeG1
A+uAC6C6qyCReghyrAv8j4q3V25TY5xnlytk1kQWrsmn3w/O5o9UTzH16Rj+NJfwNAvVd+dAuQmC
AlVyh+D6uGu+qps36WgrQXGRQeIm2U0fnSq5dk95a6sXozX8U2NBVH+WvhvHl4eJq5ASXsiJCx01
c2TEl5ODaOJvKbJlmGRcvcMQsRTT+iPcC7mVehWr4LLBaCPWDFJ+05GOXy4eik2DZPZsdOkRwo7r
m//dClkbFZZL6VhX8t5fni0mqjX0WGnfkJ7Xg5XkFU1WIdplt2sCBAoVgjKeLWXxjVNUwNnk3o3W
XO9orqQ+RAx3FYo7QvLzVvZbb1owKjQaEOLlpVfpD3UXnGpJ/RN+TQJJUebL15Yjcvka5Lr1GrQE
WSHB7UBkSpd3HF35+sN5x6nSuk+832yfIL3zEwpg/QCo53ASFpxBTwZ9C7W5auOvjY5pwyU++iXb
ok4JlW+pUK+BCEJlx9A3KBkHFn7aLXFu3uF2QRPXptbeaWYhQAM7xKg/BvVv589eCVc1MFjHxgTR
yPlsttR5w00WLDQagKBNQoj7zO7GmRZS1gnBupp93mIuY/4EMm6b1bPJgAPOJl7MLpD6s0pjgqVK
jSHYAw2s+sqgIBO6qUB38XU25s4FmrgUBCU1rC5n1+LYCmYOearPyheWVd/JF0yl32PkMez04r94
UH0DyR8Hpi0vYT9vd/zNzQWm5INVkaDiieLMLxpwZBxK2tTzqV3O6plrldMhLzgHwO1pb/3HqU7A
Y7ZgQMnD4vBg8qe9R4Cnk5/DXGONH+lOVT5Q4Lp95x1CHWP3YrPVLmzVd+VjuX1E+kKCqOy9j71c
d0YZNWpDQtfk21cLBQh1+H+ZDcHQBDI2FUQ0s1c6C62GFixzn9qwmtD5nIT5Wv5QH4ZZnliMq/6z
Wdg8kTjd18qRjNs4yxSHhoPs2F0gZ4LxAlIjBHTI7VR6ktB0fCdWEikwpn0fBEstFOKAcAo2KDa7
hjQjhy2Qaju1aZqkBfrONF+J8g0IOQ/LdH6OfH3rFKr61kRajFulBH31Q47IE5rREcCEX1AbJ31s
Eezf7T+8r4+02pbJg6NDPHAbI2+UiHQFHkFYK6/UC0f3J/JvvT1xPNObAUDj6/RFyA5Bd/DTT92m
5F+AdnM+qSAHmUpOGkvUeE7lwlsx3L6QuKOHyhCC+CDFxh3cTEspE8n+I791afmQJ84bA7Y4DPPD
B5SoVnIHEUn638VmmtGE2bibDEzp0wnCAauIdIoQfseaPDpuvPaf1KbCFKLc1aRsbYlEdkgpPH1M
IKtEdI+VmpKbWy9r7b7Eax1Gsl3kIBmj5iOLmTP8mQ9zG6FkO3AN/V9w2KnJvMi4aBbrCXvMxtAk
KeaMBrbxrH/O23fslV92tg9pEOECIgVKH13e6fMK9cbiQwlXYFt68C9zS/DAqHkLhh0MB4I31QHm
Ac2pdCS0FS0ewVI+yxvDF0Hs1r2mGaA5iJXvEds72nwdHEBkvrhXz4CajWpqfEQ3LYHpV4dyAXYJ
oDyr7L6ERpgyLk1BjYQ/+59cKobTCAneVPb0277s0kUeU0V1GPABkkMVCWpJ2abhhebX4F/mlCJV
WqTTI4Xxk2BrSfrNyl9aYxWvpTFEvAb/DnuIr0eleAT3EJBK2gleYPfa1otkivu2NiNMUCDq/AJE
/r4XVvUAY+Yi64e3MrWXbiXRWvZznVCjuXCQInLrr/81GDQ8jo2beUV+eyMAu6VqZJR4qt3ICyHE
OdZr159j4mfb2NTT26mru90MyyTpwdT707HK+OBGSzU6zuHiQDwoCd643EW6EkndJ86zvS2iJ8IU
bFwI2/GefnO9hI+ZBQR1GK6QORw6OLK5eDsVtHNTN1HuerWo9extfVmaLNc6Bg5vihGBWAvALRVK
77HwpKTvA8A8IzR6R8wFlF5iLV+s+i0uFjTZg1Jo7FnzptMU5VmvwpnycS3wZIM9FQi1SBLocnvH
1GqMDRRZGIkqtPwld16kWtSmgdKQuqGDL31jTJV4zYVmmEV3KS01upmkc0Ms/zw8fjq7RxH3W98t
Tf4R2cFJLsfiWgfECwvwVSpoErvY+kIkA/Zolgt7mWK7tbgR1y2BsHAMIhbJfwE04tIFBfTTyGZq
9FTJ1ZIrlhnHOI7Z6numQwPo23QNdm5DE6GNoDeL/SoUP7RxTL3T+fQ3ZeNzLrX8weZEqG04q2zL
w/mskSjGYzFcJXKF2tI/yGnzNLbkUTleilP7M2zjcNuDwOeD57xOh5HwS89HoZ2IpkueMtoy41Er
1VEOF0/MjPgzoe8YOxXDgKGjpn7InyWGFQMPMm+n34b3gso/S/eHMZn5OwylEaAvaV/9sZbqr6nj
uK7Lw9+u+RjgyBR1GuvUW2tfA08tMcqFZCx4ShZf5ZduzhEjQgCh+xZxEAcw05TICL87A7my0v1s
1A4g0LcAhKDVQY8Gd/dyadDhVRQ2Qb2n6Ll+CDlYea/YE4mPYz7MvUEaBUgea8uSu5kqt1B56DMA
Xc79v9ZIQPJwv9tRbSOg7B9ToTy2yW5Jh11NOlwqXK6OsNzs7AKbGg82brqVoJgM1TQexgpebEp7
Ij08qw5NTj1evIZy61mWU6dzIxgSExP2NE9OILzgXWJUm8QsOZ6dZ2ZBk8U5CtcpNYbDbEZthoEL
Nz4ORSuqF/R9FUGs38+LV82YZ27ZTj8QyTZttcDKDcxj5sz9JMpqBzyx7W7fDomIIDwVTBN+ThiU
mE9cYh2as2WS7aH0WQdimXAFq+PZzT44PK6fHNj2QiXKOWxmCylIUBthvbBOJff8PyzQ7eBY2UjG
NuUH6e7qBst0tX8ktbZaWae72+EtgwYe19TPPiQmmKIdefrWTp1+maNTaC3YqD93BSOZLz5vogpV
IuRy/ILx2CKQYev/r/VuT27S11WMhXEVgt2SXyjbIl38fpeselX3ZvvLlf2BKMyLQTvqjwxZeGDs
LFAqG1edNQnECa51W3oDf+18dekXZlPt1qYi0LRa2279MMlR1/uIzyEzHiTgwIXVEKLf8F55hKX6
aIocxpWgyfVePtsz99noyLWICqWFm5Ui9NzLOsWGhSsfTklWctZB6qQYv23I88sM+yoRhzuMcMJr
Oy1ELsbV6Pg51vp1g9Pyzlt1bMAh8XZWTTzLmMhYpATKQRBGIS/lCjkkH9H9FVKCri0DKT63XxCH
6YeMSzVC4XpsCl+agMfm2ng/wuD6ugyuwT2gZM6hBEK6iPbphvfS5F5LzyVc74zpSEjgiFdGX/Cw
5EQ4B//exWlIj23sLPCofFfz3ksgoS7q4Op/K/fF1ySDY6m/n+SYfqBvQtOrSIxwnDOOmE6VnIiJ
rMWKnsDVgSa3ty9XHkF8gxjrobKLSR6/6xXho4+m1o31YE/bklFYxHSb284DgsRihA1+IgUsWxh1
kJ9PKKbv1RTbHj8AdtJ0Wrl529uyAI81oKrIfuwg8Ytp205qPfMmZOb2QDDN1yGoVJLqnhgttBo1
M8o76M8Jjr419Xs2+Aah+Ub3gNQ6bOga2PhjSeL+5rPzzTUws+zpXcsHQugm0qh+9B5GSZYK7jyu
SsKksECQhxZYY+la+Zpr0w+Jy0EkxT0DqyQjXof2y+f4MfTwGzOfGAemncnsbgHu3WY36wEhqvqo
DjLgaQDVkmxbRpU//GlfIUaAJNsQYw6tXIQw1KepmmBE0dOMAXgUbd6ZWHTdOYxo5yqBdRc2mSVF
XVVI96c/RvSyy5NtrrARjYxAJ26Ld/Ay/j/9L65zukHX4D4YQl8S8oWhh+xYwdJdPMh1toN1e9Mi
tQNHVDeBWmseIZAThl1DriDktv3aKwrUS1y3IIwMIbUHRTns2J505DeZsNuIlfVyIWAipXKe+36Y
C4GiEtrKrgNqYJiaR8ggMkhrAQ3K6t35gHkhs4SZK57kwu3hQbavMCXMraVpGdEhSFJOBO/moCfp
wt0Q6WaM8du0aWAfbpCDAMKBQd5l1wrWP3peoCUJRn/Zn0LuMZL5wmQ0ZAVnuo44FG1VpjS3S4Lc
C3HYOJn8jYrLTKK7B9YcYnOCz5ipgZE0k+GHsLKvZXEU2DoKk1zWPUh4M9YMD9bX/HBh2MtgqCCd
ObecAHkh4vDnZbgSzeqgFz2hb4RBmX6NO7M0UKjLSI/uODKCL38toAu5uk3X6pfTDHbSiUQQjkmU
4Fgh25sJtK+ggW1jDgP3KeUlrHM8h75awF/p9oLsR0KOwf1EbjInDyLOOxKAksq5qy5+7GjgMJhr
WJ5tOlRCoEKRpWO586S7RraACCTh5WYzd2Ij6QerDSJciWWbhmEXOQ7plyZ4VealyEWboJUju2ix
eidj7Ru/NhsfQLsd3qx6Dw7A96zdPqd0aL9DF6g/mDB8PHtWdok4LmLttEXeOkn/g2EpiH4QNMXO
8s3XrD1H7QXSv1OpgTVqjk3DXg4DFYkbPs5zFKBspIy3eQJXJ5EWOgWk4TjAbW7C8bmSQkVLjE1H
vETVv2Wgw7nMZfQysJh7UwGU7Dv1TokR4rkSzmVWSwNSBvNmR9aZeFcdRycUzAFB5DWRUAHvs0Ok
PbwFuzOJq8LQTYFzL2PADpjOtabCShl/sMvGJxE8jVGvM0WZC2rzkfGT0PWGN8ASj7yQ8Ipi7fvL
avi1InhlxkkEVgjjpSbTlOEbMQ4JHZ1veCxU5XFiy+SDs4bZxehY5zuGZPaTHyKIkLhuBqwA0hTg
ZBCBA0JpsjK27Qu2/KZHstAbBDmShkG1kdolXNOrjiAiEbge2xkLT9sGC0RCJtws7GKUU8e+ddzv
XRVkI5gkSKoTJjJ4ETRqVdRsmt02HTM6MJvSbyO+YoTcwQQ8N2BENRsUhc2MjrmCOBS6WWJuDW5p
w5BYJG3Kjsf5p0TI/SNArJBleTQsd7rov1hM0LBW8dxLGg6jVf2a/AB6ldejat0Ky/fCGk/3kcVJ
Shyg9texpEjy6a/yLUn1JbSVysXTSCo+IwNscIjYnPPdeWGuuh8sjVO8kvo4JKP0cewUed1bUcSz
iL6yfcHUtx3V1ICrS7Abkm83s6UL29dF4wFvgteRaT6k3It9pmHKbwODDnAlq21WUW5LXsu53ez9
7Nf1YcHdF4zIgelO36Vd0g4l9nU2IhB/vBYNy6Tr32SDV00J2gIGpibb6isIvGopLCsFBfigU9Nz
q9xAIFisleKI3t8TAOnB9ti6APTZuJFTjNgqtMVg17htP5KktaShOmKzmkDbr4MdWL5QHtSJhSdQ
qs/U1sHs65dKCiCnKUbR7d/JX1qberEGs13oczaHzYi1qmJdIEHQZdTsRmpMCoZQ7qQHi+YbgYB6
QINqU/UVYtzl4ZYBezJs71kIZB+8d1/HEGVpCBnhPAp9eHBt4Q2xIAuS/Ni+dluIBI0cSbHyxWBQ
9UeqRfvsJaVPirrCnu++8d3eDo59Cn8v1WtbGC303c9uQF9Pj9q4EVy+SIUK8wp2ioJIA7Qe/nUz
4C6mL/G5+lpRwfUySOlXIuuvz1i+nnbck1z3lwCKr/7P1+moHWMMOicJ/+vkGenC58i4m3xNdmRa
zwEwsxlWYMCE4f7VF+gvp8FIBQqKTw3syb/taq+rqzvXkShMliK2LiVaZF75CMSXCcoPxVV/FCk3
3w3ff+w+HS4q2LyS+XxhKpxjVARGZG8uQwAzANVEPv7cvsyhsopkMCyuFZgPPyinxK4lcjkDHQDQ
A/8o19Mq4Fbfy0l5iTDksgIEL7QGmjcfX7MfFPII/efT/R4u1/2z+SQbRSvn+RyStaNTnR0f1J8G
7Ts46lg+xbj4NfeVLd0ezSIB2Zd1hNgG4mZyAqTY1hNnwdtAH0VG6FeTLModhETXXdV0a4Rvei/J
q7yomKRXPJb0UiQRXiehyHVKuSVzRe4+IMUgrIUTrxUJFBlo/YQx95IXAY8L5eo3Wy+fhtNnymxK
ob4++uFydSsabgAXXYq2XIb1jP1YUzneVQWFTu/l5Ea83ckLUz+AcDHyjqOqFYryunyIF6o3aJfi
X9sh2XMJAGpK+rrtpWFrrGfD8QKlsaNhUFuhVnPo6DFav1cINdsozLAZq5bAXRfO/I72OnvV8If2
SerKXOkrRsCEHzaYOeUwIJ5J6Djuyn/FaOZzsFOKXMo9LjIT6WphHUKdNT6CziANHf/c43BNRVtj
02BrgpMVhHoRKKFN00Xn+JIGlkwUtUETHaHd2RsXL/3SJzfOIUwRGXsj0OIzHsFrdmfobJdgS4rz
1cny/EIZuMKS+q0a6EhACqz1ceFTqONLIFEbd7638WfFqyOmJzml+4XdFp19cvkn0JvvvltcOCwi
cnyOGJicy/FwEPJfuT1SmXiMyDTdVDQzDf4ss8EWFL+TpCu5FUMc1dRWKkt8mTbnwpToAnsgcBKA
ihsYjUL5pJW4KFOeY+7xDFVzPAHfs3YHTchmhSQ4ZZwBY6eGNt/rUyRJj54zKPIYD4iowFpOnDvv
AfRsZnlxl95JahQ57kbXgw1ltDFOeDdeJfOciocmmCZ2mRB7uZnyRTfh6eTgjHvveSBemhx4453T
bYd0ngJb+qbb8KHkvKRrMsmKLPaVDJ2cy1DBp50SlPB147jbaoFypKqpdPzU1UzSAcS/eA3FGMuj
DP4bypiB9SaFkwunmkgk6t4wrqUt2XF3r+pjWWeLWjWHljaU5AMuRefb18qWcPikwhSevsdaCBrX
foEnr8Jc6rKEuFAEOlv5WMRaK2QlErWbuDKt2tcaa8zarBqB4gxmRayLldABxaNHmbSQqOrVf0hA
wbTlIXWG/NruA3JvkcHB/6Pi4dSGyL5s5mJ/ntYSLidF5fz+CSHnxTT1YIp50iJYaI4H86zMCbnd
jNToiJznhVcsT3CQ8uR+J94b1P0TZVprzn/za1vLGiQcYD9YfzzhJoY9xUTHjqFTxWBFUNRtOg31
RxA7Qr9iwjllABk5PNzVcKRyfAEzGPOynnerkm2pZCCir+eeal9Os9X4KDG1x2GjURofU0wSucXZ
6abWrnOc6ZsOexcKYx0bOlOQgfcxX5VnEYcVrllUIdqQ8VBS8yPOI00b/kCk2+ZzozSaTe8wiae7
NovRpRk+qpZz/kJJYAuPIqnb8nPs2wpWdodN/rU7VbjzYRWlaVq/u15GF2dMDDgnxrl3vjqLHYEX
1GVR0pkVtRaqhkAHXC2UnsGy03q4frvkFOAtI/nzfGa7S+Whmdqfpmp+Q2bb40xI87KALSIoVK+w
fsqj7You+ZTQHbVmyjcvlpUq8sPex/EQHUwF7MQFuRffKphUmrpYtKEafG1/cB/qgHPi6Hnsr1NO
W5BzjK3i0f8gXPlmaWzdCo17XIbyanQgN4YSbfcelUwlVebx0CbcRAJsfloB5A8hLvM0WO8U4gdb
hxqS7+eFWdq1dWfJs/rWd4fe2lm/LAkhg0SSmCvvwz3jwh7AEdoJCrGHn49LnP+VvvxeulwFyuy6
WQcxOwYvhZKrEiOuqlqIcGE+3X7W4ZU0OXjVOphaIO0Pu32DN47IUycAynfu9pTFLHcFDLOcy7hV
g6UCwSggvkBGc8T/2WgD7DOSxwR8/pFx6+7gHMiRCApPDC8s6hMtAZZHXmEmvOI3IEGk4bSKfIu0
HxH76hNsw2U7jwAy3kG+7ui+6aWDq3G9FNSv2+5qouMFED9EMdsalCJPrtS0rz1geRAx3fJtUrj0
q9ERpinrvQ0fYlocmqwUJPGECYy4Wumd1zrrwxXEHueXuBGeDpVHYXnzG/hgF6HOmo7aPB/wnv/1
5cthODd7qCEC+BwERjZucEa+siWsKvMRxWrBkm27/URXEevmaVUl/HsrgXCWIaQlrxOP3c7GCvAA
DkOtAYrk1uHySskeUCwemp7cKz41l2avR+slSpGG+H5NpQUEes1oPxFxYjWlhNfwLAwxPWLak/Bo
u+2qDVF5SFMBThu+meErPBYzn+KTdxUUZQkBaP0Y46hIjLmTJXTbHJmyAGzU0lgre/uQV9CKkkLT
iqL2JZLhwfWqW0LKsBbX7sbVVqyTvz9i8KygaYErmO4f7gqob1P70y0je/P8F0I705puZE51Jd5j
H9HzglxGB6oWsIG9wkX+Mx2z4h7YrA7moFYXAy8/Q4faw59qhAGOqSe1WdL57xzDnjd5lMh4YPbi
JiowyQnndpFCG4UNLAvwBQJ4sXFLZFUCZrPXvRh93t6GjA6hvfeodSV7zGKzpr69qqHpyP/nA2u0
FJZs1APpaNC0o6lG6fwKHptCmRMY394iAliyx75rebfAj4nDrQdUnU6TCLvcPIhJAmfayV+pqG20
ke4q71YzYUeBFAB7vFU1IbpnwlpVjbWgc9qfogFVwtPf4LDeV7IJVTcEtA8GGxFtWV7r98lM6Sl3
a3ufMFrjGbyTie2g2DXxrLETeC82Z/EwI9Zfpwi4bd91dUuJ4tNL1ZLgbN9Z9bARjodlGB3iRFyW
ipGG4V9k9UUIpqKNSCTa7GPbwe2NKaeItxn9FJgWwTEkFRu4xX/0w+lp0THvhSvsFlEQmorW8pPQ
gBZW7/DrE/gBzQOH1d5hJE0JZBdMubAtj0crI6gwBfGFUECAvkMWb97v4uavfkf09mjCqCC8jJzP
FDX5h5UfgW0deNmjB7g03Z1/EYzCC6gFk4isaPTbCfYtbNilBsNbA67yb/hIKT0L8YoYEcsCfwJL
f9ptBtyGTue1kAdEkOLerbjQ8xAXSVMjKHgiN7/mHBt1Vid9E3f6/8gYUQWFqHkoBKhiJk1ZdyII
tkEEnC6oN8uVn3ZLBsfn0VuXBHift3vGKw273O5R56X7mXrSJznrTpyzHBtaf68kXdnIz17oNQTp
hKEvQ+4b9ln/1XtzCcH0RWcYyIMHrZ/hHfeSU0059l930fx9c2e7awQiaruxCfH8MWpf3SFm0tUY
xyXpXodRVrWY9DATY2uYYg6oaoTBCJlFjvqZRXWcVVse+0lzHtJ0TA5eOqf6hxS933wLawel2wPa
r+/HMoTXR9ryKn6ZZ1GiDD/3xAHHYBkhTYUm4xlkp3DqOQYWU0wxvLxqVl1Ta9HB6xAxOwW/wqoP
mckfbveKB35uv3Q439A2LHmHvsZ6MBtwRTv1NmqYf0aH6M0b3pDiBkbzkdN8TpWscGwdoEcAyrS3
561a5fcJcqugA5rikcwzZy4fAAnuL8xtXGTGBt7GR0sOpqlb4hXNhPk+tyyZrkXWCYV91/RLb52n
1+SlKXiNS7aWhKyTznswX29BZLVTAsRBhX2IJVdP+Uo9JOJ4NxV+Qq70AVVXnStkE9Mb1Ey+5ALD
JGmmto1W0L3j8vT9DgrzyKW0NreEELGMZuwyzcUKiV37DBkgINTYP11pcMdSn0BxkB7IEKfBLyOd
xrNmHEolIeHt/euYOf/MXSgNeT26Yw+hWSxEq+fyi31brOzNy+vUstJ1cud41YdvFAsK7Y642DI4
HYZgHn5r9zBWz9keYrJ7+Z8tYNf/MKt3uPFuySS5tlukVCjKq5G9zRryDlTd+Afa0tMfx+2tr5+H
HimVzXXptjvPnRuimsd3OYD1aWeEoEdL6HgatxcjiExQ0UxPKkjM9TVe1i009KfjTfUI/WPhIJd1
2F1r+L7N3Tn/PjzbUUg1BDRDJmWuhOGaZsV0V9+mAc9KRiGfzp+uW8/FI0MI1BrUzEzgpdm15j64
EFJU2RYl12eYxAClmFxpKV5s2CCIc5muK6sIo3opYKOHDuvuIxDYxVfaGIvv9VwedOut1cIN3SQb
DMKUZckhvMF3RvifQzzznEBRZwd3eJbJNHDieRTT+4JoP1X8xL9vXLeG8zXejZJfwTLsKjbHe4lt
BveHi7xmOBxXfxxknHOPC+1zmQt59nIkyhWkZ+HvwzKkMG7vOL/pVng3/xyh6tFw4FE1QIi0OtkX
8ZHJHcFRRmR4mpeCJJvwmhOawt8LCKS4ODNlk69FRw7iL+0+zZQmaKVQgyeJ5LVnPucwEMjxrkuw
LpuVWkzhCZGlnLG5+YWXXduBvht3W4dwo19/tuL4z2R3ahGjowtgOBTi0cNSOjgsR8pX/9taGIEF
0gRYMq/wc+0jbOWrdq191mx28eNtOTc/SDztpKOoymsoLAsItrVnJkTQT70keQLNZzovn8HuiRW0
qxSMsaL7Lhi/jU8vol2iV+qGyfW7LgWcWXNYWduiA0NBj9In/Obgy038WXykJp4Gh06G9fjbH0Pu
KMRyuDnzTpiqnwa5I1/A+wc68JT0EWDL6NeUeAInR1SRcyCPMfQy0TxMtg3VFo2Vo6ADoDGJ5VwK
ZHUK6qqo+1GjKw6laENRaAqr2bOTa3dS6pb/POxvpv2R3MyyA6/zV4YsDzhNx3h8IQvEyLFaDkkG
mK1joI+EJDlvJoPXxaIWdGOvcYvkEC0dgQl1oyk7DO36mfC62uVJERXAX4AB8dPJQpa09CAEccWG
2Y/Auvgr5Ura6a3PmO7GEnrk1cokgxnOJXOtxcgU7LPl3TxXXfWO7t1JZ+sAOsyeHfpjsivuWGH9
KexujCQQAdeunQhMojzKlTtyg0cq21iOlW1DbbbOiU+dXjLaL7TZAWhPyCKgNEgpY5FS6xtpBNP3
FfaKr47f0O+gD2/h4Wc8OB2Hnm292pcAxlXm/rYbNG/TdMI2Z9z7h5bNG5CiVHlcxGHGfBthSiUh
d5UepQ+fMEAGfxw7Tl0U8UV4wYZNZqVsk9nobCtv/m5OF0Ck+Ri45SoK2NlxIxQEsArBdO4jPmn0
VOpU/aXcYXWt3qO0k4CRjBU/URYrAUVi3EMra4ecBNCoSrZ9y2T3CyFtnK74apSYEAwUBg6120ir
/eov6d4B8HWPL+IScOjPsqcuTSTcym/xVLC0EN0lIxVsF3S50866JQopnUXFcrz+rhACpBoP7G2P
UbBB0jK8m/FMsumVPGi5qf1Xo+OWzgbvMH7//jUoKKe22hojFFDmS7DtK2QsRpp5x/SmZXwfwJN+
agM0l4bW+NTRXOq7GLYOZiWA0fzCfKwspyFwLuy8qZb/Q91hNkH0127SL8HogDPOPIJhvP+ti4bw
kX6JQO6w2dr2QeCOWl2Exq5/m7XMuJ6yQY6slLG15sWaGoVnAgg1fMx1YkWQE/OK6qYwTR8HSm7k
dK2XX/xbbPeEGF59mk3u9yg9hRAAzoPRe2KOFFXm5BH8L7vqGQUK/ZrQyyEvDIAP2mxcW3w2Sk7J
XqgNsq0fwHPAd1aJCJNWhZm+HEQjzbcEurXAqWYvh+zcqzSia1G9phxQMOJA6/U/l3/XJfpehWrF
FjEUn1K8wC1MAYVukTG4CHLAME+gopnF7WPr6AR5ZkoJhW/ncBwdsmrDrQRVqlvAo+nEQ17OkUUT
dRaXro7S+NNKHKRA0zSqb3pP69swmLSKtIQxxwXGAlC6Fv2DhINpCmIuSOpMqO8I3Eyia2RAx4BQ
h1BCN9Z4G+C0wHSL8kOixlr5Z9LJWOfl8GY/M5e8eMd5c6CbKHogoTf2G0OoSmz3eKcF4ludVERC
hxkGHvI+WeNpck1rzHTMK/JZOD7V8OkUov8LgU+MbBOby/jgYjGbgOAUPe+88oiPvs4f7+fWy4aQ
dMdgCO1e9gW45Kb8BIESR5szczMNInyk57kO4SC11c0UOQXceloeX0GcO+GBtfXPGoSP85NdwSs7
nDBEOKCcSqpr9cO9N2Ftsrod+J4jUNsYItlBiei4uk4GCykqB0kuWlHLbTuWIPn7T/Z0++VwIfSh
UO7YGvW/8eaOZOKuplqsnQJltyteA/s/NmdA72NfQrazw1RlshN5Nsix3fa9CMQCBgCQ1qdUflrM
/ZczVASSwjU4DY6+NTaArLSUGEnf9vqM9vrp6C+QILey5ROZxVmadxNloxU01zWCpwRnzBLfXmr4
9WaFij9Q1FkIJqM2IFI8HzW6Kk3mdCxCziICGTWxJNTX+bKYvxBaYEbEh9koCQWbm3rYqeaOIh4d
MIBb8DEXhRz3vR0/yqEI4VTObNbcM+S6/D1rbjzqDZWjwV5OF6C0UsHMcJELZlx0dPJ/wFQgAIDi
fodxh7JvOxePscz32lcHf4Wwrx+Or/v5lXYDHFvf4jo+sYpGCrlycwFwiE2l3i0OKBTHJOKtzJaV
2cc/xC/jHpnk06bkn/LotyxVPkslwogEP/Xp4T/9mSaR5GAixP9DWrZFq/hF/E1EUWoT6Oa4TH37
oBCYjAGTPLrQHPsAb6LOCD7BrMwGccwNHf3hVhZ72m1dAuXR3mKJ/MYv5WaycDv3uafJ2P0RIAC2
leeI6MXRy9hnrT5loMRr7w7l3s9pjajFHSU7ODQIO9mGZEr4IUcETtQlXicobYI60Z3iorVJ3UdE
js3ETYtDx5l1eEI0snlzw0x6eYE3pa2N/wDsgr5Sd7QqMXu1Rq0rsVxLzSBXPqOxtOYNrD1mK6lK
G6dIPNZwXosfys+ThxeVMV/XA7O43GyOlG7/g56d3AgswvecA/YZHDidaPDblbOwd1wgUcj4CcLV
kY6oYPWzUQGMi5nWTdPp9J4DlBq9uqkUdxwLHmR98vbDxTe+o6TZ132xrfKosWLOwhmP59Yw2ZhQ
Aud/2UCYHYC24B7xL1c6f7At7ApihKD5rBuIsXEaveU++l8gYveH/S/RnFWZmbgQeeE9OrdMzQku
UJcICGZmxUI5Z+79Yp4nI+3xIEfhY9ouJDnSRH5ScZNA3lq9WjbXULde23e/l78AR8fhWiDCrh7J
/oA6l9GGaNVIMmeLEaqzEFpjItpDAKiZf4xM5W32xjxvJPbd8sn/WXHXQsyeV0wKGN0SRS1yGUBH
HmH3/3RogfJh3SVmztn154gGjT+rfup+k7TcL7FzMcnhe9Psgt6oz7wi3Wtx2+aMIWD0nXQ8norq
y0elLHrD1mdQp1A3em05ybVoncDdipyyCyEr7wXp9zckJT0p1vIC2rHXanceMnlMgoAeW6LixGAS
RH933q3R/zIgmbQHUzxj+DJJ2iKL59XfF+JeqeYdDumQ6erIMMHA42vZy464JHaQopudknGOhQrd
Jkf+ObcOLo8LQZ0YvXkTDbySQy+6RPHqLB7UUM6MUeO63Yr91hgBbruQ48e/RzErEvjJFx/cf2hB
PCAbB/yyq2eFHFvdLRjKqHma8hGKHuG8EWeSk4IIUZ/eWJHzOrP+bjBVwRcbcHSx+4jy03Z5OV4E
vwZZY7p6oPx7ocNEFKxMfV7YV2fXmLK8NvJclQlg3iS+MdDeE2D/31DOJW/rUuMfUB2yUgajRpz7
VXVp6QVk+x79Rto2wy/p3CMkjBi2DB7UX2zxHjWssz5sWYkymA/qPSHaaFrDCcME849/dzEkqTIJ
RFFFMGuuM3LGy0KltdGHoMPFmbowkYjhzd6O4X73g1T98at6ZGdxWhePuYl6zCZdQb25Vd1z+rE5
85la6FA7ojDHmekma/aI2QZa/tIvHK8vV6P6daymcYTpUEWtb0ZzzonWsR39CP49abTlACTFjnbs
J0NBgoMfNH7gU0jqr2RXWsUH3des//3K3Xz8+S4TjRLwx4hfNsl3N5mGzZozyoGHVs5DNhbIpaSi
UucHYM4FuN6sKZRJi8M1MlyrX4nUScnQZwWjrS+SPkqfN2BeA9CIUwnHopMolPI7B3qnMN2PEyh4
vmGHurxyfdKOGhp3zaVC+fvV+N8/d/HHX5Ewluw3880v9GperaV+ffGg+XqjMfM0k4MqeONpkQxn
8UxFoWKyLcCs0L+niLmpe6SCgPMIu6rC1jUVFrciB7OupCEuuEYQqvMlzdJksdyqw8FPIy6VnBWI
wVxkXMCelUphB5WxhZtk9Aey7wsrAzLH/U8jlIk9YtGDC6f4d5A/EKeLPAz/UdSZ2jtdiyI4MML6
9vfnqK6+7b9jSgBjxX1jLxGiheleskofRRdEVt89HoQcvdrypnS2R/DNcr4mex0bLWfOTRKadCup
iPyx2i16EKdbKIPLzFyvhbR/rwyDK4O0r9ZPk8fF4LDttc0S0yjxgJ4Ok1AhLMfIww6tx9WdcHIe
Cna8Fi095qKtZ4CDDHnGfBjPcenxIqIeQr57JazzLEnKyHzStim/gUgEIJOPJIuZQy5G+j7XkV2i
S4wUifZYZPSljaFFjem3kyzLzKf5CS4TthwRncE/ux0Wwut2e/L7JTc8F0cAs0AA/LXyG2cdYfjQ
gMENEXP+jKGXgui2StvACXvIjgn/aoRiZ/O9NhXq27G+jjjbdddKtRa1gTmHlclKDUYHrZjW6wKs
BhS8R1+Bu6PIDUGVVnGHy6smPI6gAZgdyTOjjKKBskM+8HoqJ8ZL4lFECLyCbXcstD5xbDrZX4lx
mfO1H6iAK6AayK42wYCOMVFWcSwvPYjQJ3/Hjy8TTSGb+mU1PEwwNLRPy2m1+OajrYh/Jv3h7Bcu
61wR5RaAm9sZHaOcLCot42NIXtGf6Paa5iJGgGjysgaPzzILnbG71hOnplCC+mBSJ4EUF44AAnP3
JFSpEKztHlp7wBBjhj2sZkYqKJofJNrpFCLFLEGsKXbXMtUil4o00ij4mXKuazDmgmd9BfgCFpXp
BOh6umC4c39XRD0zZv7O/eT3aLpPIBhI56RYP91nklN2BfSq/WXKvEOkYUH/j/eqiBw3BwsWeRgp
9dJ2qx4v6LG2NX+ZaYBntRsoTmb4i+FtPdS1XwSoQB+VeI+JPEUek3Jch+N5TaeQvSEK8TlSoz3v
A0p3CdQbWajWRL8w84/P71AzLG2Z8a43nWGkRtCyATIfotQgVUsRCyfQ2yjMoaoymeRak43Afr1N
DooUryr55ECAdSp9iVvnBABUYjcMK0GaysZW1nmtquxXogW6IO8YgLTYGkWKOtCRbkh75D6VLmhU
X4V0QDt8blDwwbxKWGp3HrgZenvg/BBllHqImmbSdhcarLkIjrHpPr2Erg9gxcbOzaVn7bo25eKe
Zuq3f+6y63yPzQHpl2dMTlsc8bbt9vU24Dj0cJOFxnYs4bEZbPFNCkDSntAXhu5o3tp9aHKuvrd+
Wh3vR2HEJmD4Mh+H/E+2Gc+z21jO9j5SHr1mTv0ZgXvFWrrKCPRcMOH2+n6CBJVK5VPrePtkWfeL
3zxDwJeVD0DFsvEhYarbMjGZyJxk1wjZMgojTFJCkkqFBRgznNJvxSLUmCFc3DnidStKH/6Qdj/L
oFJGSWhiZcpaQIrPqyvPL0QzQI+Z9g0to9eWu38MEW0InKScrpMwwH0Z8ANf7YyUpdJRo371R9iE
POO4tlveCIiRpYQ3yA/xnhe+FW09yNs7sHd5QsySftAboDDcGXeuKD+5MrsuuBxYNDtf9v2/ZawH
31XZly8kcybhxpevwjPQpTGte86l9XmPgM+avDggscq/PUC2uHNRL1osSOaS8orOlUVZtSIodIF2
sF1SzodTRlqy8t+lLys2v92sw8Y4BW7frkn2AD+psPMYO6ro0YkKg7QnLP0m3RGDOHFGCzBdIBzs
qiYCLxb53qt6EKYkrRbclKNOoHuf5pjfRFPiVRZC1FeeZ6HZI5IXJiIzay664+xvAO17gaUSfEV0
HnkTErJLARpVDk+cPXSLyj7DkNFRrxHbieQFMRWqsrNba04qHQvYvgoXbhMhmx0F3pVG+i1mDnC9
TLY0SUm1mecDba56sp8Fh0Q5UStbWhGhRGScCZHr6FmsAW8d6tv+DOHIgoptWFZEXvZFTnYx8Zcp
dqBEQ9giP3HdkBP9J6RyoECiEo670LTC3ixzeIdvX6zu8TSpO71LnOIOWsRBpd+gZDtI86pBCMHP
ppehBRFZOehBGChmVSkB2Y4a5iQTC13ANv5EgSz0RpJOGvOjewFbwNrUiqUTG0iCt8h6R9YOuHk9
JG/r62q6eb2meLuZtcYM1TcDX8J19PSf7bs/kz01oF/kJ6ffyCCsZT3R4WlSMLlJB2a7v/j3R3WO
7xilGluQNursYh/6HGo5Cgx9GuEzdav/YLBOcvbiKXkghBWfKXqUULdSOa0N+Wc060F5lciwYIam
cjvphlvMofKjpf0IGtx+BmZPcUk2MlT9t7oq9ZkmB8EWlGHs76UjzlldETuWg/niZftbQ1ncJgmH
1vG5pExl6j9R3dI7RiMMqyqU/TWDnEPXHE0i15G+9zBm0I/eksbptSLBsvywkjetXmZv9uL5UYf9
J9aIoVAqSF3ShPesJpGdH9EWGzKNOzlx+ELzB7ASSyLIUHf7y/j8Zk70uBkcF3UTsr2vF/dyBF83
Mr3Z+842fLxX1emLz7FKRpRICbL3jjihZw9007Uw+yJghdmEY7+hCZysVVAgWIUZTYwf+AusbrLw
rMBZd2FXSrzBD4RfrvlwAP0F5gEsz0JPCnKLGMLVKqUAIJYFdRhP4wZO9QSyCtmo3O6J29KaIiIr
1Wkv3H0FVl3/pS2kSpaNUwnLSatSSlJ2IfChgI0MuQbFx4yhMUTxZkhsSwv4Aq2enRzX2aTaZPRj
/8yDd7eif5F55fyg+OWHs13cHQx9LPMuTcPAouU1L2JyYtDA7U7ixuaIFHB3u/NHwTOnOOPXvZ60
vdDj/+UKAcA4+VKTG8EDq2EwUCAYH4CPPZC25Qio8+0qaDSTdj8FXrpUc6crGcTk3vc71Lfk5bJq
Xu/8ud/nAn5rvmEbtvaJpnsyjpOkcvVe6NskZN3x7SeBLqZrdfat3KyA1Nb1/CySfuvsQYJRFJjE
3WV6qZkTQQpqqaTs81tdlu7kdsTZsZvmIm1ufXN+jjauVV04sWu6Ue38u5XapvI40QYaMuVQ48Gd
Nznbu8GXX+gaereNF7E5mMQhqKX+BA3CP0tmtM3ev/n1AyZU8M3eA8JgA5hLfHtjEML7jhmN2lUC
iBcx2ZDbYD6eBt+61Ce4b3MLX+9C3+Wh9MjkLVtS/wFV6jvZdiSS48+vUrLksTZ+LYyM6zHjOaqS
Nd3YSOZPnZRVrTjBLM5+ee+tKuG1fL1GJRmnaKSpQVsOyxHNSAELoIaxdtoxO3ldBxdzNBQkyVRW
P5GRVBG2W2W1ja+LqiuX5n+mpO2b1f9KgmBO8U89O8CRVAyPoZ1rmDfcVQ777dU7S5ZyiQK7UfJh
zmoeWArsu6iZFAusnzqQRxec4fy6tnKwMYP4FoChyY1F7ycYdPPERqLSoEselYe1UuGtjPngZQu1
JrHmRpqqVxfV+pCCNHwwEm/mdxI1NqmBJCSFFgx0tWzQfrGmuCwzjw3gULeEv0DgLd2YC96wVI5z
q0XZ/RDfhnKu9W0gjVy8VyrGV55ruVjPdarjrCQDQCnbJufC/+/XbohcY5QoIu028J+ivEfB1IPm
SJVrtX0BaqAF5PyxjzXK5sjqpFeknQOcMbKWdymAy2UukqHmT8RxYqPIUz/ZW/g24XwuDFpGbOz0
3YeZ1My92rHlmeFDjvSD8EQmBfj/I+i04BgOm9NI6uOJi7V5Ql+8Kx7LCFeld+8FZp0635rkdZ52
ZXq4gNf5wZgA13ylaCfEOYadIcj3mStaY12uMa/JVV+k8Ijtdjruhxh7CL9fo940TOVIFw9DROz1
UzglNNgPdoYe22xJvMYzH7FU89G+nFzMrtLJug2wkjqRlLj+ynf7kAMu+UvJfoofTHgzY7B7NWpl
UpduEi25wgj5J9xJngmcxpKrNtZI36CR3/GwZxmgKQlm3DM695hD//lvv610y0I3tFLaewD7FtSX
+I10F9nnyERKrLvGcFoxScaKsRh1xlc8wauCiF80PvFlPROnZkccfiKZSqx8/wR23oUdQaa7IJdi
AKVstN7ICARiDwxjE3r1RYKfriZ9lDViAAJKXpO31ubsT+jduxAm5PRuQsYp3WkHciOUh0xzm6mt
XIwk697+FniM3NOxOEuILDVDjCejofBAJwViwDaQChYGM8ioI1Ti7VG/Y41G5ozoTNsDKL8CoPx8
8aC6YtGAwdo++oEcijiWDGYTb6cnMh0cIDXoR4XF477tfVr13FFEWC0VFiQNKyAGNgIv/dY2ahzn
kHCLmKQOTr8fC/lvI/o8hgr6zCOojHYtAy6BchDxoCUpJVVHKIj+G6L9dIykCGU//Rx85W0YlR0S
jP2BYI02G/tFYZTjBxqot2y1f8+95it655E53vxG7lIl74zhdT5XFZ8vwDKgb85rSF/p4Cq1YnM+
jCDwOhqpBNgf2FO0n8Nrll5hjS3Q4g+Dsh/TwZAoSwmt7kxGa/rYwkECdaXxhBVtXubq8rFWb8xk
aSQf5oz/Y5eiC5qkl7PEc+ha2fwR9a4upIPPbhJclghqVevvXWluda70iJ9IYQAswbd0MBNzZoOP
8hDcALAnlIPso1ZsY+NYJJMr72CGg8POZBtTiyNkUr6U0Ft11DoeL6VU5jP+LZtwJZuIRfJdqEkg
H37C6B2n4f6FKMGHR+mi6baIP8Vtx0sy3XCHEv6s3zHwEQucKLiO7QGmn4bm4853h+btNTFfjaqw
fBzSES3SIcrRMgjYwNiBz3ZCQnbBjFKQBzuO2MlTYGRN+0g9hjORCGIGAxkC1mQ/hG35FizOAIKH
z1SmpbgsaAxw9gKeOyuvQHCw3u6es3xfvJDk1RLUEAEL1G9n53/tKwCLkfbPLWxN1xZS1vPOaxL8
ObGFECK+ZEU+53Tac94ARSDW7TtT7OdKaCzQePitLmUqWyCiw2X7V5qvm/np+g72sitqE8NG0f/d
WMljmSAShFtVPJclA1o+z78zs0lUHObhU1QvrOw0iJQoaJbb8/w5dnAzGPl0PxTLy7PCVUi4ErQT
4xf5ZvRYgQqXuBO4WlxwmWl4AojVoZRPLUOwc3bhgcdBm80CW04xssYWGuiq8eAo/99vNo2muaN6
rDGhUfwieqQuIDFzzN8hj4aKBHhhzdZZ3vZzA1s1ZTi93bhx5qtqv0Ts/pdnHhkYVG5cqOkWz04Y
l/uzPclVsSx+q93k4Vw/7EwH0plIuXDdGRbx9QGCDbnCgpvHCjR4UCz1+A/OmHqhRnLj5KxrhobQ
vk7xr87a/7XvVMNpauEWRTgbZqi+V8CXV1CWxT7NyJMDDoyhfdS9ZpstDau9pipzRmbvg7kA/GjS
YjKMOsTqLIis1S3UzDeF4zNQXMBTycpZWgs0K6EkSCDS3AYO876UTlmN0hulny70HvtfR+b4XH6h
fmR7QVluppDDZsSbkMzOk4xPql7F79bg3U4YdGxT9SXNmyuHR2nJ6ciHtCJyst6FBHVTIoVq0AE7
7zwsSn/kFD36oFw9Ymmc4oEWHjX6dR/aXivJlZYhpz+QF4o6swCy5z7Xh+IExMCzScTmlJouPVxp
BOAvVefoAnkJR7Ksqd8et7mSvvnbbXagDKAgHhQVODFriK+lM05LzLVvkd7fnmOHovEdnTTJp+Vz
BjNHVbhLdC67dwgVmiL2/O3xXbZAxinn7BgiFvUv7VpeObeZEohkQzpJoK2A5ZtWZXzjx86F9bca
rsBgF9z282gzUacCdWq0Khn31Twm74R7wpOUNfL8wUzUHxxzSGyK549mkuukU0boqHRtno51haiG
+2amF/04FN3zDRt8P7JzBGERmhiJCxQDFVxUhOHMVuexbDTU3Oo11xDrmHMRnGm4eWF8GbpHisPZ
4CxGxsl8S3y1AVsMZncEg4Q4lRJfBSFUo1WUKA0UroOaUFcTDBNJm7QQlekZ5oHhkVuJ014CxxEF
MI8jEjWgkCzcql81F/zBrhXdFITsLuzNjTSnzJJZIaq9odwAcGi5VUOxS/WL9uA5DERXAFg8SKEY
X/UgFCvUQCXsKHfKK5GF3kxdiN2B22RDMppg2htdRNXgshzXGt801W6QV96gqa0IdJTReZqOwUk9
w0xDqomoMa3RLbgvQf9FFNgeQ0wBSGqMWxoa0kowDLsgrrXwHzinTbJ2irZ/9GuQSz4wAQCb0qlj
zf+skqW2fp+xwZvK/wN0pRVP7xtEcC8nVj3atFghkRlA3b5wKVmwln/vwKGFdwkGLrkn2o+VddoB
RNeyHm4ks/Du3NniVmzBT1f02qxkusxtK+Bm2QPNQJdBXH8Vv6xBYSdhnIe6q3mSLQKYQi7qfYPp
paPZFSshUPp8Y/zPxtOWRZIra0rYagSNJ//11FlDdnx2mJTUaaxtZuuED2H+jOd61fpvqJB9gyOE
iEbLTB8kS/+SC+3DXx8vkk3SniXOlsBIklLbHP4kbZJBbv+nn1ZFZKlMbTq2Snif0awsu8SMYsX4
wSrQ7YMdZdH24hpJl3zjjukjzktXDru/ejjfqBKr6mdy3Y2F9uKhUAgwK09qimib6RzljnInObaW
USwQfpfz3/S365o1qKXTp6nhfl2FLtlaai7kRH5Zgtikh0cPUsHbZKkjh0ynwY0PqBOJ8x6Xv2Ht
rWsieaNAJ7W5F8b55TRq3Uh4kEX02R0EjW2gV3Zb8VVbTiudB+pNZ4B+lSfHKRFRQPiAdxS2X1K+
aegqiDz9zoZ/u+sdHsmEMFJ5uVBybQXiDTeuL1VZIw9g97kzN8pQt6KfCUay9SKGQyHc7fdvQ8XV
p/wIEV2Fj24eycUocT77Y1cW/6RGZs5G9/wOWiHZXyLq4xzVz6nMEHvSX4KAOL2hZcQIW5wlkNnb
wqz/d+aZTZ9kOai0U+4tIdCkEyV7b9KnEWpJc7BUV8PuJ/N7AABIYd9XwKKILaa64BBRgh0urDyD
I+2GNneKJJdfjaLNdsxfPrTl08b80V9EHaSmV1xc1bmzfL5oZ1i1u1W4o71OqlVFlFC7CoaPLzYV
lLBzwHXnsywEGPlHOaQNRLO1wEpXrYog/XUkILVOMjxstD2d2oYnPfjzs7oVby9jB3QVc4Lj1hoG
AgH68oMJKl6nmngj7HAfUuz2w6aeDFKNSmdelY+ruaHA5tJbtqx5gHOzcSjLO+FBgN+YzmwqfdMJ
irJ5gEOzvSTLVe7koWVbcjRASpcuXl0h4QOGKKePnoKLhJgGUzsE6VGVTQl0deOlSQW5AJZr5kjh
pwNT6Usd4j6J9C06ROC/oserYFY8qj66bZ6dGeZuqZiecdfxsAuR61xm9D75ZZtvti8bTUh5aFcP
3BlRtqzGXhJ9xf44DMkasEEi25kOJIrTj6CwS02pj9oJnyd5S9GWrtU2diKVIY5WLyDukxHNbHRL
J1MyNusu4FKw2NLfyiFV7oGQVmJL/GoAgV+6GGt5NrOc1KaThBv4Gvb1gNnLt3paOV2ZXVvJBFtR
7xeyxRoUGFn3dCRaoOadyiEe7Sau4PWmz3jRh+yzLvKT7/iIxrD0QFbScU95/CocU8CuZIyFUXtM
j1WVYj2QVNqMhJwi49G9Do7TbW4Np2ERxR6xkvjwEx/nCZtz9A91sVQCCKlNpMd6C/fhOqWUXd8I
bpN64lmhAVcZy6MpGgEqBzi0jg8AoqaEAGoybe4K5wFBXCI3PsYZ6evhXhHdU5seFhQZwA5ADHCo
J6CkJa1A9YLxdXYu0REV/29vWk+WGgUpGCpff2UqgRmL7q10Jf0R1SN/sz3K02ux+tc+9xiROyXk
DVNvjwBMoPuQvoCVT8E3xtxEKsjW01zoa3icvjEI1BvFk8myK+l9J6BKAOmxoiPNCth13pcSi6ZT
C/Q+GC44rCIo/QACBAnaexMjK1qVCb6/UhNIvplLOwQeXkQ3HHBWFGdTZ2Fn2bOylkAGCN7Qp7V+
6PsUVSFaThnUzSzf3IovkpWl1QB3wwE1N+BaYXvyZB8ATziH8BqywYvfSLHuaWVS/v+ZP/JH7Dvc
H9F3H0HZ4+QC/0/cuUHzyCjKtPJhnp74w/FFeuO9JPZkbCozykDIV5eeRYbOul9uQdzBJAKwCarA
3x0Mwf22mG+NDjzF89Ns//uTM1yN/WECed20bGeP39TzBg24au7sBe2/eDLPhWcX/tIyWdjsxacD
GFpB4XjKmXkoq1GF29u8ciPHFTOVmCeYHhuT0qUfoG1w5u/c/AvfrEmu9zgrRcl2BzyvzMnclh+L
BMLqXMddRNc4uaK2UCIGrkAjimhwTfZ1Z5uX8ZKtl6E6MyfkerwRvAHz8+R0Are6xQXJYAlRebI1
sGsJhqP9kDL/pHy+nHCnQ3inRk7xbR+8s6jOKCfHQ1vxCdDUMJC3dlzEVmzYnYg5c0f3luQjWB6U
krCDdy8W52SilgVyPuXVwA+aqxC0sH5mBDnxLafJhFP7o1frS/yUNdnmjkvjXSWxj4J/GLIc4z8I
rsOplwmw2wJRpyQByz3xONc5f7FJtGbB2F/hbHF/Ovco+FKzwP9tMtQk2D2wIlyKKXyiYZWp9qvC
wPAGPY1ouVH3vR3F1xLYcGvLdl5LCtU1ZxEdvZj+CJWA+Q1ipfEE3ZewxrBzz6EWDw6wVt6vi/F0
xp7238vH2rmmtA82klC23SBxPUc8Rlui/0VchyCZcT+AiBDu9HxPemFx28mxPyuKyJGEgxb95MQa
J167BckhZ1GrxLxzSlN9eCmeqlKlu37gyDYY2CSRWqkCRVXS0LMzPAgc4WYdZgp3xy3kc+4n0eKA
7Kwk9RNgdA1asY5fct6dKaDvKr+M2UT0ZDMhxBp23aGsgLss56D1EqyTkqUy0mwnQoIGo1w+Sj3C
PKH8LwwOD5DyyCJVnPO86Aq0R5i31Q8jif0jG1lLRyPDOdDIKw7mDidZs45PbREo93uqZAVGb/SJ
lAXU1YHYchWzmPkW2aOtGIk9YNQemrSCWOx2BJAdJ6eyhnmRqbYHUKMidH0NndqipKyPHpBqP2Za
5TwmokWvlLQUXcdnwJJCxpqahoUEPQhrUG16pWJG/cRgmxMIm/IIqbNFGFEOCmq5nY58z99LWVHp
aBurFQwfjY3m/jbGdU8qjthWyyK/3WotTTO02kWU/iKpvY5MPOTqXz85CDgR49GKc2bAx9y0aaMX
F1CgVgq9WJxn5wGzGMFav+ucoQSZ/Y0bmA9Oz01OXO+zAHFcKQVr3oMPOfmM3FNFEBMyamKf2pEC
GPUDLEENU4yLwTv2IqdxWFBY+pFXEn27tMw8XX03vjDQdSxFeandHU/mBUS37BG8tYlijQdZ5Pw6
Mz7gvJ21QXdoBTvd/kvtMkw+KjygW5wfuB2FYJW9ZWsLoS9AMeubB0ke0iFn5Y8SO99OHKqbqLVv
yAhUlkg6C1MY/Gapa6gAo8swuN5Ht6Ygh5BiVRP7z6WVWVLhZB7pcyxLDP3cWtw18106cTA0s8MJ
rDQoXGh+1F02lqOLM7GZxeIkK7pXJPYGeAZxfUGvvTisxZoy1bMXILJYTCFa14fo9gDd1W23oETU
/6rSQWmHEUccGMlh+ONS24fyW1GsvS2+u+JHXsQ8PzYfkNU2mQqozH/IpzlhpOByfbL606zAKtRj
fD6h+yxJob9SdVYHwtfyYJOGdTl8ybnRCI4XPX/KBxQXeKeAfhVzNFIul4pgWWrBpSEBReaZdhBO
sYEaz/F1wyeEYheVP/X4UoY9auSLcevBHBMCF2ecbZxVw2hXpyZ/xUYIT5AwXh5hgp51c0juvYHz
5duCXvON/6Fb4bEXy+F1su+wNi7XdujsoDPeM31kWE64Qy7vjwOXl00qobPJqkEo65jjXo/jv15w
+MxZN2WyyG23Xf+74G7d2Zn9CtT3PebsHc81ELmV1sHZ3ceBAPNNtWeqUll2u+yqcmbY01vlCgT1
sVGRVtyCd9BDkHnrn0wGW5R75ffzjt8NCjA+b0pgeckOhvaxTJ8P9K/S7Cs4KUwk9A/WjCohiOHs
XeKrjREOnRtE6FC60ReKy+K2uU87BBDsH848yRAJDleR4DTSdEhlXd8z43zMJCdaN4xSl46fIavS
RGXtY3GnTIo0ALkeWMDNH6b2fIVtzxzXxkCE8xJpii039u9dtJzVabBqm9jlfWV1yvJoBweIcXLJ
hY6e6GY8CfSntI6o2tX+p+1yhbo4HWCCtw46U4vjmdNkFU6zPRnj5R3eAOhGRfATqOLEuMFxrLWA
fxG3tE6/CFCQZZ5FU7lFpJP6y0kVRbdODc+UbblF+LiByQ/qAYVTGAS7ydXkeSM3ym90QqofV1Kn
rcoR7T3JTZIwSpR1Pv63o6RLU8HWFKOZuEkL4MAfaRQOa4vOw7rSW8o78aPRtgErMPJL1LlJGwF1
+PKA5rBJE4medbwah5/6XSEgXPKaRXOjycr6NBPBQvokVcTNwfBDLVQEFdK8iIqpjhWxNW/45ar5
6TXg4yIlmEp1pM2cSe8dkqOxxiqaGm9CHngvQQhD9iMGnUPqtAciZanGwH2mavISBTsjL0V0QR4F
mP6MNpZ/d0RZpBVdk+1A99k4Pe3EAFZ/UsYIf2GjkciifV3muLIrrzjh8wIY41TFrXi5xlDm6Bk4
Lt4yKuTprKByQ2vjPXLqSFAm1aF+FlxwoORO4qeaYRBZb2WqI2kQe87ZeA4xxSYHa8fdr5Xk5+kF
2qEinIP3DopVGGf1NZv4UvOfnEzjrFIXbPuI+OzUCEZIx9FDOOsa+AYhbEmicYicwnZtwIHvCQc9
aiESs2FmaenUfefZTPZMwvc3wUidYcZgL9aP0Z/7NenciEwUBnJyaPKplmDlS4hb01ADmp2DcVq0
cGjkKpFKIFkI107Sgp9c1ygECsxVn0vd/YIgNSx4vDYPoW/sQoIYHU8gmBIzdnrav4scfAPaO9pi
3Ia4fPnoZmamLba1HD/1QTKtuHNkZYrCcZRXtwFT46pmPgt47eq+mOXeYj8AwZd3ASrGwnMgLxX4
mnKmf+jX+ubZJ7290ZrYfawQWpykbKy+R031OQw/8uW2m43datUzYrXRrmLUB/IdSMOpPbY4FDx7
8YHNYGZyszPOcnIAfmC/pQLO4WnSsAbFMGYOEyYdLqjcjUuju9PfEZmPJIQucgTHgbvFu/BgR0Do
8kLD58LPd0Pm7jnJPJWoAAKUGNAysjSUqBXUfxdiEO+bAyS0/0COqrM3/xmwWeiwTDC60q10DCA0
kOMWhTEDacS4fsKA1CeJfp7nmD9x440tCNBjxvK/aoiQESsFj77NJXPmKhZOLnmAa7D9rhHV/PDo
OoBNKrdDS6KAk/6PIbNNQiUvyjM1DM99WVOtd79slg8/yhs/4AoIk3HQ0YGaR8uAJb//6tQkpVXO
Ka8iS9MB51pyLIp/rD5CqnN57f/5Pf/GPAfg6IJejTy1OReqU/YnHKlumWSAo/KFPFUMsb9ZZD/7
s4gGMjsPfr1EkvWjdmdZof8lx827KtIVRjGyMaYfxNPEjFspfbYMIaTterdZ40wttkNm24o55oj3
yHSt3+5KF/xtJLn4J9J4sLblJucQS7lZmoWYBD+ZpNmnHweBHOrp+hfvhGdcnuSz4wXSVwUmWZbB
0/t7mjkHEq5PKI5RFLPOGeHBW8TeXQ5KtGiR4hIzvYDsAMdME6xWl0ciDyidkd/+3ru/pfhScZ4N
jNlkT76TDGRe9qiKrB8ZhC6AQWlyfIEA22AxE1TgbjXzga5tG/54gDHRV6ppc7zfU5LQrW1aVzpy
amZD/FKB4aqY7mSn5rL/ySvuc0b71G6wEqlQBNDCoqgJUIJLjyyfKHEmSpfsZgLEXKFbU9HVVeZv
wFFbq+zcWhvhu9K2rBwTCypjZIcqvtB+h+SAfPyITCSL/4gog5nePiy4JddjQZalJFDNJhczEqwq
nY10C7Q8BiHG6lcwYzH/n+xUygglic4S+dsSppunv1ptiXpDWvP2In14yTG6KYTtVrioIx6pEDMN
soIxet9gg07D9wfD80HSlGFvWhqJsHwcwKUOq85ABZLa/9s2tAAd1ngOWCvL7ZOkIc0MDliHX2ZE
XPEhyPDYpO+vPrpq6Zo0ve/ZTL/QoKvoS1wv9z7Uz4YU5dcGt8F031sQ3hK4TW52qFFEhwI+mRwB
ZNSAxEz5oRbpiv2mMBKuK5VQZFWtkFkT2m0Ka8fKk6EPL/sFu/bJE0Y4v9ZIjCzcggBU4XtjQPUh
6e391YcLevxJAMC1vsMoCieeg1yiZL+jCystSkND3+V1+Sa3/HL4Es6/dfjMw1mYadnbSpX4ff3P
5Tg3ORDmrWf2BDPUKiD9gV+mMtr6xdTW46SJDvpbtjtyDdAQuLPOboQ8dub0Kp184bWGHimUNhVb
7oEwsup3BKtp8XaEUsJoG56zQbdQ6VEMlKYkXMEiCQ30k4Ju5QPb1d0zoIwHftfQfrdX92JHLkkC
/ZqTwgJ4DAOZw2MxTOe/smJPFPDe9bbrx6sn2af6lzd5Jjhc2k1JXNIBFhOgyPiiYkLjBWQhm59m
hE9q8D5rhQMVXS/AFgoD5sU2cDt+KxtZ37C4WOW7Y21I7YRNmuct07oTVEvYYGYamQbsVu4jKfij
VfFHCkqK+pbEGcYSE7uOJXxuzCkbNty84/812g6O0sriJQbIvSIc3yVGRTUtNuZb6UFX7hNYtwsY
vswpYsfbPLC3DXXBHNdwFvs6760eBu4eoc2IUeMmixijHFwUCsWS/2XVB+tsaypwI3Zl9w5zfviZ
6ODQUVAomZ9dadhEtgx9f4HV+w57X7h5XJC+xc3vTZbFBlXs5VbTbRBJTzkz0s54vedQUam8pIvv
h2ADrhftGfqAH55mRu72D/mQgWpPIS1QFLax9SvrWuL6a9xpA8uQbqdO8eUaF3HBOzSXXSWAokQb
y3xoVjGFuTnRVpY1u3xQAt4Vj+3ldIE7O1Om72FMbCZMdgpBP8i6xDYopoBNT95JIfbjAitjG+ol
ernj9I89lXeXFYyMn/eJGKzVSHdvBnYryyymm+Df/LcKQPZudTFq/bgqhPwAGdkx8IMIlQ2RjVOu
8hQW9JzFOfygFVuGXATvK+6YEmLUabISs328OIW184DvsVEljlSkGI7DD30PzmNV+0eWYj/AW9EN
5eHUOIMnfc6B6I7gU7yMi0oAUPnENsO881ChRXzfprmgES6xC5haUFvvD6Zgle43a0k/LlmhB0IE
B7YtkMHEwmgqLFafUcX7pVAd7amdchAVW+h+jBVVaL0IWTpx8ZLwq0qfpEWq5OsqT99ZdRTPf1p5
CvcGsul/xFPT64A+Cvkz6X8CKNE0dZD5nr+s1Gdm4ezhoQvgpQmxJzYkQhdzenF6rWQi1z/kVcaU
OkG88e76kSrm0+c3KuPF55y8vlPFMGe/NTCYOeHuXdrTcZ5Fe147Bi3nEx2A6e915EX7ByIf7ckN
uTEKEZMHjOeaSHXAo+kA8WbAozO05jPYU+YHGhV7cRdmLGBUDZagv1L4i1eKJk3bGVwalkU4XZpq
MjvftpqeXaPNmsmRXQVRP1zbV7Og3NkeIJc0G+80hZKQMuGgLByUtKys4DWycVx3MrL2uZbV6VFd
W60/cJRo1uNDjuR3SbgZkiCPNTqKbwq9SZKL2ca1ME456HIRnIDeP2jkEPxXejdoSEUIhg6hGRNZ
wZOXhzMI0ia/UQnwGa/BF8oqiZsIMRWaCbNGIsdqRQeyd4q1ur5pU8azpZJKrYFZR6tMte9O92Qo
IqDHWjXO74GrMr1bumgdn4bzOYowjnbkH/1gIaL0YvBuDIB4+ArWk5nIuwK3xwhPTYVRHmERgNiQ
+I+RYddDIo03EmIUkXZ/zOS1c/MkxI602glTBorFs/xSphYRtJYfLADzgSuwND7GF1kIatUwyT1R
gKNDryPEuksj+zqpiXdDcpUpzY4VtTu5i6hE9DSwbc1xkgNWqcNjWoF5xfGkRsSBdZwIomR4yvjS
bmiVq/DNQZRh8ki8uF16mirpwuCPlOCijhANlFlRCNdUx4vFuyr8aRUlYo2i1R8ynCWYdCMkKXxr
2LEiKDxrLctarIgY/V96HFUNu0AUo4BD+J0T97HAt8fm3Lri26XECHIaL+l7gjAU7SG0QHMBtkIE
q0Eu4RP8Ox2eZxwu5BlnTw1XhjCKvLgUxrbwwrKTNeajgPGLjfbgMMMhuls1e9pDP5W4BL2Ux+Zj
NffqyyCDYftX1JhWRO6tDMb/Yp0dtILSyjiI1E2yN5oGKw73+QS+rFmEgt6BtZ31NT4DepneQsTi
oBG1hdJIcaAUWB2MvR9tQVq0noF+e+m/tcns8CbjCLYMytMAHeHC7S9iaesA7Cz8gEu1qOrSE2Vf
Ek0coZwM6cCck709i/44efJjY4w/gkRWbZ1H4SJJm1EXrG9tV1EcGYHm00S2NnS6Z+huEThMhkRT
d+KQ4cyNiulDBRYwIE6VttKn9OsQcaZQcN7B7ss0F+cPqVvB/bpTjd/4KRAXcvDZv/TRmU9R43Kv
ckDHorbp4UL40kL0tBiLA7O1tuYiPHkA8yuRihZx6KafNBwqJsCoHLJyDnzguKOhFQ5L2nWlrUQZ
C9i+Y2ifaWOVCUWNBCMz0iKwpC6UC0AkPNLp5qI8lRvVKAj1zaRcGzm4fUiJhgdgJunq93Ns0c54
bfEa/o5N7oczx5r5VFVOyBmSmVOsBPpBuSYRCsDvzM2H8nzy/oLNfL1+5qXMAD+ifevf+7Ol4sdG
bvgSb4PxfCtKcP4ViE8p2LzJKxN6h0EPyCDrhD25eRykN20f3KzZbUa5XQO3aoAZq9va2FkbNQft
HTaw/dhh5jhaKkH8zruQOz5vHyiBtyRy2dvUtGztbcijHVQ+2CrHEc90xAQmhLKcxVczA+7weH+V
m5xuEX/YD82LDkfqPpwlnda+uoH1jm3BRrPg2WSfyyPkD6/p6aGLdKCPyEV4XYDNCOeTMNeO8l8v
7O2Y+KjPcp9in8U6tXAepFPM4tzZFqkU0aC4AYQ56QHl80GaNzeDEDzJGNa5r1cXOoTMFLbBWtlY
/erpRDBQGe3gIY2AtUKrJAExPjoZwpoSyEHAI2h57JvhXbxwoRGiQQc4qg3l/YIQnuEbl3i7mRwV
9Ei/I7ySHtSXUG0+W4MYk5waJVYFTB8B9rxPm9mSGMFoi0YRj5ilFfqOdBfFb3E/Xl9yV+I9ZTp3
VGMKxZtOIKEbbeqHXLS9XSFazEL5L43XD5B/8629KQ/uFt5jzC0vLcFqLS9JFnFrbzwfw2m+t1FI
wAtKuAd79c5smjFhqO5qKPum3FA2kYUCVZkq4e0Q1keYfNhnAXxM023o2rlGgM0eYfDp4kdfxbTn
V3Fw1fymSQj161cyGYiwC35MjVEjs+FDCyUYLkJoSE7+I5qlzo4Y+1C0WQCUonbuTn3+Cp1PNs1v
5yCPu8hZCIPaPAL99xS+6r4eiCXLIt92nOm6s9V44HRNFyYXP33DBlo4Cyhe7M+pCJIs6ZNB07mu
HFgZok+/yxzKrLlQl0Gp8WwVclm41xh+qcaoCTEN7b9sXOV/V6l/LuQ/u9TfXYm66EebO6GK9SQV
ciZm3CNxdlup4qmg4mfDIoFYo0VyIgbqLQ9SOxiWtwF3myT3+BzkyQlChGRsGAXFsciEGxkjuUlm
ZoZUMd/brGT1TfTRbngrNWHxEkxFfDhYt6hkG3uodROlACMeO7M78Q79o9caQLUVZvJoiR2vs4KU
WuZz0P7Qq/1lUdaa1BHH57fBQ4NhPNqDW8F5bv1teBWnaRHH0C4YJR8Tv6IUh090xPyUQCuO0lBH
V8WrNn41VvsQsoQCpgmttTyV4iQwTejQczwGaB/Zc5tMpdBAMdWw/oV/y8SDMvyWivaWSwrdhW23
SWmUJc7qvDXG9POOrQTNcbosOoCth//dINWLF1KEn3BUflnh/Tbp1G9Z7Gqn0LH65mYJmpBQHVCO
K4ly+wBOYHlMWcupjUT0vi1qjYVs+McGuq8qEqmHGfUCRi5JPbJzTPs4D4L8rZfGrAzhW8981Yhd
M/lr+HnTtb8vkXhNylzVSCwJbsy3/nPubKGvcG8WunOFw+J1Ca8YWNtrjSBruCdKW9VFzkSo1Gbd
IJ6UlLjhzRvm3F5zThP81UYE3Rh6I1guqfNwYnW1xGy99K357EYXr06UPTPTQvl6PFGfAmD1pt/J
h/Dy7C03KNcyAPUEYRXHu6I8dDt5Rrl7MWH/QyO3t9QaKXC0/nbMo7tuwbVsitRD/At99rSO1bCP
nscsMeNNN15jNttdLC27U0sR0rlqSRuqv/SSgMdjIee0O6XF5O9Ejl7wT5VuX/PvTgVAxERc3yFd
1HD+XUTtTNPGCf7BLiBLpBfKk/zmkZ52hvm2BA2J5C598lnoD74E3ECCBoOzJehLE3u+rE+mC14P
GGYUR6c6pPmE5w/v7kT4RtcGJkiRmCNH8TFJOyDCXYLQGxwhrQ/xHdeCYSYroKWylvMZg6cWGWNW
22v0wwRlXaHIcKsx0VzxR8VxX4CjQ2CACP4tt3gtkTjNxjl7UAPBzsRrV72s0Q7BvKwc6q5vue1m
0NXhFStZiJ+7St9A0l22u0e3OH8fWKuclJcMkg4uB5vTRT03YWavQ7hSCqShC1qDCjJeFr1ZyLDg
jMD16P3KLC7dQTMAoM7TmUmlrMYi2iQAgOccQDQU++mfRWMM9js2YagRnxkQWygFFMGYbEChqIez
o+DgmN8e86hi5HHBYdrAkGQrZxCLbomTX0GEeuxi+jPtpYs2uvN4X6gxbQeM0uinSXGLpEhgjpn2
wh+lAmxJ/v6f1cnDcC2KRhbpsElbcHKsd3pFypNfzEYNxbwh9/5w4rcxzewIGjS7/Xc1EzY8j4TW
YWs8gbh6sgTnQ525wxP9iHNX0H0EscngCg8sIS1FDLHJlb8eybgXjr9/lEhx3lwFiMVQQXGpAW6Y
nTt9ZDY/lhXXqaKH0hdm2nELn0Ok4EiVAg/MyIlBRSO5Y0FPOAJsHQfabbm0TBttzZASKpt6zXUN
pZtKypWmc8KhUHzlqLvfYau/Y0iAXqz7t0BsF9+HjSbtt4hzvLMKo7+jN7QWjzSHsVerVJIB9O6G
B2i42wyjkm1pMyFx2IpVR+KYMk84ilvtMze6N9MyiL15O01xB1A3jsoAyvCvMEpo+XbFwTt6GST2
kLn91W5/rT44idBNbhjHTZetn2FJoK6vZzPpI4wEahL+Mxyt2ulgk6RNWvOyVzilo/NDwBoQD9Ep
UacjIQUA7fSvyiwrYJ8wCFpoZOwdNR+S7ooZCEjtE6aRsgB2qj3/Tgvu8/+zl4/D+Sr8YNkDK4RF
1G+BfylACmVSrdgxq3bD3PqO7xZ+IBCMfQkeNn88Meeui0g9L553xA0XXr7yu6WuXAKAqOWcTT2W
ek8fR2j776wcXLowIg3v1OiWjjm9fTewEYpCzz5G2Cup4N9AcNpdegThYSJbcwnAEwvBoKhGdGLA
5GInBA6vFFnlckZd9OSkqF5pyuyPtla9mAM3K0DYaQKCIIgciJW4S5ONTr4pOmvsCCl1qmdiQsbg
OGXIwAhKA6hRXulVoxybSfw1YVZqxjpl8E9VWJO1+TO4O5El4qOef1Gzsj9H/lwFF36iQuVp53Tu
k5RoACwZ9b8TLHIbrqF0sp9VNFXTV4sW5AEu0n+zsFNPed+CqJ6dPfNSBGY3ke7yCVKmFxirhJZ1
fJNIIE2Fd+tDOAY1mwa8U6IdjeI6PlT4M85isbifNiQbgEbf6Ba8nM3eiRn0U5/gbksx9HBPoJff
Ktou73b5j/txzHVX3kHJWyLB8hf+s95C2FxMhCTkk8UMnPf1UuyD8ArFWUXgh0tJOJ/y6tzCVL6G
tn3o72Hez/IE5bTmrAL7ZPo1oN20eEuQvEUAOjwyP5lujML9G9GOMeGJZAbNUQiRIUgAYRd1K2mU
DFvv5B1CjLAjUDvMxc6QK0e7vHsruyQfl0Frhdjtq7T+qUI+JHG/f/V7D3fjxixae4cNlsxBf06C
oKjw7VFzpwDAkJQYl3lePS1Sm7kLSDuyHVi53B9KDR6LU2AWgPFL4zOMxzSRv+7xGpxMNGckYZiR
eXsC5zpx0f2Bp5UYLmpe7d1uOx74aZN+p57MCoNZNkhXyLYskxyhQCe1oYwcKfzxzRjb2JIMJCcd
3Ogr4AjILD7Q8m+GrvwcPzWH+atkNcMXK9HaeHBGQ2Y1udGsXYcPuyK4gpGZExzO9sCI788NU53m
JUrlJ0rCIrw/0Jn3o/n5qu6ki87CTVR0jkoBEJVkYgLkLzmKGPTIiNaO9mGy9I776ixPinWlHXjh
TYzT1+8XXT5x/Jph3J5nArWpyHnyp7vpmvrKYzkayBfuRF+ocnjVmOTPziED4xWoRICansD/3/13
ZhNvFZwHEJvrK9pFGH/6sTqN4CjiCD+MUB+qqvoJljg67cUZ19y4/wXlyK0CBEi8QcW2XmhmkYsT
VoXxenn9BWpe/lKhOM5FKI3+dEBLB3/l7NWCLbCC+Mo7XSkC2kTMZ0v1SY3c5M2b+skTA4sF5hO/
sGw4Hc7ONCzgs+B8lSiexgMg+uvxp3NIRjDDvCSVhEb8cKE72wmf1Jwj58Iwr00evakku+IspEwd
X0Qcb4XGMaNUbZJiYi4SytfuJh0h1qqANDmfPs62GGr+zUNN087b194KzuUHnmgY1Rlqa72zoTJw
mbz+GQPHVzeXAULQ4YwSuBYeIJHiM+06VETB+x/283NtTJpAW92drDbCwWoFyDR2tmO2X1OndRke
V2edSQeLaSPOc9BlDCCwU/8I/fBj0b/19J4fUTJxp4SYoCdbiVcz8jlpvQhqiOQ1pxfUUxK8QJex
ZtjJlJQiFbKn8TYkihemDzUsMF9j/F1bQoPl0kNgzu5YyGHaI/8YcAvWrjWU9+iZ6HGoiTZb08px
VmzXbZhr+RkiCSvyjiuRyLUDOBp+Z5FCw+/bSKGJHeN1f5sg6fOOekPRZtOUaA4Q1j+NcB1YgwP/
ELyPxAiRJlSV+4dUXLmwvGnj0ls0TLWBKrQAzmoxIR4vqTjzzyrWvKOh/A+iDT5261aHKuBFPI/E
mj9TcsyZ/WSq9FEHuuxBJQaR1DMcXn8aMVXpDRiJyFaxINYN2wGbXCyv85jE2EyMTsvXxPzrZLSG
yf3U1Ju6zTfJNvIgwqQcNLpt5dTQ0pm4ckC+0rsrI0H6XO/9N1RY+ivEgjwH2jBgcyGnrR/Ms3zk
uFfzBRFaFLYnJEtFGGXsd7riMdYAG7wWkAYCjVltjfW22ZAe+JuSfZuW9Y8WDtIAFGiruQQXdPn4
XYVEEXtvU4JAhxHOlL6Q0a3LfEOfty65FdGYEF/VDYBKMYQWSaFTF5U55BVJ6JbdEi9w06mJXrKG
tjLrEVlCwyW/kN/ZSwVOtm5wszeaWHRRmEQUvj8K/aO4I0k55ouq4YOXT3P41wzZGqMSSQkhlKo1
sU4qazOgLuaE5tuv1FVDZ9w/sm98TPKfaFqsGpPwOgX0zotCUTKZAi3ds94JD0HI4CBVPdzXMX8q
scv6pAD7SSUoqyNtTmkfJgUAwwvECi466E5MnxGiG+TMXWOFaaOy9gGfRHFISHskQ/LO9JV7Gv3N
cxOWhONHGgq6NHkKhH0yxEGGxZiB8gmAKOOoELIlQAilMoXJDGgBNi6wakUjk19iilLwbvaLki7t
xNr7HRXfJrGalN1PW+zhhtWv4Sn+WzGHa3BNntiG8s7oT/Zo/EIVC6VqJ8KVh0+JDKqnnmECkT3I
evi6aN9mCd0pLpuNHn0WK/HqXr5irPboDWDKx6wvWD2bjQ24PvbSeE9fNGr8iGueiMei7CbluuKN
ycUqjgGaesmZsB+7/CnyKKW3BqtwIIUfgjYM9WwVhvhGQ9NzTvwAMcHdNKnQOMd3Jdh4ezPkQe0i
BmfXxfq5Yw1Bt7qxWolcBtWwRUtAbhrTo1J571M4Fu5r1NcKsdGLWgjvIfiyK9t8j6qq+WAesHUS
xMQRa6S0zEz3KbP7VNgA2B7VRFnyZEBg938GDtAz21ssDZwgasxHRdMrdzuHi5gYkZKmbJ74c+mn
+8YVogpmBUKZG3zj98C0ml7KEhDs7qM9xNjVrcu/ssxzmy2276UZRAHcX11BuDwIxoIvR3iMaB96
AbfkZSxpaniHFn4i8LIov0oSxZ8lTjW7+MnrYGwcE3DG44QssI1dJiCUJdl/PBmbOmSYrQyNnt+l
oXlUjGsKUQQKzJV+30pIZSBWtDEeE5CQFPKIs3beUjaj3xEz3KQmprR1I+Y8Zy5sN0NbG/4YOB9n
/3Nl+uXtD4JpaUwgAHOrALaTqeS9BHBtohSTs5zvd2O2RcEOwwIK63e2r0tQKIKs7/OoSlZpb585
FOhOzBbeQ2RsoKcgwyUocodUHCBzYFG91iX2Cx4QsvLKkknZW6DiKGmrHYZZt5pP5LPWr6HCb5Ki
3/+UTAW4kN6BAkrjPfyb5Ey3P/JyOE1SKPiOLhOwPzaxUq7dR7pPUqnSS6OTk+PT7RV1IgPQkcsG
Pfhx1BYQ0NfRsppFzBVUVq1Ad8HvyiJmhyPpO5qOp1+Imsxju9A381KiMvRp3MTl5kiFZOwoTsHu
hkiEO7ZHkT9t0sTNJ8MEcHIfWR+LHEIkuxuCKXfGgEw/gPvrhoXopRNiNhBuKugjS5WPAVdVTLem
Fe38kwLQcQx8s0bkHyTXdk6JRwkAeDaey/sCdWvsfvmK0z4EzxKgF+Gr2GFrZT6E4tKqK7nk7KPu
PbK8ac/bhZBJc0siiKA1gvBew+/6RmprOtmS2KZjD2NTXb87DybVsSH7fFeQpGBparnByr1YEAIA
Mk3DF/+NckKfa6g1FdUWSUlfJKO4BcLvhUF9yTT4mYna0lOPCoNsIa4WChYmECol2FqJPuA2L692
x9zQns4F/d3qPn3FsIK6IismMsk+94du5jEf+nyrGP/w2kYZksHhzM8KXCGqWimX/IlYgkg7Je1i
5TTbe7udAjOGYX9Ar/qqEXRdv84hqMtwJHAkp3R60BIO6R+7mdfrVv2UPTvJCzgTQvWiug+/SwkA
0Z7mcVqMAsLMnxaJIc3tD/SmFu1uj7SLujdqfhv21BVe4AOR87Eu658LBZPSn+XtLKStHnyZoMwi
3GHVLalmHmMmDxFBA6D2U/TCIW/kp7N20NrtMjipcb3IjOJFmkrQwczCApdYRNnX2Jkt75Alzn5+
fcW6OdousXIDci/i89hCjQl6jERsTVB4lyBq7vNV2Rd0YG98zgQfMBf+HpYJb5Y9U/ATnMwDpAo4
FDnjF+GquGjRuFH2C5mh5xMZeS4LIbEss02FUGBY5mW7BZO1Kaiho7Mim8FOQ1+E/lM6fWfAunj3
S3W0Ob1kSxM2gQGm/T9Hn3pEfVUCZbecWfmS2FJUslRokGWAU/1iAvn7P1u4sALxnFVU+rPFlUzq
Liy+k+WyBQzJTSGeuf2YwED2IWJomxjSvLglzTmqaBEveUBrskxOUKfe2ZiO9qRDNlildEPdohmv
4OdesKPT84sMuSGCnaAw6JX9h1F3qUMntEhbkadfF1ogb4h/1lvqEavusBQNpWTuPaKTVB6yn9DV
cjVUICLNq4vPX87X/9HLd3hj+kOKV8jvFmnIPmr14Kc2FQtObfmOgIc2p3IdRpNcBKqaapL26bhE
EyIOBO7ZL57gjMXt7ixkNPjW235bVDhsi9iRn9x7EKfWKRiEW+FplLD3thRfE5JhUh4UnHCqw44Z
HA/IWGKF1xjLZn8bEtPCyC5jyMHfdOGb9rKxI0GTYChk33o/3b4EiH6xxd8nQGrkjCEyw9XKBpJ/
h6u1FgeOIpkgH3Axqd0RGgQ6/XwXpWK4jTtf63COu6BuvArZxrrmoh8PDh1cNRsXBFArhOwliSSn
IYLNC7DNMBd2UavjJBPiYwDs+pByWsm5Me09WRPnalW0u/Kb9A48NDSA4SZfNS3SRLKNrNGG2LHI
yYt3baJHnNaJX2EENotk1pnUlqYkJC7zmcj2goP4GuOb0dyxm5E7tpeSfaA0lz58EG1VFrxHFXYM
AQE8U6etjyQYA1XsxyqWsFnIBIBhAyxTEHFl/sSKvZSPczRI6YCUpzH/9fu7bvBxU7MMfixYpWiG
8pjw7gdMf9i3ny0ZlqZjUBaxnQRmIov1xbe5OQPz1w5NKrvZY4xAYkbGvApRGYjmKV04an7p1vId
YNxnXmqExXu0jfXGW2xU0e8MybKghZaK9xWla1lPPRCbu6Hqb/B4GTrKOpfa8VgNlJ2qxGTlSfdT
cxZ2Zd01Fbt5nF7CRF0IT5VvY+fl66+/35R0tprH9xf7fxgFFr//CLc741L+EXAMXdCMr0C6e8OO
Jl03SnzvINcXkLra56PfwDwLrw9QqgoXnCp+viklxhvE4pzvB4o+8pT1vbmWofy1YQB8X+O+/+CZ
PuznVfMC38mU0BVHWn0grpgnc4Wkgk6ThFXwrOqKbH4lxDP4nv6CgzwRLplHWMGnnXQzWnWmYOYL
r2AIkdZNg7Z4ds3lU7NlU2RP+GJhT3C0A2b52BadsD91oPKdd6TqWdVo7cMtCRkOCIKNW2NTPpYR
8HA4LY6V9qIIkEKDO/yrvQH64SDrDHDcZ9FDon/GkmsxQVgdr0jmsZ62cCD3W4dtbiF1QeW+bXM4
Bw0jlZqEyX6MGwnNZXCsRnTQ6uAZ8Jc31QC1E5j7vj7tg8WYGrPV2SMN24UJ+y5aciRYTbPktcO2
EFHbDKLuVqojVAmH7vCakCmrbQXjmiO4Artyd3KAqTwEsd0cYPN2PFMGkPFIE05qBDgRXdeC/dE9
kNXjzf3seyDd5dD0ofWMKnNpuGCO5u2QRfQVN8fP9lHRmncy7jCNJAiqgmdsJbyA9Jm1/zwAlmzb
TpynwakoosHYDhJ0T7lxP7z56ppP3XnGZpMCVzRNo5Q/gaFZCmKDfNIZ46b07/npf+w/B4S0hn2D
2hCSW2rvwaZAj380om0kMt4+e3N3jx5vlXkq8xhRylRR4jcUx12DmaFhF4J2Hp5v+h4pbR6Ch9nQ
W+dyxerW95p6H6ButCOTEBJ/n1F/M/KY6ErSni4KxD4t9BBuPfcWRXmoQniJQH5IQ6R9AqHD6lAB
zpid2G9lgfXt70GYImEMKW/MxHjMElW1qVbLNyuO7LSUDzdRZTUx2SM7MdFekS9+odmZ7oY/JPI7
rrSLbxzIQcRZQtBAehCdTZflfZ3dgSvzSSIOuAHcfrHc+3QGtLV5SQ/Q0goXYDGXb1J35cRuBWHt
XVRgU2/aZH2pLwvSt6orDsF7H2jICpfk3uNXPYMPPotI3eew+YQVC8T7Gbuiry18ActuWvny0+ib
FOl8baKsozCc19rwrZIBVQhahatMvvyi/bDhFM7QCl9i7t0g2dF3f2WPOIHrvei64OlrY7yCJsne
ZMBAHxKcg7WmEHxac5qOWf1tqfmwHEfhTOYKMjft1nK3YeQWx9K9ejIcgLv8jQQtK8Ecojokp1Xd
U4F1PfDWeTsjrEjkAONN1oBG0Lp8Lg76WT8nIHuz4bcrCG5w+kHFjrw5RqcPv+sYKTcIccTgqXb6
5SpE6jLaHVm/ll51+xIkclbPkU+A+tp0fCHZg4ow1/YfJioPFKLQnTN2+zF+EzPRUrpJIYx6nKug
xOdtwORj+9/jh9grIpzOkkBED0AtQY9oOvbk8FCiugpVukeZ55ayfDQnbQNewJxaob/ORLGqEO56
9soK+X4N/VoubmOx3mkXQ+emlz11fqbHLuxJvZcoZrc8YHAB/tRr8oB3eTPadulvYBE4yHSRQLmX
huw8YhI1W2Caqy+zyUcu1t5jGtp3JkecV1hIGJxiUOtT9Bwol5Lkj9COmOvJlh2HfEL2gxjovB5V
1SKPkFUHN8iCReMLv45kMilV+ExlIg93QDmQ/5J+bNHIjowBa2d42C1+knTn6vB8UWqM2kJHV7XP
s59mXoEAr6+S1AVfLl3TmO/fLEl1nnFmGU+wv3QFVv7hWKyRO1dfa8Gvg+0MBlF3pOwTPIBzY89g
TMBAFMtB6cSk1SxDF6IEuZETAHkYK83RJ1JhiTElrO+/hJp0CpzDpn2xlamNMAKJU2rJxd4Q2zBR
gu4u5DhSZw0eLf5emPzzy1P/yUZdCj98zlxAyzhQ7SDuuwny4XB/iIZqYHhSL0NaIrgqWQCvw6RN
3alhWnEx/ZF6vAWH11JYCemC8fUwddbVZemwLr3PiUmyhvtl7uB8O3i52tjylgjvx6tiHkpSNXSs
X9EiILKbv5JJYFBHWGBrK1QSL0nVKnmSL6BHpcn9QpDBSuwrjSozbx0Fq787ubHS/K2Faqy/s/2r
5UTT/KrpIpQqkbshyKUPofxYFGQUj46FlRZalPwuBGCydHmEQSH+DCntukhjAOBiNpy4MwVdoR3T
jA5L05/n3y66F/ZdkJ2Md+B4gPspSFP6FC/WdxD+uulZZXB4BfnjVkW/gCo+/gtbEoXnLU7Uz4tz
2ZU0pA//j9tWD3Bvh874c43eh7bkoIwu/ruyhGYhT++RaksOnSOyTapre/kXVK/8XaPZVA8IBYm4
b4N7fsirnYFdc6fe4BQlpXdxwyiQcc/3BbYG2KYkeZUAGAxj4Ayw4353MPAEEaKGmO9EKBZ52q3f
BEx/cN6Vhs7s2B+Ls2sGIt0JlRiZ/4QbWTvaAIhdF6uQXHC58lKD7CbSPdcWsBQHzSqzDA7LTOTi
FzWGqe9zzxWeC5X2egc5sDO0xmPUMISO6AYGtbxDJ6CEIfx2Hkc/41BdIFA1jo40wlz6l3ETV5n8
M+ehjwisojnC9AExRhZosihGBhfx0Am+6ACW+E72NOaAXQ7QpWhWgUXmi91yRoqnr9J4sxtsmhXL
whHO+qzXUac2rbfgYHnOldBK53v2cDp8DAC4pnY3LxzHZYQkkl/XMqfHTTb4ZgEJL1D/EC6wgRmI
kF5L7XjPelKFFoYWTtSmSn2UKJgxk7QBRS/Z52ivICEs4SUnqbzXI+pGgB+p+T0KOPTsm+mtsBpg
J22mwa+tiJAzuR85trX6Tdg9erYbq1QyR3pY6ZcO2MMa8zFV9/F6JjbQEliWAYloOrblNtlrpkvI
fWB991FL2vmHq0R1c2oYcIH9K7xfypse5wlccs4qxTBPCpdys4RgaK5Zh/drpEYTCB2pgFsy9ewB
knU9hPnEEed5LedWZuV3UrKo4dcyolW7FXTQ/7pNEh4kp6rzxZTszGbbNfMzWMSkI7l2ZnDQg3Dm
CeJjkJdPdBGUBdSPAvLy8WZpsRZteB4IuHnIjk0mqPHS6aYtYIEc1ETW9LYebHh7mKjMU+DNj45y
lheD5HIOs1yyvQR6OaiZLH/MOJM/Ej5kOR1iu2LsXfv1XbmcNG99pogz2WTegg8fcJrSqd18E6cB
ALkJyOltcCGoqlDJxLznKhQugzPnjvvleT217XDp8irZG94Yt+Plk7i0c/ACRSiJqD3cRH6rrChi
ru+pDP7wWksrmj4WLz+IhEA+9lKrnS5BxiupD/WKyvnVzFusgSrjGP0R6R0pSotHWFbMMogJe0zF
LTL7kSrjXJzf2sV8EzQOeOt2WPeKjxunHDg+YpM4DvDsSy1BrdCJ/86p40E2hfH/lgeSFCjq66LE
tYQE5eBAS/YkgdH3d5H5nv8pA2dQMM+CkZ8x45YyfD4F9F17qnnjpD27c+kZDi9iZFDigXz3MHYF
Mu/6PnMIW9CcbVgXMAvPXxFacc8u6tjfXppqkNougWAAHG06bCRU7bAcmKJQZUzUULoWz1UXluWj
RWNW91PiDe7fs9ILrpdVTtbroBAe/VTZliLoTEIuQc2AjR6pzdxhcJDP5Szf72J+69Dzy5lsw5Lp
Yp3AJ/sFmsRcxoNJ9kXsyR7Ms4F9rT4kHcvyvYh6lp57vM5z+uggto8MIqrINcnHsVPSdtK/TKzS
dI2XR7OwhOKnWAQnWjoG2I+kkI1CHU2T5w4jsOR7jqI5Tyb0GYcUiJP7YtALEIldo5FzalEBLYeH
FC8KKn+AYWHL7q5EeA67mZvZEGEI8ErDEIkI4QG5j5LgAtYediBHEVXKgA0ZuHWqgMjUpaFLoFAT
i9GkYNK8QPEnXI7YKDb/A/c9oSLEWms0PxfP6b2+ZdDfWlC1FtaOHtGg50b7WW7WSyOZz+VHeloR
zn9ekM/4PV7TTlPkOLByxeW+yDQwUeYgk4wSC8omzUALAcrX8WJHpFKzlIPhFx5hNPK8HcTdmvPN
XQgsznRcdvZZss+k+Dh5XM3HDCbL1lf9tLb7j9V1mDv5DXBS+9QgkXmutwmwZX0r7C5IeIXKnfDW
eq3Dwg8OWPp37CUYksE1Svzg0D8ES/hAWd4r4z2rQwP6BZnrjW7f+HdHGa4iIkd8Ibdv8OW389z6
+zH9hVJ+s4HoOjqVK6OcgA4fF5PTxZ5FedkfbV3qoZ19lAbKrGoP167C05RwCUCHLfWTPXJTWTtN
2t2CX3pmpI3qOqTFpDLs5RC1exYt6gDhHA8aGVeVU4Z5b8bAJM2Xlihl2U9geFl53gXcDlrsm8aJ
fcj6sn5CSHBHNH0yiqqy/T0GM4OYJiTkuTN/ImUwU7aKvJj4Ffg5VbfHb2y82P6D9djQbShYsk+8
qMDzfcEFbTlokmffQpKzxPUXzRdlK9BO5L833q50R1QT1DYQHLYbnoZoelYSb3IOJysLLEHtHaY7
XXgYFkY//4KIHh/gQpYS+Ix44Ia4svCDT/CpRoaEhQdkLFey2shGk/WJTQ+GhomGPieQD8QJadcM
MukxS6xm58TrJiydtc14il2LT1qsbR88mcEaBgFHLSTaacj8szLwV7PFILpwq9anNWw9EzB/UTVl
AYCLY981bnspK+abVf3JcXL6D2IxeEXYOTyYKn+gkxBYBCVTS8lskjQZAzo9NpHD/NROUt1q4lci
98DA036bmvEw0ZgyFOtduAn3BTwvjbcRiWxEx86h9vkK6mdPCpGUz3nLk02PBXIp3D/z2WmAWSKF
sXxtF6JHSE7hxmYVbV+VM5anPvYs6h5tTt+xznL7fuMnAklg2z8L8V+/gdGf60rGLV7QN82vF5A3
13Mr+GF18OI3zDLFlfWs5ZdoeEEq7GF7yZ794Rz+nAk3XRwyG7o4IOx+40NkE/m/yiKUb8yLNAjy
BrEThyQgwcAxYCapTETVK6IFqo3sf8dCyHJP9KA9n122HnFk+wE3fuZAtu0JPHXvvYSLARi5ss4z
POzXu5qUX7kkH3o5LEsIfsZaC96TInjzzrTFglpdw+M2xQhyYlh0k1UMO0i62x1HxI+rHWP8aSEA
4lbRS4bxHbF7xnfNkxhD8ntkfGFS13JK0Ijl4hG5hreWSMI1RJlWNjm16ktefcO7/gDWe3m/I7KE
O+VdI4BlIdRFSbeEGeultkQJL5MxzR4KPzZVGkX2AmxmdTqkUa+912vJMQM+7t6cfiT4QJCG6hnK
XDjni4mMWCapalEHTCi8qMwl2n2wdznkZoCAwh+OcX0JNfEfbPTqsLLsC69mu9Kly8NoYs7Tfs54
5VIL4cyDBeOBbV9qOGhoiL9sh1esblHtNR4kEyyo0RJ/2jDZ0b+KUbQw+pAR4JRE3zTlemV78/0n
lZw4eHcwwSIhLmK4mW1fFLYdYss7Nv6WhZ8Ny3RjsKCyRcSDnSU3DbdcB9jfzRpozuOxzrUJNPa+
XdBTjZPYtVIvRXmmKlqDz93j9nEcU4VQUo7YoNqCcOBcoYO2UTzJT622f7wEmiAV3O4tjfwWr+G5
qDA58sBfAd6gDrd4++i2bQZmqKN290QiUULp3zTn67fg9JpLNpDkijLX2Ea5EG9hl6wCiVHFQRYG
mGsV9fG+njYfgYnEo+XLDYZMjAuzBWfEEGqMPi7zAq32MGgKTqSeLhBJsz2h+upOuxmNDOa0En9g
5OkKiJnuDAAqtBxIj5XeB+ms70RTJ5I2DZF/0ZVdZWqrMiExzcWC5dGw/70VpdWb45v4G9k2GpwP
hNaed+b4OgYjM4q6xXxCq+VcKUvr4+QVqI8wN6tv5FknxHBjIs8vbbdwnfqlcO89kuld6sfKu0lm
j8hCwOTNTEAUNc3E+chz2xrPJtv/adfwFRFSdKRQVyIKdjduLBbdEI06lsMgpu7d6Lju4FGp8MR8
aZKZpR39eGPPYtQN5a2DAasDPyGyohqCCsdsl8HJn+V7aC/1x4vsRt8bLBYQHVl7rkVu74x+S4au
8pAA32aOVBqmrrGdeBH7Pgn5jKSNuequUDz6Pzlf6cN0pkGndT9XIlUrClvZ5p0iMfNFtluzftTb
qZxo/umNYl6x+vPanScoKnMD4sFEdde9WdcWt2jWjxh4t+5dnOMq9CqLWG5T9KvVb9UDjmy3n3ey
jvnHigFbDjrsaUtgzJs94cUT1XlDeBpcIaeJYYYt8jTlrrTY5WdO4oQViuTBIJBN31rE4hrZkAtu
tKWXYDs0I8LugrKsbUkTY3sbLmtlLYHUMvauc8tZFH7blljsVhUf9e0vfzJDaNK8y780vy0zseRg
LLt4c2xPUQYU84xqxyUubA/5a2rgtl2dUQBzifCFXZjZLLe63RM3iWYSdlSl9rvmWJBGMDpqtlZW
v6+H/fNLzvVV1dF5RXg6X2xw53gaxWXLoO0AOXmI+jtiiBUoILWMZX3N0ABcx8eD6avF82xiTWY+
EfZAhJhyxiNCxYizaqj2j2ORjp5+DdYWek/ArEjLoxtAWgtF2RqIoFtqJDZyovmYIX0yGAmeTTBx
RcLoWxHHxqMRnTYG/yXkQ9tdChGHBxCIXfKga+Wv2gbgAokIH/NcOEZ7u/AuaN0CwHuDLfPnEECG
KGc1Vd7Y60nIugLyc+AzxB4uzsjaNEzUD28bKojn8MLyzZdEUlDJC5IAJvEOFnJzxvqO6SWeoZgc
faLHYa4zBKvrs4oIF9j+O3hcmKFk/VbXosRt1t2fOxQQFGyGqTFCDporAaQ0kd3fgJpU7sJRqRwn
lb8/ewGH8VoyiBDtjLx9M4otfXLnAt0z/QuwbsngcmQT6M7k4eiJYww73kjpANRh7NULN1TVqZ1u
LC9aHHrzeYJRcfboVkkmlPdYc8EuqYdq+zd2/a2jbzgoM+luw03rfuUEklCVTh4i9CJTYlHQAfJi
9jK0ok8DPdtUZHGzxl3m636wODNabZQoT3y7qOyBVe9W3yXxw+oqhAgWHorN2JXUFQvZzhksesj8
mMNGicq14NfyWsmsf6nKZEY8WPCFPzB9Bi6GielkxZjA1IU0DqzAgA7xN6TqWb2F9ShppJygTX+D
IGpc3r72BxKyxNjZSZzvsW6KJ90a4Pe4sQ6i5IaWz5YdTaqBFAbpmvjasfilt6/Ljf/pCcO1McvD
PzIBLBZ5nZHdABarNci2XcebfEXnOABu2oZ5IrMnc6z8YqRQnB/IbEnMZ/Jl+Q6YVJOePPNhivtz
SLtfA/OS+yHBj6SLK4/98cq/W/v0mRFciPA16oe6VOGEANbHDtWKpXSglxqFzcIPxjjF5FGQKIpS
ilZM57nmPaGqZX8w2NErgnAJRpvZy7yTVmEAMbZT/aZQ2AmBg6e9ArOqPZ+stB3AocLJ+GrKyiBy
eAUKkAxXmqHjaG7qqdbOaLGAwgQc8VQvttDpFObULew3ZLYt+1lBqrBEhJjtKmdegT1sypa9cJt1
DzXfn2ghh7ZIl/FHK5+TALA5c5sR5FoBEV76praK8Dx6HJILDbdu3D6oJ0VGJb6wph0DEFOq+m+u
vjLrQqPqepGuHYYA40d6VWHbPajuCJv1CkdemaIxjZfYFZhLdEFm40ss6hKR3rbAaR8yc5SfhvkC
va+QI6lcwCiBLvHxQHE2Chg2x47ZwD68nWsdwaSnHLv2QEjDah5zGp7jNkSEwaODqSLnStbPMtit
M2jk9cMsPnBhlvd8MyiJb8vuRL/0TQmSWSzFh+brOSrPQf5XteGaDGtOsANka3UaYemUncrrA0o6
vY/GkcHwD/SSZhzoue2K+Z66P2EESwV+YmmIf9+1M8sYHeSMQjyt+oTQZUbt3XAJ/2BUyswayGsZ
BeZ1WouIHQuCSpkqBzyxOJ4lJgmjC2K246RyOwmKUnV7a29khIsDCGt6haGewutBNNioCd0l+roT
xRvRr2IDpTJHpvhVzHTc8KO248uOfnXqkccR2pb7D7iv+F77RZDbYCruoXjOK2pwK6/pr/IU7qm0
Ix9KqZO39J6DolaA+sJ/D68oBdE6/LDCuPGmRMJeVZqUBoO2DHfJJ6eMJOUXTUplDLLt4L55Zb5j
/V/QxRLhua/0GtuMs0/wL6+yZFnfFNlvx70H1WQUjk2SXPWcmgabGe5kwIO0lG6yiILmIUDl6a7P
xkTzhXqKBaxLwe9/nxrwmqix9j2/Nml58JWM4gYNUR2aZkrxhAg9PvZ0+mvBF1gQeHhOxCxuHMH/
y6tRmOWo1ejJiBIqQa7rmZjgxM1UPO7vUYFWPkl9MoRd6R0kTQyhVtAW6iobrykAGF/zcUGYjmfp
XY3fA1LiS/Q8lnwduEtoSGZgl3pW82VSItfJWHV2T93XRmdNYlqrFDHSrb+302g13AbnCiTjn7G/
jynCQPoarGAT95+qECtrXf+r68IXiTF9YTelsePTUMi0ZTSZ1pe6QU1EEwh9rs3qHzkAGF6eywyY
iwvioraWUq2LZlhDnJkLRpPTZSdrN8glLDqSgfNhbT0CS8HQJpL5bDaRcKywheTBZ5axcqO3L6bS
zTgSb2EJAC34y4GZ8os96YpFm5oYQccdANwV20uKwtAMQaXL5tXWFlgpvMmgNIeYZXTjjAixe8dZ
FwdXj3PnDeOY9gHwLa90aRJbI9CXPYZo2D/pjRDiUU8EzPcz6sTXMqMv20kFfsWYJfs6BAe9YCWa
6KT4i4K9PTrmzfZmn2Byg98Vj9Io7upKrHqx9bnPz2NLEni2zQwYH1wVfD9WGxYKY9N4Fw+UoKk6
DiV8YcbrKieOriT31g7k2RilAOsdsywnWXnkBovGNBKUfYx+ObMR4B8ObawMD+MrJusCb15DqD7i
wo1TDSlMVhqVZjwmg488ZGULxNjzt3uxRrThDZSSnS6vwytQrFbkcH8R6abfuTKT8Dd/0pm5r1AN
bBAn5WmKwXziFbpcH/XEtERbVr4yIs+8rCuwRuxXL5b+76juL7gG0gduWDTzvVEAgMYYUf/eUsbL
LrbQKhAirAavamGYJVu2NzuDwFVKfbdwx9a4IhAzqsugKo0qPb0zmmoxWzpQgd2xNaiNZkKRBtv6
2K/HIPqph8KCE3FGS2AS9mfgQuHh+0sq00GV4JnEQQAKWBmJN40EY+w0eTxupu9z4POlitBKZtWt
IMK8lbIVKGXYi3fKjub+yY4eXnu2TicaGT6n/JPMdF7y0Nn2XOy9e5x+P71qbjuUcfDFuJCN6+4w
biBgnTgQqWeFWiZpZDPnl1kjB8edbSrqBDbzOWQbJZQicXT4sNqM9zGaTmBKqvoG3m3F02hdwPo8
hUZb/N/Wv9oxM5p7xQUSduS51Z0CrFXIWiwXuWSaFDJADoSb7/NYn+ioOsXgY4OxZDcvgpmrghTa
/gt2ki07Bo1CXa7tyK8wCbwVagn4leyNZzIigrIjIgPn2AQPgywVFZyC5Cc+szVc1XuwEnKh/9WU
o6hxRdeGDQ3klJZdkdBP0jDnv3m4XUP5BmM7ue3PYbYYMMwv+PccszxeQVBedYTPqvhyOvCkkLc+
t+1wZvf1YEQKvr9MhRkengghFMyQkdoPxz43sia5N6oven2jp7ovZaJmDxfte4ivm2v5CKvsMiel
TYiWn9kuI7ovmoWMgFZ9nKjHcZje//Ch0T5md931h2XfDK+S0p/A6LvhkgqzBR6zES+8qoYqdkSf
Wx3dFHrwaEUyfdy1vgF2cWpcvUg0hMk0oqwVWnJfJTAwzg347HZZo9Iru8gxeoRb4qjl0d5ZQVVb
bxYZ9w12zIBX8EZY/Q64s1BWrvEJ4hblmpDKcAPugtKIcuXQqrPHcFPjWIeYudgtOb0EZeZ/Q0ZL
vX+gFmku+B2LWgT7zktTf+Mws9VSjvQgfWEuk9wRjcM5K53dc4MaENjIqoHEIVjHZqlkf/C0qUiO
H2y0A2XOvOTHzhi0GtoSa/JMQBkvMxrRPBZ0960QWz5KrXhXJ7hCpLMRip9nTsZq71iTIA077IkF
IJ0pWoDK1cBA0PnePswPE49ScHs2SOzkEvc3LVVW/dvNgwgb3ZDSfvIsCXi7gTAO45IWtQjdiF8M
4zlACTtSDy1nkHNX3Osyz4kxvk9vFLeoj99fLnAN+tdGyFleTuIgDWthWOoJE3nW0RGn94O14Xpo
NvSYgUxWove+6aYwYfILxgkNf9bwtV6oVHGR60ukddGV0r7wtJ+kCp/B2LuSI3oRPwsjbWirW7g/
KxBvH3GGaA1F8bZUVITzql38Pd0iBUwWvMHk0rmSpY7yFKlrcma4lWeRnwmsjbnx3sKHp4A/7Ma1
i9odMqXum2Rh9b/F6cJIJJjWA57Q/rj4bQrYIHzlXKHh6VIOQ9ZNcNZFFGBbBANbrKXjKs9MBVr3
WemsRzElfcSbI8Mzl/+UN1RtDpKV0/Uajx3UjrBbZTDRLCMB5PSFPslbfbpDYUQXMh/S5g2oGxaf
desuPFu+LD5HQrXrsR2hVLOo9WRQw58sW4qVZtdRAkpNQLnM/R+vH2Z0BRwmYyxsvE9FlDxX7PhD
n0rgAKIfXUg4PyJjbk//pAhuG4v1Xcwk2l/hbEPEeOrJbCYsyC/nTr2VXe29M4VF3faOPRdnG0SB
z5s7xe88kGkesKEVKqb3eZisNTUcbL5XCSMHKLC5U2neR0RNkTJjd8ses2taZdoEQinc8N+2bE40
nwYPdaTmbxjTGXSUgxqV8rWvEOcuebEWoBZdNPbvePz40f4crPRVhRIlejqbe8MW+m8A59bnqilu
bfp2zVy1BG4cmKHc/pxTNqvlddHckfyJHrRG9EGubPgjuDiBY7o0mkhJ2rCqv6zkTqUWHliRJ2/N
D7PT5PXsj0fmGfuX/2twvs2Z9Dc3hUzs7RL7aZ3yT9M0oFhiQ0NhDpXoxzmps6KOLBq/Uh7KPQeN
WaXYkPhm0D+QYCQRLrpCtFrK4jj2Ytjgpyc2v6VClOEHLdMHf0vR43/wJjxBTqE9nBIhh3h8sIV3
ZF1NzZZWARcPRqlw/lDbBiyOhD9WkfmL8MLdIFb+NHB3+lCQBCBx92PShY4UT4wL8SoRtk8mnJtv
ommvoM7t8NS/T544bx4PlThStEbSoPCoOVI9w+0+Weoel0V+UBzpsfVoC6fa/6APIfbTzFGI+E24
o+0mk9jdvwZrPchqE8pZ1ei+DB34zTWS4W2OFIvmY+Y4Zd69wQ0V1Q44DniNJ8BjGVdMlRVPdBsr
P+iIuSnE7nePx2uxDxhSY0pu/djW1KEt7gM6/EyQruvuNjgVLk571ITnJGaroj+sHKvGSzObPhRh
NHPV52FOAK/PdtjvLbKuqdKZ6/j8BIi9hVvKkNQJTGVJh/7d0WYQio7kTMiYRKLm8v8rouHqqxk7
8TVYc+xZ+zSj2caaC5dF6Q4jbOorH84oayfjTOFasTCpxBLBTSwcsRoa7+nKiNHVZ10743ZriNXL
yjaSiDl1/xGzNzgNYg4m9CspAovBxBEjDD201+bkm5tz5+QXWlYCIy7pqTR50qKBJK4wnNG8nXnC
yX3x7V75tOZIPwA+gO7Jco0WHMSSuPTkZObgj5VwgG3/iscaUAb/6qpSI5tNK2TsleGp+YrvFse5
s6q7ZRrOcAeRdxJe2xq6y9guMMas442Y6kDYcbZUuqW8XypXCPLc5iflJQsPu0no98cH2edYbZtq
Bwwy3m3wAt/x3YPnQyPe5FSslSQYD3m+PSm1ObwEqAahX9/BS5X+EQXhblHwaDoADLGZ/LUXj868
qZhS9psxn3HiNsaf82VaHM6JmWhf8X1J4EVJr1wlm5Tg0Ds4eQ59BCNSOfavFvfnev1DKPfGB2PK
fqFL5jIeBlJGDL3TbZQ9FI9vZnqf56PY83+nLRwW+r9v9MS3TvH+xrNTay7pdUJ/iO5D6MYuXi+s
67AfQTGwzTW9G9TM7HvNaS62IaxwhLKCID4NAvm+xnx4ZZBVVwo0g4U0SK+YrEb4Fg1NHAhVcpq/
TaH2iX0hZ0E/LRNlvipXABrd0Pom6Wx98IYu8IW/WAFlhBBge9b+D5yPCH+rti4M42oZK6dR2zkF
nDV/NMKWDwKqmK15ezH/000ivRuyg9pnfZ1F7n8BFJROMY59KoEg/DlJ6XYpR7RKt1ebVg7PQ5Hk
Gk7TWV96/nob4RmV5WFcaNUdceEt6H8KQMgs0oWIyxEzdyMIjmo9PwVFsdkDjUS/nm6N6udpP5Ez
XDiQo3OA4Nef2pyqvXjQxuxAZcjZyGAvywwzfh8UtZsNnScqlbaeaYkiXQf2rbh7Fqvelr/PnTS7
Q3KuOFbbOiyJwNYRQkYm31OCdLPeH4a6Bhm6mi+NWezDM5LcgFKUnUcqP32ASYZo5VmG64pwgUnZ
pi/0F7NUn1lovWZjS2RNhec9zH6NkNfnCCD8djf2c5vnqe9Xw53oIJOhAuq8q0gxf+kYHV0erWg0
Pcwz7dkL8Jli2+wW/V1vfNGJnI8xOiCCS2y55SUaVhIzw1BSR6cmxbeoOrvyP59q6RPS8T/0CfCD
V4zpZFn5M8mIFD6oCiptoXUDwyXkBs4t5tJPAc7KVC3+QXHN6KmeTPMb0YtXa0HGwACdGFyadkCQ
8YpMWyQuZWVuXo5wZoR1YlQiXsDmrkR1vJoBgBXrDTXcz9QuCCbRk0q/R2vRiK2Vtw4oS1gi8o8m
U3572a08Uzunkxvmj8dHW+XXGV++DqcuEiogXNVShfzVgR6cm3y9fpOf5HCj5dy3ZbDzzQ49Rlxh
hdXYJyFx7YVfCZxudOGV6sfXMgYl6SCRPVBRjlKlSXTqbzUwRHtQ3jKfX7i6ntECxgFuf/Wf6pAm
xsW/iPqIA+8ACunGNU1QnZq6Jw3MrJXCW1j9rSxxPGtUHqCMzlM02qhkBXZutHd9gnoxlwnVa6FW
baT9cXjd/5eNltFBv8RE9k6ezOYNqqZld1qfCil0txnO8kI54LLx1vD/gyS5vkMEXdFuD6CveIaD
TW3G7lWoPsCftiFT3D2dUkL0YFIm2qR6jbXxnqS0mymo0f6qe21lo63jLzDtCQmBBDrSo4Kb/O3p
gqeyLrLDSlpFiHrttCiZbwHeoQXMyrSjOnk5WZ089b5s0pHmzEWD+cfULPDNENfED9aHw/7G+FZf
A5zkVl3PU7R0i9qlObaaQS29XLb/V/mpnT5Yn3Aii+3T+3YdJt9VS7CKwB6MSgbdNtXAllODvDsj
Aj9lVUjUXNyJyudDSqvBVwgzoluPrlCO1BZ5I3Iu+LbBAzVEeSgszdNZfhvLqGz08YXDJyYWy0gE
jk/ia/KjP4VV/QuB+AUu0ewWo/lvM/Ya9FmheA9N1RY8j9+QgB9vgDp7kIBB3OgQLczKU79i7sEx
zRzS43yNb5bAJjXKsXyooE6+3GMYjvXyU90OkrA21bRuzh8LIrzuP5XloFo4mv4Xzf1zFU0N+k9e
Rq5Y6B74OIFdFiOX2NRDsxgiTy88meu2vUk32j7J0m+WHRYH6MiK9es10rbkp4BlaC+3iW9lz6Pr
4uW7q2zhomKDyL/TVEgZZKwxcaTQDYU7QvaG/uCrR+wG+JBQJvY/C+K4v8XC/3e83YfoeVFW90VK
7wZ/C6v4M6T9qj+aKq6ZjufE/vj+Z6LdelWhq8bxzH8NfQGhFHZgaech56tiyEYzaQxAtVnJRCQ0
bEZo9IT9gI7LsXXKn0+tX1k26Wpw/oCHF7FNx84qanlLWHjpbtpZck5FnAGVnPJD1XURaWoVujHh
uhjfT5x5imn+C3Z/lKv4FChFaIZiYkLP1zEm3P/YzP40rBAY0eBd0Fw5it2NM/jEBKkwLJdEt7tu
oRpby8UXC44LNoeKuHNcKUxffyJ1MWZkSsMrwNazV3CzRsTd4yi8s/+Ctf8MopUIbqmTpv1a9u1h
CE3AtOVnhdOwR4ds75xoVx3QpSlE6z28azv1YktJ3qm4T48wSAVRiT4EOmUN5IZ+B+hNbSy+ein7
RbjSmBdTPnMZ7VxLyx2tMm9Hkghz3anrJtVGR5tndxSXkA3MiUB2e5gLfmi9XrQsmJvvAAAPOPXr
jpvaKyoT35gLylIRdD1Wmjbx4JBUEr8zaKIJuvgvIOaBz8/ALCCsrqqh3dnBnuYtgsT4JQPTDquV
Au/zHXHCP0zNn+awrUO2v9zLf1ek1i8uPvxS73X/j6cYmPB74lzdCdncNO1mxT7oXdsSbsQSHkiU
TlGNxtZGRGZfcz+a//WO+AP/v2pgRJIDvneOlgWfybaxJrTg2tSMFVu2ZqKNd3Xpn2gcY/k5qOfW
1PcbwcJK6PCqpwsQrdoCi6xZaF9xqIHL3mpoGmG1VpHtzB37Gf6guC9Njrbn7QoVXjnVr6Gv9P0M
jfhEfgRTpZJfZUsEx3ORbKNykgTKFWbkMQVFXYKeKQSkvMDdSfp5sHkUUAJVqWtNxQ6+3DopKJjs
pJZdmY5Ld7LOU5tVnNNd9JiLWCoPgPfrTtPyMoRThIu2DaTiIL9uh62YuSeGcpkkv8VYKW+fAztB
qtzQu83YUb+/BC0BL2VT+iyRc102pJOD9811P1DOfGY9HPGcra6djJpls96dJREijvaKmrowlq/Z
xeqNHbfKu9P2mtikyJDqumbRlUZ/IlpCvK7m7c2Tx/dbkdLv92CjXPNjtEg32gbmCrSxaoJY0gwH
s3vLK2+bXU84z+JKSzU93FAcxQpQLfqYjffNeGQ6PVszBRe5mAjitLpjZlCcysplArmMhYalH4ku
iz9XzEtSMcOw9R0Y04cVSEYhVE/N6fXlznUuz9eMR1J2zp9Vg1ajDQdL8NhLPn3C51M/JJHUQL0f
U5W49r6gYLR2UUkgWv3QwN9Zs/mZarDPYBmRli/HhQbKFxbz0ZzTMU1eyesZ3H0uqTOYGc8xPFXK
YrPlN0fk9XtqwTwlAOzVWUXvyGrUAhOqXNfDilz49zvfIvplxncLsSC+Sln0vJg0/Vb6JOKAUQGd
VoLAUpDhXbnRwz4RSDY7XTUdaExrB6NqSO8QhrMAeYFbUBnjL88jGe/NJYJIvRVy9yrsbTQLmmtW
YbUX3jDh7gjrCw5umLHnSDIggYoxg5cG+z5Z+7VAPPSVinN2zGF/th/dOr/XcwaEw5bDw8zyEQFS
rDWTjMgtJFmf9bt7OHgwqeF8LA57oDzu4lwjaNEhMpvJelGaIFLvx3QWCr2sDwqZsu5j/sKb9FRa
/yy1hfq6Kh6Den60obzcgGBwG1iUsb0f2HBPacrXd1jR78sSBfl0YsMboUp4o6es3ue8auKgkA3w
J+aiG1+BiBFnEwJY8arear5265EgOAK157X0EtjVzXVduq8KWz5Dm5Na4ENyXYiRRtjYwFMA0NFh
61KUNw1SexrLhp26MRlXQylNkI6WTs1gukjyL9f3ybv+6L9Te8ffdQxc3ajbeQPo5hEfCRPgGvZK
jXAAcL8qagLc9C0sx25qoUzOF/cUCh2kR4NjDtlyY+1TA06033ehNVJAVVzjbNGUDSt5MllyDpKx
3VvdzRI00jPHuABrwGngeEMzR5GUQRRTOa/kpJ5Vr4UFuoqq8g+rlZBgWKDUKKFsEisraRPBiBzI
Sbo5sQGFk81lXmsO1dRe/1KFgF0yq4ck0g+/hQpq6Ck8hcxH6VnYq4eNAxWTKVxAIN3IjQrPFBI5
ta5auS6cVe0tHrycyYGHyhNBSzwXX8NQ7c6WXhTgUgjq12Lo0s/Oljuny4xlSNCaWF+I45M8zibw
69LGfucoMNjCR4wBXWJrgzXOAlIT8Bc1twNIXEStflbGQhwE6ua6tPXraSV6E+qNEyE/vCj5x0kr
d3gRHr4EIwTMn0qqgD5lvMxTtwmSPTmGdbM/iHD2JO0Gcw92Sf3bZyY1w7wbxCESI49FbELSKG4z
lrOPHRU5FG8CfvO7uFwNe0t5Zm13gePh1FXNiefe68zKSHv7mz6wKCMjhL2K1FGZmi6+mMY/dTfh
7gzuPbZ9rU+9WpJU7zsmqSyjnvHmZGQVHqoHyVN2F4vP9rL9L7fPFjTO96WByH/XzSeSwh+H54OP
84KIuO6sprjJ5jd10UQo50u50hPSsuPFh5ydDt7tz8lZTxlGPrKfzmD8OkNQ0DoNKw6i7mD0mewx
3Ec8NvjeWnJnQVPGLesSMsqYqK6f9SCLEcg/tBkf7UUClrCD6GipJB9S/tdzLyJbzmkNCeCi4buW
vOXcHrAhBg0jk12LGqEK+PT/va0LzuZoO/vJHC7IYwTEh1O5FcxENKnkuSzFmDAOIOAQyOp+yqLC
s92CXx7OeOJx58Qx3yv1MtxknfEN8bQ2KJAFazUBRCWZUDfySdIsjbGFHkS33xkgLdUBdUrkiDtF
P3IsvTdvshtidaccAVRv4vVs06eEoW/9Qb4Ar9Ajm4gG3jAhq2e4I2izjrySX3U4XDa9ho9g+09q
eXcF0Tuve1Mn2gij0KgoFwAlt7ijZFEh05Xd4BhNKNw9AvWZX+98tLQfjMiZM6VJMovhbxba7m1O
I0S3qc2VbiH1Hv/+AhmK4CC24JC0w07T9JWs9yDXD7QFmxuzHysuBFzZIxdHDypRZtRHS7CTN+4t
Cgi9Kv4xWSNIx7PX1JWzosWUR4mJXIFA24vtRJe08OoMwchyC5dUz3BMWaPnXgeIyT7HRN3mdQLQ
C/Uv0xdxjKM/2xzaS+XqCiwqopGlH6PCMwdeu/ydV8zZ12gNLTYYO7e25MENXn3QdgtGsANbGitZ
0NdiElFLiE8ieOIJeiSU4P+VFfrwoeqMSeVCFt+p3l01TNA2Ig6wWbhCbDKKnvz8aw1lwJgvKOZU
ud6wpGB+PnBJ7593GhB2z2e+SaLal2eaGbRI1zCf/KBwy7zWQ8icVW4FkEHQWczBMAvV2swb9FKI
qbu5dt74O98AC/z7zAPdcYWJjZjgTDMe8CMBFb8YmDoA3fF82X08k0QkbUosnnAURt9fDXi9BuDY
OaYNO80bgfiaX3yamL/p15LdliKwIPhnnaJwk9QU+wTHkMCWEf3wLjookGTOVgOK8JZObkK2si9f
Pis5IBJNq1KzjwFTJafxMp19xuXDK7xtcnBXheaM1Hf2MRG1Sk2fhnZzrSOZGymJ/D8E4b2JfGlN
LpLbpke5FWSADW4vUxrGjxz3m2EUGCz4TXYF+nbLRC9ctXC2By04rwryr6eBjXp8sHcImCwtDnF1
iz4zurlWbFpx57s2uRtNsErB9efg+PQ5SPu35TSmsRcx1cigDjXM3Ul2yTFN5x+C+C89bwBK7C5L
OsDrZv/XIiWxKMo9cSEVZrGIcUblCycXfcMToQ1ecDUNSRCQ5GwG19+LECN5BLOMI5yHyEkR85+m
YLzy3TQuJ9MTC+dASBIT6e1AvCOI+Cn9RRyUJqgMjBMsUfTO9xOu8K/IFOtrBflNAiroguEeohec
3uLwMxcm/ceYmMwWyvkQd4avfz6IzsvsF+KYPFCKlrwgs3vzFEXO/i0xN07sqeGbvyYvt93F6vlR
KfxbIx+Icp8X5QyFpIUWUJN8QFTudGnVLY9h83y+OARQ6PcjhiSNf+1jFRu6mVjYC+X0/heL1Mx0
BEteVuHLjeg5aZMtkoppW2IVMISBQhaUwVJnbVwi3ji2M5SUPF3olMHMiHo/vvmbucNaPnv6Q5+l
qNzg0CO4GdwKTopD1wqjc0U4s9l6EZAztCQzNlJGBCK/Hf01b4vY8F6OMW+C2/wcuDGcqTjq9A85
KuzJot0IDG0Bawe2PaPV0pLlp2pbqtiPCBzomVSu3bFsl1msXirM82OII3iMDPlxE/vj8QcDTYQY
W7WWmTLde7dU8aFUw7zWZr7OR+M6qLxG71P0elCZ3buRK6ssoUtP5M7rvL427rhJtZaLJ89Syasn
E6G7Onk4WfKjcbTeu7JF63Eu1BnOWgd5sfmS9jchIukdhc/zykCE/PU8arDe0sQhN4+tQccnHQmn
38LmXVqgRKuSiKB36jVRwThJNjgL/WW2ybYY+fcCX1BY1ekLd8KwvEn/t+agU7osuTWUBDiQYvP0
AvICj+cPPmf6bjd6Vs8Jxi6COFTofZNb5SAr7rDT/semFfZiZNcivijBdoUODec/Ba8M2WewE2OX
XMdZ5m19MK9YVvV7YvZhgbvVtgy4cWkHcHMFBl3FZyihNxXc5iGuYgliHFmRNGhfgximOxAgoOKc
49WwQYu4AVAz1TiWolnm+/rNQB+4lyBSNOfAPxEqFeD5lddeHrB7teMf/lG8OFEZ4XCTgTAMa0di
30nRyTP2COrXU/JZwpjLIToJKu6IHctn9s5wGNxQXaDs12WNlXm2MMWLUKcvRFwLLZ3O4t/cx3C7
c8oGwjPcYoEqkPkatVizqCPpKGqjFTdtZGIcR37iAPXGwFQXvcw+pt0xamVxqAA5LMmblTEWN+f5
iyCFToPtdAG/icrR4ed5MVobh/s8erSfERHteS6biR4ckAnAnL7mFJiRvTrjZVBGVafTAW/X1fc/
bgr7TQpAYFZK4QP2kmqswaOLNUuaaWnbSAvGoMfwoQohosmZzok/wjYLZqIwgpDE9jiDmPGqzGg2
/afOAlCNeQDD3AqtOzmT7cDiL+snh9/vtUrJjEL57McNWCORLIpJS4CWush0xGHemzWehukzRSPH
Fb7+GDUnCMhLcYOuKGm2uBppkdOzzGNoxuFZtb2Qs0YEdVkW7nvlyMpOwBQ80T0ILnNDU2tepts/
LTepMmsbxJ+yCmVt3vfdVUIWznOxo7SY7xccdbGw5NmG3y8oobCkeIDqR9x4AUnYhGGr+3+jwmx3
8lpDMJitAbJrTYTEjkTu7rQK7syQTpTNAlAACUlgFs+HWmzj2fI5W+fz5NXVnywLfglDMkgwO0X+
8Yh6LBokHl+tEVUc1W2D4qEVQw6oS39oBFxTi6j29loznv3Y8WjTxtMJvke0mDWY2pJqSgxlSOOs
djYo7gU42cIY4gNsS/y7FZdK0wuPw/dUz81FdHsDBEOi+CFmnoV0yTeN70TmuoUyo4dnL2e/mvO6
oueyR5MOFuCuo947QF+e2LVdUg72i59g5pqHd1weY5/a4jMSMiDBZtr0QyeKQRKWHvHREdr4R0U3
xk5t8+IH1ijb61qsf+Hc+VxscwbNob4VBoqDLRwXPUoFCq6e77RrQDQDfScFllrqQfgIs9ESacR9
rfi6FFl9pxysmuhEX2+BzOhSP/QwAocdGvJPQfLfstFm71RhQvrkW7hCqD/I2igXPBQvXZ1pMDah
prj82cirwf9M+Dj9HyZtGglbWgCFfUawtjAySAow8uZTppZGlCrEdGp98yU1GN8TjcvXkQcu4TBk
sV0jQBHbqeB2QxW1YnNu4x6a7V5qN97WkeafzqCURgWyxp92nXk9I9maekQ4I2Hsv4GsXZl0dL5r
AY65fcfEe1E5wEw4awXp02Xqo8kCsDJGkyGGBFBlrPgZu4jorZsUnFG/JSTeBChqzHhwnGZOouQd
oKx3xSJUO3OHkOUJddIg1cwonliN7cOHg+s+NC6R5OLiQ4tVX0UU6b3ADaVGZ2QFAHXmwBA+avtR
hGVEJvYze5Yrg1wemP84O30uDE7RIXbzFNrxna0ChwzGPIrYyoELyr/Fa4KTG87p13Dxseg17Mqn
grh9VLFM3zL7LuK98W8d3iSbxCXtRZRRowi3CgItmJb/tkA7+hntBa/4jD2JFFn2qAlTtjCRn1Aw
B0pyj+5X3W21AK2JDc5ahb30qtKZbEsfFxeTlKv/sm1dzxDas2pfRMtchWL4aRabgbf+bYlpzSdk
GcSaSSRammNPIIRVsuPhR0D9vLdAbK60ZeY95+QZcXV4TTDJ42gvtbjpmjKbTrkz/ki5NgV1rHYe
UBZs/hJ/R+CTvvZ1C4Rahn3uZL6LIVPnHo12cLcDQzsa7ZV9smzPp2whx1hLfQfOQ7dVKqHmOg0Q
68oEpRpclvEOSSKrW+4FyOh8CW/FlV7oWZB9prJZ+VJR8Y5OoV3vYuUMOgVftCfsJcsWk59WhNYV
VErSfnECXTpi1AFjxlaGDzXZery2W8m47kjVTfxh/aHTFmPcrh8ZPwCqtkreItgo8nC7eJuzZiNS
tr8TrxBpIaSi5HYQqKPXmvGTDx88m4p5Gg6q9p7Q2LQKgHy5THpJtM1FzrQYeCTcc2jLqn1PEJVT
4FW7Fp5j79ZmAuPQIHoPDw49DneRv7yZ7SITe8f0ndARGyAaShYNeL686ICIdNfZyaqllnQxARJQ
tNHXjr7Fql8VzGwHRzP0Jj/O0fzc1BmmT3q+4Cm0a0LyMFJ5pV58Ou6n9fXxViM8MT9xl89mXP9j
57ncHt2sSFvNmDl7QHim4dEU/vcGhRYHlqsWzdWVJbZmd1t+VQ9uhgC3bClnQKp5tJ42MbMWrPfL
8/r1M3DYzl0jc5tS4HJdiA/GmFev1jru3o8US2/IawyRkvcXWe2eKZx8Yf+UmwD09vf87dENbP0n
2XGOfcD+w5/gbzrvmwIn33ZrKcrSQpp4/mQM93MdQe/n4OvDMAbcqBijX7UEbz7yNOxuByk7UFMq
kfGcjPwO+3+VrVQAu+jFym5094tR6+Ny6G9qhhiINgPQP3qFRs8pU8iJzDcBVjy0n+SiSIaOjGhp
aHcDgtUGxGumiE94X4Fgh8bwrI/+9nEhfnTVVEReHJPCalNIZijOcVSIhb1Cukq1iLFMrs815bDI
8gZmuqscK9r9xMQbw5lJlj5K3LhBiyIjXbFm0AsBdazvYnibmJGHtvRXOgSxqiM+1J+YVIwLTP6d
6eWq/S4BaXu82Ko/ycJpRAy+kcqrFno42uBsuQ5e2RN3zFOqmz02FLUMhrmQwl5RR308k1BbcU8g
mlgN7/eiagtL9J+EBn7aWPhfXWVEgApYbf7NG5tBLG/z75zUm7pWodHdB9uJscbRIAhJGM/XkEKI
EtdTzypzw6Y8OzgvUTy2kUPSa3mPQPzOWG8wvnZX2UYXvFgSaSqsT4tPvF9o07CFDAt/sUv5nycT
/+lfFrwfDOUpxa+mA5ldCmiSr+QAmL9CTxtf7e8aqk/MOsEMdSANO/rF5W9JLkbkPabbLIDV7xRZ
iu1UvqtDF7u71+RjOYKp2Fsd52ObB6sFKDqjcWTgSjpIoRVbaX4ZJ2K1P0/+QfOptO66ZHKERcdY
G3V9ZJEbHiYXY1ppRVMSeFXJFFT3cAw3X1Dfq2Pd1IlOm6bT338FM8lqHd2UhimpHGRN9poZwS7D
kqBvvcwZxWj0pT/Jd5c3EWM5lIlXzvseNiZFYGZazLuF7ehOLXtnUHexStgda/o9jYQnJ+7nNVyV
1tmNBAxegc8FI3rCJL49V30i8jrJIOqSKt3Z07Q8Jn7ePp3kfbe0IMlB/F9Tv12uOeO2DOwfIpDP
EPkUsJjHXEXkIzDPa7zuPr+AzSp9c8B2lkMxQX7bMXVWXSUX+D9rAwwrnlX5GQEVm+VablwDo8oR
4VF8+xlNDlGkK1k+d7WeLEOfHM/z0NK4xYLf0vrVkIi16bFMxPKbftXrSy57xuCmOb/ZE2uUuVqx
KuJCDYMbS6tqirWiQnnvhQwFypcnMIPTe9nwUicRFVNsb0xVhtv6fgSzphKr43VbtUnEoCZ9KKu5
DFZyPL0MFTsRB1FH4TL5a5pf13EshNEFOZD70dXcOKdNohItr/XhdLkOLGho+XWDsBxFE1NCx6vv
Qu8+IW1ewduGXUKM1LmMY9qyQD7VTYLGpTil5YPss8pxb74j322wsJBMDlxh5IbUz0M53/2tZfbU
H+UMx9SgQEEquxx6PIw6cyDTmya+0LqHiy2B15o0dAp+35YY6yDvI9JlnSucoeniN5lQtF8Ulxwn
Uh/eSdoN23XiStO646jHgMjZECdB/DO1OR8/szs2M49+FpN4jXfCtXvl+8S55e3IT2PFCfIxvwzq
iq758lw5m7Y01HCwWen61WZI3BVn7GCHzZzLEmC6Zmxv9gOwCH33KOK78o6hgj4xvqziPb5CJ/G9
yrJixp4EkAsSSayQ0mft9O49oKP5UoAHpALrmBC2TI/JRExoB7fJNhCUtmHqWT/I8gaCRlGmEYIm
rLO0QBCkfShRrcNXZ0dJX4QIJoXZZtjocPAEpmn8T8c8Yle5JxoZEQlVQi07YaMxjBuSIDByqp0n
38cn8yeoYDvcVwWYMe3OmwYuN5FZhvjLRF1xe2wnD14fd2xo7QjnXRjBW49bqtjKG4TmAoqvnWH8
zogOsT3Mh92XMNARkTA1SCvJh7CsPgl+ciwOmRUVKzO8yDH02MSt1oAY117BUva6q+2pBilvDtsL
tKiZV0DYqz10qeS3l24ALUs8b5Llnfk9RWzJWv19YZ9E/uOO8DxVJkX/X5lhBPPfI1amUox2GU8G
V1chOTm8eAGx0fe43rAuxUVKEozd4X30JeXYq0IQ70HaApLwlHeA4HQuppDBOS2rYFzjBwxpK6Q0
mYSVO0Qn82y6eTS6IXdr4SBNn+JqhjK3fwmCyImKZbT75WI5AZcNJ09UP+iTEUALtCMGeRDIEUuZ
T2M08OgmSIPIPnaH5Ob7/ae+rOHJ/p4Tela4amsz2BTw+jVBLrbeYaibmdPli2rrOktoIVyV+Bvk
8Mk9uBjBn5eTO/OsZCOo6t2tjQrXuuITN7z+xdWk2ohTcI33Ne9MGdENUCyiWYGjdOy0D6sYWHK6
CcZfXzdHCaYmhnTcqqQFywWyMQsiLdCWiSstmTiWJZ+oMB6f8mFLS3cp7DN9DkIY4cwBHNFMjC+T
rRzQLKij+sdjPS3JqV5TIwNhzRainG2SDC3Xzs3AkNnYHwBrsH01fyJDFc5u0M8CI1t27LugyRUK
MeXDOzxQ2qR8f70/i6wA3J5KWXrgk/Dsukw0DAPnmOuZzYIrVsuqVFJeLNFmEK6qbx5/Wp2h8mxw
O6cpuUDm+6q/AVgZ1N/OabM0i48deOs5IT2qVjdpOus48+vm9f7++DI63WC9/2ui4hTKUOXVRRQI
NFev0XbQArniF9C+3HJ2vgDa3D+4SzXrQq3S3D99Y21xuqEhYCk30bRpB2CtCNIMcUSaavh/Kvjr
jR5tSKDtpiWIgzpzqY5nplnhV1SS+PXB17d4Ix37z5d6hlJvJRXXesJOBPbL67ot5mQSSPyHYlHT
nqJwmRHSIM5iLb1Akt2+fytxhck7eFmmlqKMohoiu9yGR+UREzyRlga69/WTriaYUMJ+io4l4+SF
EkXZ2radupLwDVDKGaR4X6LQt0e58LWyZhI9ARGoBk8VbUACNAc3EcwSngNELcDm9GR/pFllSxD+
hqdrMVIQUP7aKJpvna4Kd8E41kS61A3zQu8LAoCptu9pE836d8SbXOK6o5eLiBv6eCNH7eMC+qNl
oR+bg0O684EJGtrYwiPpkm689lgM5uRDJFfZD3IpnIgwDpL7DeWo8xQZabhiPAPAzT0MDPpDXJ2j
nGtT+2NfbnbOUDhxXpvqeFLFH87C3Sl03YFlfDnyzHKemU6P3oqNOPfAEmQ0cXsqpqVXYBB7t985
5lPHYcXzcvubFipZT5SCxIdqWRCS2o3inur4F9whsqETsqOqdWtxx+tA/8z6e/YOydHGd5O4Su2/
h6K8iUFMA82hJE9TfdqPsUEhOXirKDa8nJna0Z8fpbFq1MGE/h1Mb6GMQ8MKzOKiA0nR7slwlj//
RJMyakvnimNEBHGY53svq106KJ4DkU5LlxAs+3fAu1G940PfCpwMo94GxKOLDfX/KIhrzt5Uj60u
SiXYyKeL1pOpSAqXS1fMRilD6pBG/EhaJeV5JgAnnrcV9FuGEWBeL9eAkukIvMIBW/n1HvYTc2vo
DOcSANI1bnJt71PTocmVOrvtUpKIHaOVyWlgq58fATcyqitvhsyyvvgXlR/sMSLfnJpuH5Cp1F8w
aDi/b9rJeHYbLyoPxy5fznpRPPtTRNmYm6PR6CROBTVpK2trq1x+bJXQSTFh4mICMUOsSBxFTmel
9EAoDvkmDokZIRzCJJadWiEPuRTwgs+8K+qZsfIq1Pc4f+bmDFNfqjMsr2t/ZsyxQEai3+IxmZDi
UVALCco+g1P6m1/32O3dMiYJCQ8ujZdW+MgH8bEu0TczicS3AAgp+IJ7PO6KyreZtjUQ4EAEhwRv
IUgUe94pN7ZK67CbjMWyHdEiRNA7tUy45ySpO7TGP/30OZOyV2HQaNii5I7MUaGEW4ZGmlC8qUib
QTlMgmnqHeyX7wI4+8JOkdDvA+Yx+/J4mQg6VAwqNKkzH2QCR8pHSehrh5rI76Xciemf4AWRYN4O
Ovf2JSSIeXTLVHHAgEai4pgv0JfCbcmhvMoGxqKUQn9+EyeRUEY1Q/sXHh6fE5BCSuvSjZdUsFXn
dXjBmlWl9m6J+YmWqwCkPtjC7C6Jn8kJWxc/jW2YToDUPHwlowrdRkGhIu+DQ1f2trAaRCzHHP8g
a1YKjYpaDvgMx7ibyHNAoye2G9v1oc73iQxjfGvtxYfGA11zm9YBmVqxSLQYm9l/3/Zj7pxvDHyC
/YkhqGpQK1xcesmqhPAfXrmtenTV4yMmvtYjIInVCXYm9WRNy511wU+NoTfHr6KLkc8aZnlJuYSJ
efgvpQLzrPmw2FIWHNPtLap+kdYSDIrcAWOYAe8Ne4d/a4WVH7Cq+KmQKrxS/hkSWLm5dP2G0hGk
xkzSEkp/6mVBpMnCPoaIjfhFg6OmrM3shcGgZKnWQeh5rN0qTrAmgo6GXioMph2RYHs1YQsOuukz
iR/1psX5g4Ju1eZvRyEggXaH7Gmk1hHyfumTBjtJ+c3ewRpHNyTJhoA/qWPc48rkbQ2UMXNpy9aP
zNXLdcbCbGEJ5qmZwRehLiQJajMXSPUeVNeJIzUuXRPpUrae4pFoWS8NZ10tZRmLrkglZIv1lTjz
VlqFwva41Yx3/Cz0laxbXzsco7nl5X2591RypmLU6n7JaiM13O85CgB0RgaO3+rZIIQ4P5GgmS7X
+w1V1UKJpgm19O1sSuPeygXDcAw/1xVUUZFVYQBaQfSusJAEAnEZztlQxtGR1F03Aju+rGbRqIMw
TtCdf3U1BkBbA96hADd2lpW6OdlM5agwgs6IQ+vn7WykYLJGvSpiwNSy5HhpRdaWBZglOx+xFAIi
XHczoFx3HFED/Yq/1SJ3+Kq1Sbw1KxtnO71yjBTcsbQS40v1rYQMYnrq3wI4t8knTAX4YtiOs3sV
ZZBmoqCSg34OlZEtTyUVJCKPHk9Ir+AnUTrHb02/yWb3jaaPAYVIlPF45YaWLZQDDoqihnv5fUDV
NQhGK0OfM1vLhTCcEi2d3zfCO18xD/I0fJoZDm7fSReXPQHliAmKrATNIGdtckse4JHGbMHmSf4u
sB8X47rbM7vGwwCX9zemLfHcfhim4UNPqHRKj81ofHz7CpsqugLQEIBTTF0h5rkMkalkCBZTZ6Zl
xFlDOf+lOMSQznlQETSlMQPplbwjd5XI4EKuy/bkm36fAHc0fJ+2+0y7y9M6qxJGvFpG3hNsk82e
5218ATdrlCn23C//bahdV9zvTurax+GItbJuNElT5GcVSjyZEj4zv7QQlbmx+qTGxPTbmroUokn9
wGmczshhJ08aUyY3mQ1/j0OZoWouWKipLl5bb0JEiIzP6qR3JqnGxWih1iBE8y3p9vPu4iaGj0K4
2b/Wlp5ff2m8cwfJao8vTe1VHnC4ZHdguLr/K9wvc0BkU0sw06aUdAO4TH1HoweYClV7IE8rk+y2
bzb0G6p8KmrJby3ZR6J+5dsjclAlX0RS7ZFf5qdbzk1ARVvsuRZhpjfpX9OyZWkqtGOMxpet3T/t
8y+hL3LRGTdPLPHY52w+ShoMaWCy33ijpFGvvE84zI+eFHRaEOaRUSwLBRf52DxFBPsQA7Cs11kc
PE36vcj2mEbwufHO4d9iXiLuendk0QIqEjc/5zYROiI9aYPR/cTqK3vnr9oiXZH1lRMZe/wIAp9Q
zReKpeJXxgrdDhLP2b5Pm/dhCM4ePIXD5bh2SwRJ4Himu3lUSwP0uD6s/JLMUuT2xwrMWEloy4nK
MXGD2KlqqYERCkKZn7VjPtWaPX52EdOByYSrdjcein4zfXlNshfpIZfl0zZhu2Y5wYNklSZOaWOC
47sjBV4b72h1VTCclDaIrKu9joN79cHcK4OO+q0lAEzI+Tk30Z/BWviLM0zRv6f/srRBCZyz7J9g
Nxuu0w1eR9G5qpT9xp42jB636UhTRuKrF/8jceppMkc+AXGPhjak0mT8qX2/kfgKss2Z2p6dM/h9
OcZlmFrnUQwjVyJ768wDeG2//YY/ZFyXb1E3rZDVBpSmPpQUvbe1+6Qm4R53m+bXi+hBSrPgvYMy
iruz84ayTQTN8ayKTlSY1bWTizAwDnIHCZEEkdrfgvr7PFh4G+MWy26uSdtN78N4e792mrajKUFZ
Qf8qu6ITJ6FF0TcsKf+vDikCN7nIbxY6t8v2dKsD6PtV/hpHiV9D4tIEwf9hrWxCOLaob72rLJbX
3MPcZb0Mlr+whyRypyMSRxEfd7OuV6lb0IQlG4QGqYr7cdRSIDxGHrBqbTH+s5J6BPFFSY9K/0EQ
Mi6Z1pWbcWxYK3HvF1g2m2sxJ2tuPdrZi6hFAsbeY7J3cpTXylz+/b08x+BaWFErSEDRAYNEex2j
9SDutLh0Sa1XgSOkPPFmcyURqTVNv9pKoXiesIk0aMa7NqVg62h9L264HvAgxFAy6w8cCEFF55M0
C8k3VpP30u2yRRDKoU//5b7eysNh0I83w0ctT2v1PC1pC1jKQHF4H7wqivHNFoUBnyPc898a3Ant
oOsqxTarKyfj4yyIAyihsv237GUNtUzEVSljqDPLVDNkpGnkmObC6BbryuXLV5w+Zx0tGdfFheS+
2y43x5SdYuJsZm6MakByemZJ4A5eJR0Mm4EU9QxhaNo/wxLmTsDk4wErsIudJlQiQpYzxwAnc00e
uHpWZbc8Fm8W8/RJIEYgvaC5B2QzeXbzgPDPXqnMqi5ALDRZHZG3te7bE8nNxT0xntpSZrFt4Wmf
PuoYS4WRensjOrn+HphNKUuULMe/q4VvD2K5jb6/x/y+hwQslNIj0/a3tL6ISpP++2XTx9KBYoOR
Byoo/m7Q34k2hbvx5EWmeXh97V86e0/ysj24Vcyyf1pkMBbD8UQl2Lay77an3vXOtBilCVObOTIT
l9b2+iGtdlRnJ4Sp7+kk2//4F3At2iejeg1w+jrP4fNCCn1mrO6GeTuVMaPtPN7P0Ac2O26LrQiV
Y7OxX/odhYM6r67mPmj1DE35eDrU0NsYbhbRuldEZKNCD2ZQoc8E8kcqOa5JqRJGCr2N5rv+ZbOz
7nrMQNoVz7uVCApsBUn3EOGbchDzz5DzJ6cvhDVWy8dCR+ohV6VYuYUqVgEaedTWPGMRAOFu2TcM
OZluG8PCNdb4UUwZ57sUmqXScau1L2DbvAA6z2K/hk4XmNUtn0mkRzTRqSBJHs+OnR8mMY6WzMVm
e47u8aKLyPmmz1nstT4objZB4fSnuunT0OmSjF4w65owSjGpLyDCq6ZDWr++pD6F2eFY02+iwWOw
Hhs2ANNMkCPha27Qd5LvxlvfwgFsaavd+/TXCZPqO1whT64Z99dsrWxw8aXNxPeme5g0gSrjxfSu
pkO8/AzC3gnchdgg714Pt9IsSnq3Hiy5H04vvrxDhRdttLcnKhDhkRLNBbEaIAqDa652MDuY9rx9
rhXOMqPZkUCVwVWCIi8oPPmGg099zDnbDwBnXhKWaa3PSPKGNrzaysxcD9NQHmKICvAeXHRYcXpS
EI9Lb0DiOA5JZsrWU19JmTjWIQvNFsQN5hVY25gw81qrbNongIjDr0NtL+IMqOR/a7+znnSOaNmC
anp6iegoel+Q6Hvzl+Ltj4nx2c0/bmU17oW0czh7bFHkNU6n66yUxmNdcJJOpFCQejejd/f+D+ia
+L0DBVeD1lJEuU49hqgkykMv40BaImwPnQu3MdCycoGLmkI+ZlZSSZJ7+w/bDhVCTcmlZNWAlNgl
6hR536oUJa9W9utT1tVAMP9H07fNvb3yYhn3w54VMXFTbfJ7VV2njD7o6osVskvgyOj5E7/k6oJo
pzQqcpTq5Y8q3FppGZ0ZFU+bK3TDq72g7V6pMN5IR6Mq1D1njdnKl78LlhrjvCKnYwzqlD/EIoRW
sEMH1Kk0ZtJrj9/00uQbupM7mCVQdRyQ51uaNr520SyWuhG/lQgHPI9DxXHi0hGMhPD3bkpKmYiq
pyO/hM6cQZupNNPgUupr9G/0bVmXE6jTJc9wxPW2iO+3KIKNs/H/i2loQseY2I9ZAekT5dOSZCMI
1kPAXTkatJx8lhQ4xXw4EowmVMAkY0Nb5Rb6DUNwzrFZ6WbwtMnsPNqN0f3t7ww6v3UI7TNhmqB2
g8YGLiBWPS73sH367n52/oKDwbMq5eghsuyd0Q8mlOpnfgT4BuSQ2hQ/7PKLlyWbiJ6808NctgxC
3o0lsD0gekOIUfQ17O8vVI9TH6OccNhovFUHc1L+paV64QiGZNr9ALNYHs5yU68mCmSn4eS8+5r5
XYX7zyc4azPLzu9jnyabWP+w0gFf2+3DbLXuDj9twdZTzU6j8jVQEEZgDRdqg+VvUWlr1P6fr+cK
dSyFOUKfYZQdzkMsJ1THkVQmfWHEYw6CmiMz8mFGiDQky648ocbkb2oRFl629QjnjOX/oFBYmz8Z
qWBfcKbLRkrczUOp8Jh8f09jyDImnUbZWNXrOiz3lVEKFYM2R6gl1zGTikMFdpAmGjusUHJ4XZ1D
bXdfJAukQF3y5mObTRGUEcLE4Rg5/qVKwNAQO5u5PeLPMDRStOeCKcM8FfXCXB7pmwAL8LGiBzJU
ndFIsnGx5vDxjJXuX5wC85NmB7EB1FZdSPl33IL+0vi+yjVJPfHBdow1BLgQs7FPAU9+tOOf4s1j
bQosH5idS2//Gu74dZkjtjrG+ua/MzpRc2Tm+EWlbDFt/WS02CcJXWLbU4boGwbzC93rk0nKodaV
cLvty+DlRGB29mlEXUORLMyDIszzZa+jIddM2GxFmvmzTzdlIYOI/1x7Zi9n+lR4ljL+M0QKr2OU
wNmjaWAM8RVUuDALvY+Wc1HzLuqzqjwavdDqM0fetuk8NTHAQfgr+UdJRhuNElJ0jyajQde9Unab
WebMCtsQxVEdbU4QUEURVUmYv34C9KmJvB7S8CcTSFMixJJhnsrkrvlbdl8O116TJzFsTzWcJfsb
u5Oc4HOBrelHE4q7935tcdmr5sJeBkMBWCqfLD12g8ChKgUJJ76Vt/XS4jMXPuNuFI3LdvDHC+u4
5rWGlmp3ESpDCB018yyPR+gVEz5Jt99SrnLOfGSw4gODId+ea8IgQRWoohkhe/slDN0Ho+V1+iSX
xLC6PG17RxKNTL+2xYugOo2LY8aZgHNhFbRTQPmgw0OqlNJ4OytmA3F3M5wB5Mo9XLKtrLx9Ri8U
zt4828orhyRbOjlImFpUJQWEkgvlIQAjAwVLiWsq3SFCXcuxf0N47Q9zWwHRIsQC/gUDFiwfC21Y
vG9iDmDfrg0Q5eGSX9+fXJ53emeJg7JZI0HriMndJ4uz84+f65DEeC1EJT9alZly3suRTjcY6Jkz
h9eI+xbuzK20YWb7SbaHRrVt1DKEFTeo61UIEE+4JhxlM4o7KkWx4C6X/crXQwqEZQFfe5PW5nx1
a8U1e5WMUO6VScm0VpDchMs40nIkLl0a9tVAKI880pUTMQ2WRhVgnSE5tGHPFu1VSem7y+ABk45m
ntHbwqYYlIIdigNwZXyQV9Lx+hZC5/qHBhz2kT9NDWEtt9YgaMGkjT8LoDZPQS6ik7n/LnOUhmOn
GoXkJiy/SoJzQVR/e9glwy8k7oXcSOKBNaojbywAjb7kHUkxQkW4FxYBq7jmtXtfZrbWSbc+lGsg
hTSNCnYqgk1Jwjy/OhLALkbJ4bKABQaLd5SGrFglpQksZAGDEgjCufenheJn00ucVsutWQRggPSi
BkZ4iRR5jWaFbYc2SwIr9m7LIDnmrFLbb4pZL122vJ8hxA7G/LyDWjQOkCWK6e/G/nLZb9CI755q
ssufyaN6KeIQ+90BV0cdYV6pJt5cvuWLX95964CDrZsLKXk2A5VSxgJbp/p+zQOZUNt8g7khKk/F
/XeouUbX3yi+zfa+okZpkaDBQaJ7OiRXiAlfPfBd+3jS5p4Ps2dFwRWHC9BGMebQnx2GG9DglOKg
y4NYy2ptq4+HXlNeM4Vb7tUhpaKCTq07m+LulHnhItdC8g2vLilQcyi4fj0w281HyLzPQLs+qejB
atEVhyCS9z6K7x2cqjksmBiIw7W67mOcAAcweYe33zDv6bLs2zBRVR4XEO3OQn5PwfAVH+u7dbDU
qYWxxqDOtM/PQt1SoNo3V7meS0PjbMmIvgTbP+6KeynRzKqBXw0AsX89NDT1G/qtKR9rFbTZBMJD
XJxFtGtwmaVivSsACvjvqjIUCvb2n4m/AN6qAvZCQ6sw7grmO8adpea5KXAomDorkcq45X1BOdL8
6DoN9DMSOnyPrBSPqFPFptlQEmSRkrIB9FXRcFDp6fEZHXquH37ZS6KvOYzhiFemstYBhzQkxt2Q
xZx4Huo+Ik36fCxEqcQGFwaB+rZtGkUgZ6msdeYLBt+oJqUKimBQC7pnVTuzM7pA9WbQDN4vZLLO
uZjoQGqwVxJz3SFW2rtKmSyCe9x9HVA0ouFdT57zhZr1OKJL4KWv7AASPw49jP8jvtet+t+yRwJQ
ym16ge1Q26oI9sf9KyMBilOgJTU2Q5krZN2Rn8imi10A8Z9ypMXKowsfE3zFReVblkgFDXjVIN4h
Y5J/F7LC6lJ/BwQQgoh99eYMCXiAZ30bOd8SAwojNlcUYp6zsTzfAeyHCv8ubA10wepGQVTTdg29
5vWgnrAO0UQi+7lgW1RENO2LG/dG7FxVG6HTzioQR/25pbgQRN0+nHetNc36EednmbVsbRIV+qn8
Ie/UWFvkYnja2yjGtON+jOfbMHSnJ+4WMv1YzhhHJWQ0dfNV8JkTrP6zeSwsZp9EZQAClvEO6b63
49MJy1AGLKhXuRWNgQnY7Ymqwh5P3c5e4mo/8CWhkPJbaiRHkoNA2eOSUuLXlhMlVDeaEaRHzoQ3
PeqCrhfRqE54GlNuao/1lleR7fNu6sT/JPkaqJiMp8sxsMacAn9zxnMvT1qqUHaxG7jzb7rT0Fl0
DClbn1n+36Dki7FtaIpUR9cfjqyIE435LkMYCiWylQuUzfDG5RYHQrDUUy/ixjEt6YUO2AseCYbS
M597JeLLl/s4TcLeRdTHDbymcq9thHREhwX5NeJsKdrbs8r9z0OK2+T198NPtD4BBBpdM/Mrm5Vi
7UXoViXtVlfLRC4U5phF/Ceeyq2hkXPqhSyM1+k3tTRRVKvsTITw32xGxpY3CQbmgLudn+UacMFS
pYDdcRtIpgGLOp4mKyPwWn855fDtbpw6aiWMBm+/FishwQOyK5hOhqZhbRxtETniP9PCevPj0n8W
vDnwtzIK3TTLkm98McU278nbpPKl/zeLOmwZBLsRT3/EDi2/n232JcH/2pkSIYUvc//06zJfl1Ut
uaL8o91rHbPRxBWA6oNNUkFv+Wx3fP+cNmWJK9Q4T4nfrWAu8ia6M1UmeUGSMfEx6bTJmQHTUNEg
uZ0VkpsI6uxK2jaEMUUuIIg7vS3z95YxKnNrTMP392PaefLqcUGAQTrvjZgULX331eeNUEjwWFv2
UGULJjfw5YpJXB1ozsUARA6DRo1d4hozQaV8pRtafIp7fhlI94gaKyDafFGCsTCS6WLDbGFNTyfv
ZToEybT/0tFShU46Mo56RjGawuxFDTU00JEfCvnmh0QlJ/d4Rwz+/MRxjPWJiGozJI2UI9UZYHq+
m7acajx176dTfyNUcrR+V2u3g+EDzoRXEHLYNw7QM1cfnDvCof0JFzUbUyJcgT1/4uMMhXSq20Sw
NBhrlTN32VYxItnQ2yuY1mvg6JGzvg6VHIgnuNjCPmGqCN9+BSgfgIvwRZvAIowkpBRhog0IBA3a
0J/SQkhUPoCD8WAVWY61bkZ369vFoNnzPn5tsqw6JU+zbz0WWXhBUsBFrNTZcMrTsqFtpDNB4zSM
j/SM/9AQUn9BkAnvwmR/ZS/OFKM5ChtC6EDfzVI7ogfAXyDRkGwV9iI9BQTMwMzqNQAnk724Ydg7
e3O+GGdZfcF3cVFFQHIzp1JutEQyudUOsoah1J86dWYpl4Pnmjwrtn88G78xJObY16Rslh+w+Rrb
GMnfdPS5zGRlH7XiVJb4OSiZmQwlszmdZ+j2Yh3THeaDDxAlKM+QJYDrH+NG+nBJAo/5o7GtK8YY
HOOVUwLwuUzFn7zxDdR1EzR7SpWKir43gYVbvkBBsVci09xrB1/k0tkY8o45DMODJtJ6FldKpkDv
pRHjO1Jv1Q2refNlBoBYQmIuKbKqD1tVTxaT6lkXS7RHzXGofSqtLxgUXhkxlG7F/pTGf1y8oKXz
KLIuPoivSRLGSsXXX49EIVjBC9H0JRNcL2nEvf+SyC6D3A/eDEr99BcoFbKArMrP+Y3qo9jVrrdq
iG3cuTwT7e/NU972kWWFsHx3XIC06Ht2yU8yaREnOEFk3+VRVt4VCKs+y8vCPac3Kw7KbTbnWKcd
BCdNDQyBnsa68PRLU9U/W2tebuJN9SFcoBhLXOeV0/Ok/gJ2riuwy8rP+XUEYEmAZEB9MFdPscz9
BAKbZyrAkSnuxlqfjvuLV/dhWqT97x2CUlOz3xPNGZIo1An1wX2yw5gPWbEGYbOk0ZYS7eY9RP6g
g0r0jqhscsjbD1Yz/mUnSZr6O+i/IVSnb8jz4BcdPtyuNHt+/TZjTUeV30Qgg4kM+6ktvTgZpupY
H2j6WkDi9oy0uNNvfwJwdxiDtaaB5lIYM+sSP/m/Sg11VRG8coNhOa+paiccY4by6IdyNxrclay5
Us+qGNM4pX7O4jlqksZkdKZhN3Fz2k4t1yw8RvyMnucJSRNiclTU5M9MC5jkYFpcm7tTHNQri6HW
p/UTW4OfgNtJmlS8lYwwwo87wE7hik836VQMNI0o60yQFcFxO6X+8jdiSSKqLhSKIfNNumBrOSKz
NiojdBVNFx/RMauPlM836Kji4TGwsygUrbHoNMeMEqWo2wy2rwcI3mDZF8PjU8Bk8yALnv23IetE
Y9EoKOs4rnP2oVFbtWdHp31LeI3KDoAsitrU+Qx41rt9NcEsdZLCNITHzcTbA3yLJOqmtYf3FS1c
l7BWIa6eEI9qO6V40D1RW/gaQHrfyLAC4hihByF7ouszyETbDx1zH2W677D+Rn2Upf81HZdi7lRf
G7y+pSUnj3OBo3D/QOOkCffpkxmYBVnfhPLBf25R+52vmHI5/Mi5Aq0ugVMugcbuQskww1gDH7z8
VHfHwYIS7C5F/cxhMSTlKwA1ntmrFqcfzQApLmvd/KgRujizknle6IeiYWoMvfnZF/VzNP0Vq/4r
nx9i2SE1kxBY7OKbWRgbGyJEClmJz8A0IZuXdQ2n5ae2DnOfQYGWAHfOSQ//uOfFmu1N3dq8o2tV
pA7BfsPntH7sUtQoaaPtrQbn3rWx0uI7/eDLF5EiQqiih64+bUjzc69sY5xhbY1Ls+KsI7+sF0gb
c9KA6bd6KrkQkm/KYmJHUItcXobCNWp9sS2GT0rBzkHsqTLTd7v0slVAx+RS/M4/lg3hnyLe+j1T
Nns9QxD/TdPsMsEaxbu7lI76/ZjP/LG5HOSY6DxRe8UF0BybMnpS5R2RKBGeY4HZPXUTmqGT6sEL
imc57HqUGzu7S5x+0/UcVPTsBwW1+KTB4ejl1fMbHJidyXw6mU1iKCXeOziWrRKYNljLEWi2ilfW
jZT/q4n1vBh0lhIe9f30kKcsvPyNSAhJ1/zl35PHrUgyDDj5xZOMvKsDqWsUWOEWYIT4wNWcf+uv
GHp0AIBdCPVuOlmQe8pqVctIlR3N1g4+vPUoFtBU3xw+3DvZvufCNVYLLYMDOZ9vlKbjVacxJaoR
dxSQQYxEx17L3IsoiXftVvaGX8VhhOyTr3hMnFfM+/bQ/zF1uh/1KbuV9xs7OO/n0x1E061vgdWP
ZPsXSVuL2wFPyqBCW8hF2t+GK4/hm+ikoncOWFrN0HgjIFQ/2yCFVNCQZ/m5VdQYuZePgiR+JZKp
myVjRItQj1Q5gNMhjQv8JAgyG3NpVMz5cPnp4Rmx9ZvkrkB/BlxKr+EAEzVNl95bPY2YkmBTPNZB
cxWL73ttiD0uAQvqchdEcrTxGsK7SW+683eZChhmBldvMJQ0/OYnhUI2xeMeqyP9KaVIQ7tpbCU1
16iYeTIwy9h6cZQwy8x1rJK5suE5im7UberHKUlxQxZKX4qMS/xHNoW8t5STKM3AlB4e3Tq1VBiy
Y2QdFB35cGFkVtKGbF4vZZwca+0Gf+zA1SSjqTHsOSjCs2utTyqOTv+GH7ElCzpZNN8fYWCQEosR
buoNHsF7JY55Pv19hEoASA1VawztpeHn8pYk0AFHxx45R42SlAGghT0STvsvAqilNGG/BJF928MB
MfwY8t6QcZLQeRqiA2DkRPVo5wwRph3fS74kNFY3D9C8Don0tgPkON+0ImOI1QP7p74WQD6ZOwas
oezNeBHCitQBGAc/0nBc5/7t8ozLYCr/EhWl5Y83L1dRx8p7ThOwce5xS5kqBDVUJF8U8EnawW/J
2ozkRO2aV4NPWivv3K/Tpr07zuoBB7i2nKS9aMOrFTFkoXPcRpVsR99r2nY45LqZXTJWkyB8Z74H
8tCv4ZNv28SvlEHckaqx0tpzZPh6IMLzZd5EsjI19VHT4o9P9EIifHZMznL/nv9846cRG6TXOfwp
NH8AY7xnTwDe+9/u/k4P+0Wu2biCpiePhl4y3KahVugL9iwqo0epvTeai2A/1Wb/p3Eltbq4DfoF
S98kfBU+jo80G+ZZ6B+S7JD5MDyl5qbiIU+n+91G3m1D+RKSY/uZ5/0GBJ4yBIGQyiWWsDcZi1WP
mEQyDrN60y8oNv2u8tblQyjo+YlOTYBCSiD3J8eNcgThkZkZ7t0wor6cg6RRtWzTOhqt+IW03GEj
9cBHz0gJf5BjfgRdRJY96VMcnkFObO9Tg6D1NUUeLidGDlTzslhE0p9aYM2us4E6dfNawY2pjz6G
+smrDQUiUW0lWdV4dYWhVTjWV/2I+xNaea/gLXOHnP/kT2hqjD+WtRCExH0BE3IbIMyq7qXmF2uK
vitRLs6Xnq0UgVqEneSyoZ80LTsmKmoflb7S5/RQvGuiDOoHsIxasjA35iZ6wpj/ZaC76cCQTbhR
36Jw7fq51nH7WotASQgz7w9bWIc4GOn60vHSTHO6WefcFH0pGgYkU/+Sky81p24JHFnCOeNOcoG4
PEfDgCx7rVRNMfCQJtqqUQGGwMCtVFcveCQpNa7QijNLIBLg3xIui4u1irLPdlSBDcQFbwZkaTa8
sWdqhVUAXnY9B7LnDHUWE9JCRCSjb9d6G0XQX1muMdgZoX4/CM/AbsBKc5LfCq+7t0A2W8RvsiHR
lnp375Sl8WYY6+DCinTwCbKxhFfZJrDVZLGopr6KVKCBBeB4kBrwPIWpbietZGM1JAgUQBSw4/Pu
A6mam2bWPdzFofrxnDOHy9oTiRtLm4v5PB+8a+3J6Tf5XiPsYP9JRzbZKUu58OEI/hk2oFnhfANL
6rM9gj0zDhCvUPCmz42wwB/1DLTjVqU4H0PaKmnk86zFqwn1zvhjPz4MLR4Q9S/z0UF+ERhRFOrw
EcDTlcCospb7T7/qBoVaG+aT+UxSsE2pvu3XnZpd0wG+0ipTvwQEw2jPMFJ57d/zNJz1S3bu3ZwZ
Gm5flEWFtESvGbcsLl1reMrQ1CdUPUw+9/XOPokXK6cVfpnWUN+N6JWDoQLIHLi1E3PmRTLq+U2D
bfkurMpAi6yVA71knp9I4VWQSpMHDINAwy05kW7GUSsUa3gctpsAiD0jGOO8WefHhzoLFQ7Zk5sO
HbRlZm04g/mi1KuCB4oYawQmIz8hZB0hJRjDfKR3fWF7w+IShnCsUxTp9YOb7edH6ukroowAoux4
Y8wX9PmbFQl69DRo7Zq+GyZ2ZwrtOVSlYuHEa2/rVk/Vn7vb2wQIxEXL/EUJEa6tapVDpJF1pRkh
ce+A8jsNEfloSZcBOvSdCVoYzEH+e8SQETQ4iLfnWp0inCCaOw+xZR0DDCm0ypfH9WNmG8WI8Ikd
+jI1YWY5X07Xom7DKdl79V0NjReT2nw5xw8vSq9A0gjfzfH7kZDXxNuAO704zFPWrvvTn2LF9AKl
zKLbOE2e3HINlSAqcEWZDPmx7R2hwvKEH4DYw55Tz1mGkjHVusrTQbUGIkc/Xfv4Xr3GF5XrwvIY
TiNH5uUHrSnwlzohiADLS7mBVRFrOtQz+STg61CffBg0K4U/1kYZbsT2WONlg/IR7B76FaqMTHQz
ipBWeDI1zAbEVVIQVmpb5aypZ7ZL0HPGyeIf7wvQjKBh57VXHLPAOCaEc91lU7acAyjsdOGErZfl
u4aY7ZkoFI6fmxYyF284LBG4nLVzHU4vgkvaLeAFpjhUueMU3cRbVygOgSVfR/DpDySDJuI3KGQ+
SMHVGoxnsbnkZJEV7nR2T8qr3hfYeVCJqPVcd2wbdwlad474IIfFQZAu3A8PEsHfj1w+VrzZ1l/X
tRJLofHSqFroTBFoRoWFoWeuNfjBEr7KFS2kdXKSvvW/eRkEM6LRKRXgAmGy6yY5deugwzAdjayo
v1UheqBbOkBjph4UyfsYQ7HzLIyTjM0jNLBc85EwXItkU+8ZxmgGUhyYqVM9rR3SQTwyJstlBsUL
8w3e9ICKGvhAX7c3/uWL8qAt3fgXp1fNY0Iz5d+ik4U+OuhA4OhwptX8/CuYn+mFBvQ4JsFllaJy
n/ggCKs7YhlS78r6rRcyVCoZ4fbYs1e0JsW/xZXxvqorywUA5/fYBspFo2MlSEcNAmaXSkq3W9Pq
IApwBjB7Ig7ZVzNw872XkzQRcFMVvVERS5LVKr8OjdQDnZLsFRHT9l6p6q/Lt6vcWNba11JCTlB7
MY0r5SET5CnjWtT1CwcaAIJb+pKERwhG2HWNxqqPJiN/ia7B+56lvfo9SAIKma2FKmiCDZuqqsCa
sKTPEm7pUGm4d7n6i998Kt1XhCes7tSHQ/JcgN/8XhQzagNK1roZrQg7iBnkfbF/z1nJJksSyGT7
Seqm4LWltyYLq0tm4WEgunBzH4mV5pYVIfCVjmniMajNvTuGns9YmxhGtbMG/vTzCKUpWgFZqCDg
9IRZnHoVzHbLBWFY97lu8zHwFoXMGeoayYr+PudV9ADuv4bKXeDtuhoO1AHPzlHfMN3byZofCpOr
aS+PWVDOBb0huTgASBxyNkix2aZiUHmvjKQAmlCV7GBGUiZHMlekAfK4kkMk9vev+mLAbypQusKs
rh1Eh2I0MBQBlBGKM1S6rgsUu5fy3bTeoqY+j7vSF6pkv0DzztJloku5cgQU65hqAtigO6oiwOQy
OKU+QheEo0XkrQ==
`protect end_protected

